// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Dec  7 18:01:21 2021
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n25888, data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(352[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(360[15:20])
    
    wire pwm_setpoint_23__N_207, n12452, n12456, n12458, n12462, n12464, 
        n12468, n12470, n12474, n12476, n12480, n12482, n260, 
        n58952, n58951, n12488, n294, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n625, 
        n623, n622, n621, n77679;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n68099, n58950, n67902, n58949;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, RX_N_2, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n58948, n65854, n1319, n58144, n58313, n1784, 
        n1786, n1788, n1790, n1792, n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    wire [5:0]color_bit_N_502;
    
    wire n58947, n58161, n58946, n25, n34, n33, n24, n23, n22, 
        n21, n7, n20, n19, n19_adj_5713, n17, n16, n15, n13, 
        n12, n11, n10, n9, n18, n17_adj_5714, n2819, n16_adj_5715;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n15_adj_5716, n14, n13_adj_5717, n2, n58519, n32, n31, 
        n30, n29, n28, n27, n26, n14_adj_5718, n15_adj_5719, n16_adj_5720, 
        n17_adj_5721, n18_adj_5722, n19_adj_5723, n20_adj_5724, n21_adj_5725, 
        n22_adj_5726, n23_adj_5727, n24_adj_5728, n25_adj_5729, n25_adj_5730, 
        n24_adj_5731, n23_adj_5732, n22_adj_5733, n21_adj_5734, n20_adj_5735, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    
    wire n70721;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n58518, n19_adj_5736, n18_adj_5737, n17_adj_5738, n16_adj_5739, 
        n15_adj_5740, n14_adj_5741, n13_adj_5742, n12_adj_5743, n58312;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n4, n4928, n4927, n4926, 
        n4906, n4905, n4907, n4908, n4909, n4910, n4911, n4912, 
        n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
        n4921, n4922, n4923, n4924, n4925, n58517, n58311, n2872, 
        n11_adj_5744, n10_adj_5745, n9_adj_5746, n4938, n77776, n8, 
        n58945, n58944, n58516, n58515, n35808, n58310, n58160, 
        n58514, n58309, n6, n58943, n58513, n58308, n58159, n58942, 
        n58512, n58307, n58941, n58511, n58940, n58510, n58939, 
        n58509, n58306, n65859, n66003, n66002, n66001, n65855, 
        n66000, n65999, n66004, n65998, n65997, n65996, n65995, 
        n65994, n65993, n65992, n65991, n65856, n65990, n65989, 
        n65988, n65987, n65986, n65985, n65984, n65983, n65982, 
        n65981, n65980, n65979, n65978, n65977, n65976, n65975, 
        n65974, n65973, n65972, n65971, n65970, n65969, n65968, 
        n65967, n65966, n65965, n65964, n65963, n65962, n65961, 
        n65960, n65959, n65958, n65957, n65956, n65955, n65954, 
        n65953, n65952, n65951, n65950, n65949, n65948, n65947, 
        n65946, n65945, n65857, n65944, n65943, n65862, n65866, 
        n65867, n65868, n65869, n65870, n65873, n29286, n65876, 
        n65877, n65878, n65879, n65880, n65875, n65881, n65882, 
        n65883, n65884, n65885, n65886, n65887, n65888, n65889, 
        n65890, n65891, n65892, n65893, n65894, n65895, n65896, 
        n65897, n65898, n65899, n65900, n65901, n65902, n65903, 
        n65904, n65905, n65906, n65907, n65908, n65909, n65910, 
        n29249, n65911, n65912, n65913, n65914, n65915, n65916, 
        n65917, n65918, n65919, n65920, n65921, n65922, n65923, 
        n65924, n65925, n65926, n65927, n65928, n65929, n65930, 
        n65931, n65932, n65934, n65935, n65936, n65937, n65938, 
        n65939, n65858, n65940, n65941, n65942, n70705, n29176, 
        n26732, n65853, n70699, n58508, n58305, n58304, n58507, 
        n58303, n58158, n58302, n58506, n58301, n58157, n58938, 
        n58300, n58505, n58299, n58937, n58504, n58298, n70693, 
        n58503, n58297, n70925, n58296, n70687, n58502, n58295, 
        n4_adj_5747, n58294, n70681, n70679, n58936, n58935, n58934, 
        n58501, n58500, n58933, n58293, n58932, n58499, n58931, 
        n58930, n58498, n70675, n58497, n58292, n70663, n7_adj_5748, 
        n6_adj_5749, n5, n4_adj_5750, n3, n2_adj_5751, n8_adj_5752, 
        n6_adj_5753, n58929, n15_adj_5754, n8_adj_5755, n70983, n6_adj_5756, 
        n58928, Kp_23__N_612, n71769, \FRAME_MATCHER.i_31__N_2509 , 
        Kp_23__N_1748, n70613, n69006, n30143, n30139, n30136, n30133, 
        n30130, n30127, n30124, n30121, n68987, n30117, n30116, 
        n30115, n30114, n30113, n30112, n30111, n30110, n30109, 
        n30108, n30107, n30106, n30105, n30093, n30092, n30091, 
        n30090, n30089, n30088, n30087, n30086, n30085, n30084, 
        n30083, n30082, n30081, n30080, n30079, n30078, n30077, 
        n30076, n30074, n30073, n30072, n30071, n30070, n30069, 
        n30068, n30066, n30065, n30064, n30063, n30062, n30061, 
        n30060, n30059, n30058, n30057, n30056, n30055, n30054, 
        n30053, n30052, n30051, n30050, n30049, n30048, n30047, 
        n30046, n30045, n30044, n30043, n30042, n30041, n30040, 
        n30039, n30037, n30036, n30034, n30033, n30032, n30031, 
        n30030, n30029, n30028, n30027, n30026, n30025, n30024, 
        n30023, n30022, n30021, n30020, n30019, n30018, n30011, 
        n30010, n30006, n30005, n30001, n30000, n29999, n29998, 
        n29997, n29996, n29995, n29994, n29993, n29992, n29991, 
        n29990, n29989, n29988, n29984, n70607, n66893, n29968, 
        n29967, n29966, n29965, n29964, n29963, n45323, n29959, 
        n29958, n29957, n29956, n29954, n29947, n29945, n29943, 
        n29942, n29939, n29938, n29937, n29936, n29935, n29934, 
        n29933, n29932, n45315, n45313, n45215, n29913, n29912, 
        n45309, n29908, n45307, n29904, n45303, n45297, n45291, 
        n45289, n45285, n29877, n29874, n29870, n65132, n65134, 
        n29861, n29858, n29849, n29843, n29840, n45281, n45295, 
        n45293, n45299, n45321, n45389, n45377, n70919, n45373, 
        n7_adj_5757, n6_adj_5758, n5_adj_5759, n4_adj_5760, n22_adj_5761, 
        n76884, n19_adj_5762, n17_adj_5763, n16_adj_5764, n15_adj_5765, 
        n35278, n25_adj_5766, n13_adj_5767, n11_adj_5768, n9_adj_5769, 
        n8_adj_5770, n7_adj_5771, n6_adj_5772, n5_adj_5773, n4_adj_5774, 
        n78834, n30_adj_5775, n23_adj_5776, n21_adj_5777, n19_adj_5778, 
        n17_adj_5779, n16_adj_5780, n15_adj_5781, n13_adj_5782, n11_adj_5783, 
        n10_adj_5784, n9_adj_5785, n8_adj_5786, n7_adj_5787, n6_adj_5788, 
        n4_adj_5789, n70601, n69122, n7_adj_5790, n70597, n66225, 
        n15_adj_5791, n70591, n58927, n58926, n58925, n58924, n58923, 
        n70589, n58922, n4_adj_5792, n4_adj_5793, n58921, n58920, 
        n58919, n58918, n58917, n58916, n70587, n58915, n58914, 
        n67079, n58913, n11_adj_5794, n58912, n45345, n30770, n30766, 
        n30765, n30764, n70565, control_update, n30761, n30760, 
        n58911, n58910;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n30756, n58909, n70561, n58908, n45105, n30749, n30746, 
        n58907, n58906, n58905, n58904, n30738, n58496, n12450, 
        n30735, n30734, n30732, n30731, n30730, n239, n247, n258, 
        n284, n291, n299_adj_5795, n313, n322, n336, n337, n339, 
        n340, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, 
        n359, n460, n467, n475, n486, n7_adj_5796, n5218, n5215, 
        n30728, n30725, n70555, n30723, n3163, n30721, n30720, 
        n30719, n30718, n30717, n5_adj_5797, n30716, n30715, n30714, 
        n30713, n15_adj_5798, n11_adj_5799, n30704, n30703, n30702, 
        n30701, n30700;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, n30699, debounce_cnt_N_3833, n30698, n30697, 
        n30696, position_31__N_3836, n67037, n23186, n30679, n30677, 
        n30676, n30675;
    wire [1:0]a_new_adj_6018;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_6019;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5802, b_prev_adj_5803, debounce_cnt_N_3833_adj_5804, 
        n30674, n30673, n30672, n30671, position_31__N_3836_adj_5805, 
        n37146, n71685, n30670, n70547, n30669, n12_adj_5806, n11_adj_5807, 
        n10_adj_5808, n4_adj_5809, n3_adj_5810, n2_adj_5811, n30668, 
        n30667, n30666, n30665, n58872;
    wire [7:0]data_adj_6032;   // verilog/eeprom.v(23[12:16])
    
    wire n30664;
    wire [7:0]state_7__N_3918;
    
    wire n58871, n58870, n58869, n58868, n58867, n58866, n58865, 
        n58864, n291_adj_5812, n30663, n4_adj_5813, n70541, n5_adj_5814, 
        n58863, n58862, n6901, n29780, n58861, n58860, n58859, 
        n58858, n30631, n30630, n45363, n30629, n30628, n58857, 
        n58856, clk_out;
    wire [15:0]data_adj_6039;   // verilog/tli4970.v(27[14:18])
    
    wire n67002;
    wire [7:0]state_adj_6041;   // verilog/tli4970.v(29[13:18])
    
    wire n30624, n58855, n30622, n30617, n68695, n30616, n15_adj_5825, 
        n30601, n30591, n30587, n30586, n66998, n58854, n5_adj_5826, 
        n30583, n30582, n30581, n29777, n30580, n58853, n12486, 
        n30579, n30578, n30577, n58852, n30576, n58851, state_7__N_4319, 
        n30575, n29773, n9_adj_5827, n8_adj_5828, n7_adj_5829, n6_adj_5830, 
        n5_adj_5831, n30574, n70535, n30553, n58156, n58291, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n6_adj_5832, n6_adj_5833, n45146, n78239;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n29770, n45359;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n66992, n67733;
    wire [2:0]r_SM_Main_adj_6055;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_6056;   // verilog/uart_tx.v(33[16:29])
    
    wire n70913, n30515, n30514, n30513, n30512, n23023, n25794, 
        n66982;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n30511, n30510, n30509, n30508, n30507, n30506, n30505, 
        n30503, n30501, n30500, n30499, n30498, n30497, n30496, 
        n30495, n30494, n30493, n70529;
    wire [7:0]state_adj_6068;   // verilog/i2c_controller.v(33[12:17])
    
    wire n70527, enable_slow_N_4213, n8_adj_5845, n30488, n30487, 
        n29767, n30479, n8_adj_5846;
    wire [7:0]state_7__N_4110;
    
    wire n30477, n6705, n58495;
    wire [7:0]state_7__N_4126;
    
    wire n30456, n70519, n36861, n30430, n68961, n29764, n66166, 
        n77736, n70513, n58494, n731, n58143, n7759, n7758, n7757, 
        n7756, n7755, n7754, n828, n829, n830, n831, n832, n833, 
        n834, n70507, n861, n896, n897, n898, n899, n900, n901, 
        n927, n928, n929, n930, n931, n932, n933, n934, n935, 
        n936, n937, n938, n939, n940, n941, n942, n943, n944, 
        n945, n946, n947, n948, n949, n950, n951, n952, n953, 
        n954, n955, n956, n957, n58493, n960, n995, n996, n997, 
        n998, n999, n1000, n1001, n70501, n1026, n1027, n1028, 
        n1029, n1030, n1031, n1032, n1033, n1059, n78225, n1093, 
        n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
        n58809, n34_adj_5847, n1125, n1126, n1127, n1128, n1129, 
        n1130, n1131, n1132, n1133, n70497, n1158, n1193, n1194, 
        n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1224_adj_5848, 
        n1225_adj_5849, n1226_adj_5850, n1227_adj_5851, n1228_adj_5852, 
        n1229_adj_5853, n1230_adj_5854, n1231_adj_5855, n1232_adj_5856, 
        n1233_adj_5857, n78268, n1257, n58808, n58807, n58806, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
        n1301, n58805, n58804, n58803, n58802, n58801, n58800, 
        n58799, n58798, n1323, n1324, n1325, n1326, n1327, n1328, 
        n1329, n1330, n1331, n1332, n1333, n58797, n58796, n58795, 
        n78284, n1356, n58794, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n1422, n1423, 
        n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n1455, n22_adj_5858, n1490, n1491, n1492, 
        n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
        n1501, n70481, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1554, 
        n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
        n1597, n1598, n1599, n1600, n1601, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1653, n58793, n58792, n1688, n1689, 
        n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
        n1698, n1699, n1700, n1701, n58791, n1719, n1720, n1721, 
        n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
        n1730, n1731, n1732, n1733, n58790, n58789, n78340, n1752, 
        n1787, n1788_adj_5859, n1789, n1790_adj_5860, n1791, n1792_adj_5861, 
        n1793, n1794_adj_5862, n1795, n1796_adj_5863, n1797, n1798, 
        n1799, n1800, n1801, n1818, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n41543, n61, n41560, n1851, n85, 
        n76, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
        n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
        n1901, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
        n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
        n1932, n1933, n77878, n1950, n45257, n1985, n1986, n1987, 
        n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
        n1996, n1997, n1998, n1999, n2000, n2001, n70475, n2016, 
        n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, 
        n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
        n2033, n78132, n2049, n66902, n66900, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n66898, 
        n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
        n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, 
        n2131, n2132, n2133, n58492, n2148, n70469, n66896, n58491, 
        n58490, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
        n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
        n2198, n2199, n2200, n2201, n66892, n2214, n2215, n2216, 
        n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, 
        n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
        n2233, n58769, n2247, n58768, n58767, n58766, n70463, 
        n58489, n58488, n58765, n58764, n58763, n2282, n2283, 
        n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, 
        n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
        n2300, n2301, n2313, n2314, n2315, n2316, n2317, n2318, 
        n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
        n2327, n2328, n2329, n2330, n2331, n2332, n2333, n70461, 
        n58762, n58761, n2346, n58760, n58759, n58758, n58757, 
        n58487, n58756, n58755, n2381, n2382, n2383, n2384, n2385, 
        n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
        n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
        n58486, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
        n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
        n2427, n2428, n2429, n2430, n2431, n2432, n2433, n58754, 
        n58753, n77967, n2445, n58752, n58751, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n58750, n29_adj_5864, n2511, n2512, 
        n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
        n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
        n2529, n2530, n2531, n2532, n2533, n2544, n27_adj_5865, 
        n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
        n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
        n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, 
        n23_adj_5866, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2643, n2678, n2679, n2680, n2681, n2682, 
        n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
        n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
        n2699, n2700, n2701, n76043, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
        n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
        n2729, n2730, n2731, n2732, n2733, n70443, n78370, n2742, 
        n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, 
        n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
        n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
        n2801, n2808, n2809, n2810, n2811, n2812, n2813, n2814, 
        n2815, n2816, n2817, n2818, n2819_adj_5867, n2820, n2821, 
        n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
        n2830, n2831, n2832, n2833, n2841, n70437, n2875, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n76037, n2907, n2908, n2909, n2910, n2911, n2912, 
        n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
        n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2929, n2930, n2931, n2932, n2933, n2940, n58485, n70431, 
        n78642, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
        n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
        n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
        n2998, n2999, n3000, n3001, n3006, n3007, n3008, n3009, 
        n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
        n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
        n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
        n58484, n3039, n70427, n58483, n3074, n3075, n3076, n3077, 
        n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, 
        n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
        n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
        n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
        n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
        n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
        n3129, n3130, n3131, n3132, n3133, n3138, n58482, n70419, 
        n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, 
        n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
        n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
        n3197, n3198, n3199, n3200, n3201, n3204, n3205, n3206, 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, 
        n3231, n3232, n3233, n3237, n58481, n78639, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
        n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, 
        n3301, n70413, n70407, n78567, n78549, n76880, n58480, 
        n58723, n58722, n24_adj_5868, n58479, n62, n58721, n58720, 
        n58719, n58478, n58477, n58718, n58717, n58716, n58715, 
        n58714, n58713, n70401, n58712, n58476, n58711, n58475, 
        n58710, n58709, n58474, n58708, n58707, n58473, n58706, 
        n58705, n58472, n58471, n13_adj_5869, n17_adj_5870, n32_adj_5871, 
        n34_adj_5872, n39, n41, n28271, n58470, n58469, n77405, 
        n28238, n70391, n58468, n28192, n58467, n58466, n58049, 
        n45327, n28172, n70385, n58465, n58687, n58686, n58685, 
        n58684, n44499, n58464, n58463, n58683, n58142, n28128, 
        n58682, n58681, n77824, n44644, n70381, n58680, n58462, 
        n58461, n58460, n28115, n58679, n58678, n28097, n9_adj_5873, 
        n16_adj_5874, n20_adj_5875, n22_adj_5876, n25_adj_5877, n33_adj_5878, 
        n37, n41_adj_5879, n70373, n21_adj_5880, n79029, n37_adj_5881, 
        n8_adj_5882, n10_adj_5883, n25_adj_5884, n79023, n39_adj_5885, 
        n79017, n38, n40, n24_adj_5886, n76916, n28074, n2_adj_5887, 
        n3_adj_5888, n4_adj_5889, n5_adj_5890, n6_adj_5891, n7_adj_5892, 
        n8_adj_5893, n9_adj_5894, n10_adj_5895, n11_adj_5896, n12_adj_5897, 
        n13_adj_5898, n14_adj_5899, n15_adj_5900, n16_adj_5901, n17_adj_5902, 
        n18_adj_5903, n19_adj_5904, n20_adj_5905, n21_adj_5906, n22_adj_5907, 
        n23_adj_5908, n24_adj_5909, n25_adj_5910, n26_adj_5911, n27_adj_5912, 
        n28_adj_5913, n29_adj_5914, n30_adj_5915, n31_adj_5916, n32_adj_5917, 
        n58677, n58459, n44573, n58676, n58675, n58674, n44534, 
        n70367, n78999, n58458, n58457, n58456, n76882, n58673, 
        n58672, n58455, n58671, n58670, n58454, n58453, n58155, 
        n58154, n58452, n58451, n70361, n28049, n59414, n59413, 
        n59412, n59411, n59410, n59409, n59408, n76924, n78993, 
        n45233, n25867, n28025, n70343, n67741, n65728, n58450, 
        n78981, n5_adj_5918, n79293, n70335, n25893, n58449, n58448, 
        n58447, n78320, n58446, n58445, n58444, n58443, n70329, 
        n58442, n58441, n58440, n70323, n58439, n70321, n70317, 
        n70315, n58646, n70313, n70311, n78969, n78963, n70305, 
        n58259, n58153, n70303, n6_adj_5919, n58258, n58257, n58256, 
        n70301, n58255, n58141, n51, n58254, n58253, n58252, n58251, 
        n58645, n58644, n58643, n58250, n58249, n58642, n58248, 
        n58247, n78957, n110, n44439, n70295, n70291, n77874, 
        n67642, n12_adj_5920, n58246, n78951, n58245, n70281, n58244, 
        n58243, n44122, n58242, n56, n38_adj_5921, n58241, n58240, 
        n69064, n27241, n70277, n27201, n58239, n58238, n58641, 
        n78945, n70265, n58640, n58639, n5_adj_5922, n8_adj_5923, 
        n7_adj_5924, n68995, n27004, n58638, n62242, n75904, n70257, 
        n78618, n67847, n70249, n58637, n58237, n26758, n58636, 
        n78615, n58635, n70243, n78939, n75908, n26873, n76598, 
        n58152, n70235, n58151, n78933, n76580, n4_adj_5925, n6_adj_5926, 
        n8_adj_5927, n9_adj_5928, n11_adj_5929, n13_adj_5930, n15_adj_5931, 
        n4_adj_5932, n6_adj_5933, n8_adj_5934, n9_adj_5935, n66388, 
        n58634, n58633, n75891, n58140, n38_adj_5936, n39_adj_5937, 
        n40_adj_5938, n41_adj_5939, n42, n43, n44, n45, n26329, 
        n58632, n58631, n58630, n58395, n12_adj_5940, n70229, n58394, 
        n70227, n66625, n70221, n66555, n66463, n29436, n68353, 
        n68798, n65874, n66040, n66039, n66038, n66037, n66036, 
        n65864, n65861, n66035, n66034, n66033, n65871, n65865, 
        n66032, n66031, n66030, n70215, n66029, n66028, n66027, 
        n66026, n66025, n66024, n66023, n66022, n66021, n66020, 
        n65872, n66019, n66018, n66017, n66016, n66015, n66014, 
        n66013, n66012, n66011, n65863, n28715, n28713, n28711, 
        n68999, n28701, n58393, n70211, n29153, n28662, n28660, 
        n28654, n58392, n58150, n71691, n58391, n70207, n26478, 
        n58390, n58389, n58139, n58388, n58387, n77630, n70197, 
        n78128, n20466, n11849, n11847, n58386, n58385, n37336, 
        n76616, n37335, n77589, n66010, n78576, n65078, n70191, 
        n70189, n20419, n67807, n34707, n77531, n78531, n78519, 
        n78513, n78507, n78498, n78489, n58384, n70179, n58383, 
        n77480, n75124, n75085, n75073, n78573, n70175, n67725, 
        n25771, n30318, n25774, n30314, n30308, n70165, n30304, 
        n29732, n29729, n30298, n30294, n25930, n78900, n70159, 
        n70153, n45383, n30265, n30262, n70147, n45353, n30259, 
        n30256, n30253, n30250, n30247, n76606, n77391, n70141, 
        n70137, n70135, n58614, n58613, n58612, n58611, n58610, 
        n58609, n58608, n58607, n58606, n58605, n58604, n58603, 
        n70119, n58602, n58601, n59170, n59169, n59168, n59167, 
        n70113, n59166, n58600, n59165, n59164, n59163, n59162, 
        n59161, n59160, n59159, n59158, n58599, n59157, n70107, 
        n59156, n59155, n59154, n59153, n70103, n59152, n59151, 
        n70101, n59150, n59149, n59148, n77284, n59147, n59146, 
        n59145, n77283, n59144, n59143, n59142, n59141, n59140, 
        n59139, n59138, n59137, n59136, n59135, n59134, n59133, 
        n59132, n59131, n78810, n77019, n44603, n59130, n59129, 
        n59128, n61786, n59127, n59126, n59125, n59124, n59123, 
        n59122, n59121, n59120, n70089, n59119, n59118, n59117, 
        n59116, n59115, n59114, n59113, n59112, n59111, n66240, 
        n59110, n59109, n41575, n70083, n59108, n78105, n59107, 
        n70077, n59106, n59105, n59104, n75775, n59103, n59102, 
        n75773, n59101, n59100, n70075, n58578, n58577, n58576, 
        n59099, n59098, n59097, n59096, n58575, n75767, n58574, 
        n58573, n59095, n59094, n59093, n59092, n59091, n59090, 
        n59089, n59088, n59087, n59086, n59085, n58572, n59084, 
        n58571, n58570, n59083, n59082, n58569, n70067, n58568, 
        n59081, n58149, n59080, n59079, n58567, n70061, n59078, 
        n59077, n59076, n59075, n59074, n59073, n59072, n59071, 
        n59070, n78807, n78804, n58566, n58565, n59069, n70055, 
        n59068, n59067, n58564, n59066, n75743, n59065, n59064, 
        n59063, n59062, n59061, n59060, n70051, n58148, n59059, 
        n59058, n59057, n59056, n59055, n59054, n59053, n59052, 
        n59051, n59050, n59049, n70045, n59048, n59047, n58138, 
        n70043, n76926, n59046, n59045, n59044, n76917, n59043, 
        n59042, n59041, n59040, n59039, n59038, n59037, n59036, 
        n59035, n59034, n58550, n59033, n58549, n58548, n59032, 
        n59031, n59030, n58547, n58546, n59029, n58545, n58544, 
        n59028, n59027, n59026, n59025, n59024, n59023, n13_adj_5941, 
        n59022, n19_adj_5942, n21_adj_5943, n23_adj_5944, n25_adj_5945, 
        n59021, n29_adj_5946, n33_adj_5947, n61_adj_5948, n59020, 
        n59019, n58147, n59018, n70029, n59017, n59016, n59015, 
        n59014, n59013, n59012, n70027, n70025, n59011, n59010, 
        n59009, n59008, n59007, n59006, n59005, n70023, n59004, 
        n57846, n58146, n59003, n59002, n58543, n36173, n58167, 
        n58542, n59001, n70021, n70019, n12454, n59000, n58166, 
        n58541, n12448, n58137, n58540, n58999, n75045, n20493, 
        n58539, n12460, n58998, n58997, n70017, n58538, n58537, 
        n70015, n65933, n75043, n12466, n70013, n7_adj_5949, n12472, 
        n71784, n70011, n7_adj_5950, n71787, n58996, n75039, n76659, 
        n7_adj_5951, n58995, n75037, n12478, n58994, n71907, n71763, 
        n75029, n12484, n70005, n71766, n71799, n75016, n70001, 
        n12490, n71808, n71688, n7_adj_5952, n58993, n65860, n58992, 
        n20465, n75007, n71686, n66009, n66008, n58991, n21156, 
        n58990, n66007, n58989, n58988, n21152, n58987, n78071, 
        n58986, n58985, n58984, n78768, n66006, n60808, n11912, 
        n61349, n58145, n58983, n58982, n58981, n58980, n58979, 
        n10_adj_5953, n66005, n58978, n25404, n58977, n65754, n58976, 
        n69022, n58165, n25769, n58975, n58974, n20420, n60716, 
        n58164, n58973, n58972, n78418, n76617, n58971, n68771, 
        n58970, n58969, n58968, n69169, n58967, n58966, n60685, 
        n58163, n58162, n58965, n76662, n61123, n61318, n58964, 
        n60656, n78030, n58963, n6_adj_5954, n60646, n58962, n68385, 
        n58961, n77530, n78023, n58960, n25910, n58959, n58958, 
        n58957, n58956, n25883, n76011, n77437, n58955, n58954, 
        n58953, n76658, n76673, n76672, n71912, n71908, n77229, 
        n71888, n68824, n17_adj_5955, n25_adj_5956, n64260, n24_adj_5957, 
        n5_adj_5958, n64350, n71361, n15_adj_5959, n14_adj_5960, n66244, 
        n67816, n14_adj_5961, n13_adj_5962, n66150, n66270, n6_adj_5963, 
        n74657, n66894, n78741, n74640, n66450, n69083, n74617, 
        n74616, n66644, n78310, n74609, n69709, n74890, n66660, 
        n74606, n69703, n66769, n14_adj_5964, n10_adj_5965, n74590, 
        n69697, n74589, n76779, n66791, n69693, n69687, n6_adj_5966, 
        n5_adj_5967, n66842, n69681, n69677, n69671, n69665, n12_adj_5968, 
        n11_adj_5969, n10_adj_5970, n4_adj_5971, n69661, n69655, n69649, 
        n69645, n69639, n67720, n69633, n69629, n4_adj_5972, n69623, 
        n71810, n66590, n69617, n69613, n69607, n76778, n71801, 
        n69601, n66594, n69597, n69591, n69585, n66680, n67722, 
        n67779, n65094, n71789, n71786, n65130, n67822, n67837, 
        n77940, n65142, n65146, n65150, n65154, n67871, n65160, 
        n65164, n65168, n65172, n65176, n71771, n9_adj_5973, n71768, 
        n71767, n71764, n71755, n71754, n65244, n69523, n67787, 
        n69517, n8_adj_5974, n65268, n65272, n65276, n66788, n69276, 
        n65318, n65336, n74462, n65360, n7_adj_5975, n69038, n65398, 
        n78264, n69459, n69425, n74445, n71189, n74442, n77637, 
        n67763, n67800, n69383, n66751, n67825, n71492, n78729, 
        n7_adj_5976, n4_adj_5977;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n28025), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n59010), .I0(n2925), 
            .I1(VCC_net), .CO(n59011));
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .neopxl_color({neopxl_color}), 
            .\color_bit_N_502[1] (color_bit_N_502[1]), .state({state}), 
            .GND_net(GND_net), .bit_ctr({Open_0, Open_1, Open_2, Open_3, 
            bit_ctr[0]}), .n60716(n60716), .n60685(n60685), .n7(n7), 
            .timer({timer}), .VCC_net(VCC_net), .\bit_ctr[1] (bit_ctr[1]), 
            .\bit_ctr[3] (bit_ctr[3]), .n29966(n29966), .t0({t0}), .n28192(n28192), 
            .\bit_ctr[4] (bit_ctr[4]), .n30582(n30582), .n30581(n30581), 
            .n30580(n30580), .n30579(n30579), .n30578(n30578), .n30577(n30577), 
            .n30576(n30576), .n30575(n30575), .n30574(n30574), .n30553(n30553), 
            .n30477(n30477), .n65078(n65078), .NEOPXL_c(NEOPXL_c), .n44603(n44603), 
            .\color_bit_N_502[2] (color_bit_N_502[2]), .n3163(n3163), .n25404(n25404), 
            .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 mux_3812_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5731), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n59009), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62923 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[20] [0]), .I2(\data_out_frame[21] [0]), 
            .I3(byte_transmit_counter[2]), .O(n78807));
    defparam byte_transmit_counter_0__bdd_4_lut_62923.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n59009), .I0(n2926), 
            .I1(VCC_net), .CO(n59010));
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n59008), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n78807_bdd_4_lut (.I0(n78807), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[2]), 
            .O(n78810));
    defparam n78807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n59008), .I0(n2927), 
            .I1(VCC_net), .CO(n59009));
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n59007), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n59007), .I0(n2928), 
            .I1(VCC_net), .CO(n59008));
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n59006), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n59006), .I0(n2929), 
            .I1(GND_net), .CO(n59007));
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n59005), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n59005), .I0(n2930), 
            .I1(GND_net), .CO(n59006));
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n59004), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n59004), .I0(n2931), 
            .I1(VCC_net), .CO(n59005));
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n59003), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(n5_adj_5958), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n70401));
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5751), .I1(n7754), 
            .I2(n70401), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i61820_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[0] [7]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n65398));   // verilog/coms.v(94[13:20])
    defparam i61820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15665_3_lut (.I0(\data_in_frame[0] [6]), .I1(rx_data[6]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n29877));   // verilog/coms.v(130[12] 305[6])
    defparam i15665_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15662_3_lut (.I0(\data_in_frame[0] [5]), .I1(rx_data[5]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n29874));   // verilog/coms.v(130[12] 305[6])
    defparam i15662_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15658_3_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(n28701), .I3(GND_net), .O(n29870));   // verilog/coms.v(130[12] 305[6])
    defparam i15658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [6]), .I1(n45257), .I2(n28701), 
            .I3(rx_data[6]), .O(n65130));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i11_4_lut_adj_1764 (.I0(\data_in_frame[23] [5]), .I1(n45257), 
            .I2(n28701), .I3(rx_data[5]), .O(n65132));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_1764.LUT_INIT = 16'hca0a;
    SB_LUT4 i15649_3_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(n28701), .I3(GND_net), .O(n29861));   // verilog/coms.v(130[12] 305[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15646_3_lut (.I0(\data_in_frame[23] [3]), .I1(rx_data[3]), 
            .I2(n28701), .I3(GND_net), .O(n29858));   // verilog/coms.v(130[12] 305[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31177_2_lut (.I0(n45146), .I1(n41543), .I2(GND_net), .I3(GND_net), 
            .O(n45257));
    defparam i31177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut_adj_1765 (.I0(\data_in_frame[23] [2]), .I1(n45257), 
            .I2(n28701), .I3(rx_data[2]), .O(n65134));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_1765.LUT_INIT = 16'hca0a;
    SB_LUT4 i62297_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78132));
    defparam i62297_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15637_3_lut (.I0(\data_in_frame[0] [3]), .I1(rx_data[3]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n29849));   // verilog/coms.v(130[12] 305[6])
    defparam i15637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15631_3_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(n28701), .I3(GND_net), .O(n29843));   // verilog/coms.v(130[12] 305[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut (.I0(color_bit_N_502[2]), .I1(n60716), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i59016_4_lut (.I0(bit_ctr[0]), .I1(n7), .I2(n60685), .I3(color_bit_N_502[1]), 
            .O(n74640));   // verilog/neopixel.v(34[12] 113[6])
    defparam i59016_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i26_4_lut (.I0(n25404), .I1(n74640), .I2(state[1]), .I3(n4_adj_5977), 
            .O(n65078));   // verilog/neopixel.v(34[12] 113[6])
    defparam i26_4_lut.LUT_INIT = 16'hfaca;
    SB_LUT4 i15628_3_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(n28701), .I3(GND_net), .O(n29840));   // verilog/coms.v(130[12] 305[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16267_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n28074), .I3(GND_net), .O(n30479));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16275_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n28074), .I3(GND_net), .O(n30487));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22987_3_lut (.I0(n313), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n37146));
    defparam i22987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n37146), .I2(n28074), 
            .I3(GND_net), .O(n30488));
    defparam i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16281_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n28074), .I3(GND_net), .O(n30493));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5732), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16282_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n28074), .I3(GND_net), .O(n30494));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i23179_3_lut (.I0(n239), .I1(n291), .I2(n284), .I3(GND_net), 
            .O(n37335));
    defparam i23179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23180_3_lut (.I0(n37335), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n37336));
    defparam i23180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5729));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n37336), .I2(n28074), 
            .I3(GND_net), .O(n30495));
    defparam i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16284_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n28074), .I3(GND_net), .O(n30496));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5728));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n59003), .I0(n2932), 
            .I1(GND_net), .CO(n59004));
    SB_LUT4 i16285_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n28074), .I3(GND_net), .O(n30497));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16286_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n28074), .I3(GND_net), .O(n30498));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16287_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n28074), .I3(GND_net), .O(n30499));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16288_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n28074), .I3(GND_net), .O(n30500));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22652_3_lut (.I0(n322), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n347));
    defparam i22652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22653_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n28074), .I3(GND_net), .O(n30501));
    defparam i22653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62433_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78268));
    defparam i62433_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n59002), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16291_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n28074), .I3(GND_net), .O(n30503));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22699_3_lut (.I0(n247), .I1(n299_adj_5795), .I2(n284), .I3(GND_net), 
            .O(n36861));
    defparam i22699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30353_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i30353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n59002), .I0(n2933), 
            .I1(VCC_net), .CO(n59003));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5727));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22700_3_lut (.I0(n36861), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n349));
    defparam i22700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16293_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n28074), .I3(GND_net), .O(n30505));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16294_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n28074), .I3(GND_net), .O(n30506));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16295_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n28074), .I3(GND_net), .O(n30507));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16296_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n28074), .I3(GND_net), .O(n30508));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16297_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n28074), .I3(GND_net), .O(n30509));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16298_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n28074), .I3(GND_net), .O(n30510));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16299_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n28074), .I3(GND_net), .O(n30511));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16300_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n28074), .I3(GND_net), .O(n30512));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5726));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16301_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n28074), .I3(GND_net), .O(n30513));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16302_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n28074), .I3(GND_net), .O(n30514));   // verilog/motorControl.v(42[14] 73[8])
    defparam i16302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16303_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n23023), .I3(GND_net), .O(n30515));   // verilog/coms.v(130[12] 305[6])
    defparam i16303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[17] [4]), .I1(n28660), .I2(n28713), 
            .I3(rx_data[4]), .O(n65268));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1766 (.I0(\data_in_frame[17] [3]), .I1(n28660), 
            .I2(n28713), .I3(rx_data[3]), .O(n65272));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1766.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut (.I0(n8_adj_5845), .I1(n41543), .I2(GND_net), .I3(GND_net), 
            .O(n28660));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12_4_lut_adj_1767 (.I0(\data_in_frame[17] [2]), .I1(n28660), 
            .I2(n28713), .I3(rx_data[2]), .O(n65276));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1767.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_1768 (.I0(\data_in_frame[16] [7]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[7]), .O(n65142));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1768.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1769 (.I0(\data_in_frame[16] [4]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[4]), .O(n65094));
    defparam i12_4_lut_adj_1769.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_1770 (.I0(\data_in_frame[16] [3]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[3]), .O(n65146));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1770.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1771 (.I0(\data_in_frame[16] [2]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[2]), .O(n65150));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1771.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16218_3_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n28715), .I3(GND_net), .O(n30430));   // verilog/coms.v(130[12] 305[6])
    defparam i16218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1772 (.I0(n8_adj_5752), .I1(n41543), .I2(GND_net), 
            .I3(GND_net), .O(n28662));
    defparam i1_2_lut_adj_1772.LUT_INIT = 16'hbbbb;
    SB_LUT4 i12_4_lut_adj_1773 (.I0(\data_in_frame[16] [0]), .I1(n28662), 
            .I2(n28715), .I3(rx_data[0]), .O(n65154));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1773.LUT_INIT = 16'h3a0a;
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n59002));
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(GND_net), .I1(n2808), 
            .I2(VCC_net), .I3(n59001), .O(n2875)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n59000), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n59000), .I0(n2809), 
            .I1(VCC_net), .CO(n59001));
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n58999), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n58999), .I0(n2810), 
            .I1(VCC_net), .CO(n59000));
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n58998), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n58998), .I0(n2811), 
            .I1(VCC_net), .CO(n58999));
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n58997), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n58997), .I0(n2812), 
            .I1(VCC_net), .CO(n58998));
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n58996), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n58996), .I0(n2813), 
            .I1(VCC_net), .CO(n58997));
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n58995), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n58995), .I0(n2814), 
            .I1(VCC_net), .CO(n58996));
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n58994), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_151_14 (.CI(n58148), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n58149));
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n58994), .I0(n2815), 
            .I1(VCC_net), .CO(n58995));
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1774 (.I0(n347), .I1(Ki[1]), .I2(GND_net), .I3(GND_net), 
            .O(n110));
    defparam i1_2_lut_adj_1774.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(n78225), .I1(n1521), 
            .I2(VCC_net), .I3(n58519), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n58993), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n58518), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n58993), .I0(n2816), 
            .I1(VCC_net), .CO(n58994));
    SB_LUT4 i589_2_lut (.I0(n1319), .I1(n44439), .I2(GND_net), .I3(GND_net), 
            .O(n2819));   // verilog/TinyFPGA_B.v(384[18] 386[12])
    defparam i589_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n58992), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n58992), .I0(n2817), 
            .I1(VCC_net), .CO(n58993));
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i55666_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n71492));
    defparam i55666_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5725));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n58991), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n58991), .I0(n2818), 
            .I1(VCC_net), .CO(n58992));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819_adj_5867), 
            .I2(VCC_net), .I3(n58990), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62598_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6901), .I2(n71492), 
            .I3(n25_adj_5956), .O(n17_adj_5955));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i62598_4_lut.LUT_INIT = 16'h88ba;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n58990), .I0(n2819_adj_5867), 
            .I1(VCC_net), .CO(n58991));
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n58989), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5811), .I3(n58313), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n58989), .I0(n2820), 
            .I1(VCC_net), .CO(n58990));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5810), .I3(n58312), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n58139), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n58988), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5724));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n58312), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5810), .CO(n58313));
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n58988), .I0(n2821), 
            .I1(VCC_net), .CO(n58989));
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n58987), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n58987), .I0(n2822), 
            .I1(VCC_net), .CO(n58988));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5809), .I3(n58311), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n58147), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n58986), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i15893_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[1]), .I2(n5_adj_5797), 
            .I3(n25893), .O(n30105));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15894_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[2]), .I2(n5_adj_5826), 
            .I3(n25893), .O(n30106));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15894_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n58311), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5809), .CO(n58312));
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n58986), .I0(n2823), 
            .I1(VCC_net), .CO(n58987));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n58985), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5723));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n58518), .I0(n1522), 
            .I1(VCC_net), .CO(n58519));
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n58985), .I0(n2824), 
            .I1(VCC_net), .CO(n58986));
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n58984), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n58984), .I0(n2825), 
            .I1(VCC_net), .CO(n58985));
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i15895_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[3]), .I2(n44573), 
            .I3(n25893), .O(n30107));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15895_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15896_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[4]), .I2(n5_adj_5814), 
            .I3(n25883), .O(n30108));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15896_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n58983), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15897_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[5]), .I2(n5_adj_5797), 
            .I3(n25883), .O(n30109));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15897_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5831), .I3(n58310), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n58517), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15898_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[6]), .I2(n5_adj_5826), 
            .I3(n25883), .O(n30110));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15898_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n58310), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5831), .CO(n58311));
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n58983), .I0(n2826), 
            .I1(VCC_net), .CO(n58984));
    SB_LUT4 i1_2_lut_adj_1775 (.I0(n347), .I1(Ki[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_5921));
    defparam i1_2_lut_adj_1775.LUT_INIT = 16'h8888;
    SB_LUT4 i15899_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[7]), .I2(n44573), 
            .I3(n25883), .O(n30111));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15899_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16341_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3163), .I3(GND_net), 
            .O(n30553));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15900_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[8]), .I2(n5_adj_5814), 
            .I3(n25867), .O(n30112));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15900_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5722));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15901_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[9]), .I2(n5_adj_5797), 
            .I3(n25867), .O(n30113));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15901_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15902_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[10]), .I2(n5_adj_5826), 
            .I3(n25867), .O(n30114));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15902_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15903_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[11]), .I2(n44573), 
            .I3(n25867), .O(n30115));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15903_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n58982), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n58982), .I0(n2827), 
            .I1(VCC_net), .CO(n58983));
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n58981), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n58981), .I0(n2828), 
            .I1(VCC_net), .CO(n58982));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n58980), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15904_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[12]), .I2(n5_adj_5814), 
            .I3(n25910), .O(n30116));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15904_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n58980), .I0(n2829), 
            .I1(GND_net), .CO(n58981));
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n58979), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n58517), .I0(n1523), 
            .I1(VCC_net), .CO(n58518));
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n58979), .I0(n2830), 
            .I1(GND_net), .CO(n58980));
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n58978), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n58516), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n58516), .I0(n1524), 
            .I1(VCC_net), .CO(n58517));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5721));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n58978), .I0(n2831), 
            .I1(VCC_net), .CO(n58979));
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n58977), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n58977), .I0(n2832), 
            .I1(GND_net), .CO(n58978));
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n58976), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5830), .I3(n58309), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n58976), .I0(n2833), 
            .I1(VCC_net), .CO(n58977));
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n58976));
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(n78340), .I1(n2709), 
            .I2(VCC_net), .I3(n58975), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n58974), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n58974), .I0(n2710), 
            .I1(VCC_net), .CO(n58975));
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n58515), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n58973), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n58515), .I0(n1525), 
            .I1(VCC_net), .CO(n58516));
    SB_LUT4 i31273_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n45353));
    defparam i31273_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n58973), .I0(n2711), 
            .I1(VCC_net), .CO(n58974));
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n58309), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5830), .CO(n58310));
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n58972), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n58514), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n58972), .I0(n2712), 
            .I1(VCC_net), .CO(n58973));
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n58971), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n58971), .I0(n2713), 
            .I1(VCC_net), .CO(n58972));
    SB_LUT4 mux_3812_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5735), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15905_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[15]), .I2(n44573), 
            .I3(n25910), .O(n30117));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15905_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28128), 
            .D(n1238), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n58970), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15909_3_lut (.I0(\data_in_frame[4] [0]), .I1(rx_data[0]), .I2(n66150), 
            .I3(GND_net), .O(n30121));   // verilog/coms.v(130[12] 305[6])
    defparam i15909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15912_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n66150), 
            .I3(GND_net), .O(n30124));   // verilog/coms.v(130[12] 305[6])
    defparam i15912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n58970), .I0(n2714), 
            .I1(VCC_net), .CO(n58971));
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n58969), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n58969), .I0(n2715), 
            .I1(VCC_net), .CO(n58970));
    SB_LUT4 i15915_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n66150), 
            .I3(GND_net), .O(n30127));   // verilog/coms.v(130[12] 305[6])
    defparam i15915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15918_3_lut (.I0(\data_in_frame[4] [3]), .I1(rx_data[3]), .I2(n66150), 
            .I3(GND_net), .O(n30130));   // verilog/coms.v(130[12] 305[6])
    defparam i15918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n58968), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n58968), .I0(n2716), 
            .I1(VCC_net), .CO(n58969));
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n58514), .I0(n1526), 
            .I1(VCC_net), .CO(n58515));
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n58967), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n58513), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16106_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n66992), .I3(GND_net), .O(n30318));   // verilog/coms.v(130[12] 305[6])
    defparam i16106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31393_4_lut (.I0(n829), .I1(n828), .I2(n45353), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i31393_4_lut.LUT_INIT = 16'heccc;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n58513), .I0(n1527), 
            .I1(VCC_net), .CO(n58514));
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n58967), .I0(n2717), 
            .I1(VCC_net), .CO(n58968));
    SB_LUT4 i16102_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n66992), .I3(GND_net), .O(n30314));   // verilog/coms.v(130[12] 305[6])
    defparam i16102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n58966), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5829), .I3(n58308), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n58512), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61817_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[11] [5]), 
            .I2(n66992), .I3(GND_net), .O(n65318));   // verilog/coms.v(94[13:20])
    defparam i61817_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n58308), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5829), .CO(n58309));
    SB_LUT4 i16096_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n66992), .I3(GND_net), .O(n30308));   // verilog/coms.v(130[12] 305[6])
    defparam i16096_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5828), .I3(n58307), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n58307), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5828), .CO(n58308));
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n58966), .I0(n2718), 
            .I1(VCC_net), .CO(n58967));
    SB_LUT4 i12_4_lut_adj_1776 (.I0(n71799), .I1(n71801), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n65728));   // verilog/coms.v(105[12:33])
    defparam i12_4_lut_adj_1776.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n58965), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n58965), .I0(n2719), 
            .I1(VCC_net), .CO(n58966));
    SB_CARRY add_151_13 (.CI(n58147), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n58148));
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n58964), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5827), .I3(n58306), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16092_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n66992), .I3(GND_net), .O(n30304));   // verilog/coms.v(130[12] 305[6])
    defparam i16092_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n58964), .I0(n2720), 
            .I1(VCC_net), .CO(n58965));
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n58963), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n58306), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5827), .CO(n58307));
    SB_LUT4 i61818_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[11] [2]), 
            .I2(n66992), .I3(GND_net), .O(n65336));   // verilog/coms.v(94[13:20])
    defparam i61818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16086_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n66992), .I3(GND_net), .O(n30298));   // verilog/coms.v(130[12] 305[6])
    defparam i16086_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n58963), .I0(n2721), 
            .I1(VCC_net), .CO(n58964));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5714));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n58962), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_adj_1777 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_1777.LUT_INIT = 16'h4444;
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n58962), .I0(n2722), 
            .I1(VCC_net), .CO(n58963));
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n58512), .I0(n1528), 
            .I1(VCC_net), .CO(n58513));
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n58511), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n58961), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n58511), .I0(n1529), 
            .I1(GND_net), .CO(n58512));
    SB_LUT4 i1_3_lut_adj_1778 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1778.LUT_INIT = 16'h1414;
    SB_LUT4 i16082_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n66992), .I3(GND_net), .O(n30294));   // verilog/coms.v(130[12] 305[6])
    defparam i16082_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n58961), .I0(n2723), 
            .I1(VCC_net), .CO(n58962));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5808), .I3(n58305), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n58960), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n58960), .I0(n2724), 
            .I1(VCC_net), .CO(n58961));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n58959), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n58305), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5808), .CO(n58306));
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n58959), .I0(n2725), 
            .I1(VCC_net), .CO(n58960));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5807), .I3(n58304), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n58958), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16362_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3163), .I3(GND_net), 
            .O(n30574));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16362_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n58958), .I0(n2726), 
            .I1(VCC_net), .CO(n58959));
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n58957), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n58510), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n58957), .I0(n2727), 
            .I1(VCC_net), .CO(n58958));
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n58510), .I0(n1530), 
            .I1(GND_net), .CO(n58511));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n58509), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n58956), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n58509), .I0(n1531), 
            .I1(VCC_net), .CO(n58510));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n58304), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5807), .CO(n58305));
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n58146), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n58956), .I0(n2728), 
            .I1(VCC_net), .CO(n58957));
    SB_LUT4 i16363_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3163), .I3(GND_net), 
            .O(n30575));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n58955), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5806), .I3(n58303), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n58955), .I0(n2729), 
            .I1(GND_net), .CO(n58956));
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n58954), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16364_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3163), .I3(GND_net), 
            .O(n30576));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16364_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n58954), .I0(n2730), 
            .I1(GND_net), .CO(n58955));
    SB_LUT4 i16365_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3163), .I3(GND_net), 
            .O(n30577));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16366_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3163), .I3(GND_net), 
            .O(n30578));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n58953), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n58953), .I0(n2731), 
            .I1(VCC_net), .CO(n58954));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n58303), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5806), .CO(n58304));
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28128), 
            .D(n1237), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i16367_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3163), .I3(GND_net), 
            .O(n30579));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16368_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3163), .I3(GND_net), 
            .O(n30580));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15921_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n66150), 
            .I3(GND_net), .O(n30133));   // verilog/coms.v(130[12] 305[6])
    defparam i15921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i25_3_lut (.I0(encoder0_position[24]), .I1(n8), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16369_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3163), .I3(GND_net), 
            .O(n30581));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16370_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3163), .I3(GND_net), 
            .O(n30582));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16371_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n23023), .I3(GND_net), .O(n30583));   // verilog/coms.v(130[12] 305[6])
    defparam i16371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n58952), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14935_2_lut (.I0(n28049), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14935_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5717), .I3(n58302), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61814_4_lut (.I0(commutation_state[1]), .I1(n23186), .I2(dti), 
            .I3(commutation_state[2]), .O(n28049));
    defparam i61814_4_lut.LUT_INIT = 16'hc5cf;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n58952), .I0(n2732), 
            .I1(GND_net), .CO(n58953));
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n58508), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n58508), .I0(n1532), 
            .I1(GND_net), .CO(n58509));
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n58951), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16374_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n23023), .I3(GND_net), .O(n30586));   // verilog/coms.v(130[12] 305[6])
    defparam i16374_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n58951), .I0(n2733), 
            .I1(VCC_net), .CO(n58952));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n58302), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5717), .CO(n58303));
    SB_LUT4 i16375_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n23023), .I3(GND_net), .O(n30587));   // verilog/coms.v(130[12] 305[6])
    defparam i16375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27444_4_lut (.I0(n61), .I1(n76), .I2(rx_data[5]), .I3(\data_in_frame[17] [5]), 
            .O(n41575));   // verilog/coms.v(94[13:20])
    defparam i27444_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27445_3_lut (.I0(n41575), .I1(\data_in_frame[17] [5]), .I2(reset), 
            .I3(GND_net), .O(n30591));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n58507), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n58507), .I0(n1533), 
            .I1(VCC_net), .CO(n58508));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n58301), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n58301), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n58302));
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n58951));
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(n77967), .I1(n2610), 
            .I2(VCC_net), .I3(n58950), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n58949), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n58949), .I0(n2611), 
            .I1(VCC_net), .CO(n58950));
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n58948), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n58948), .I0(n2612), 
            .I1(VCC_net), .CO(n58949));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n58947), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n58947), .I0(n2613), 
            .I1(VCC_net), .CO(n58948));
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n58946), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15924_3_lut (.I0(\data_in_frame[4] [5]), .I1(rx_data[5]), .I2(n66150), 
            .I3(GND_net), .O(n30136));   // verilog/coms.v(130[12] 305[6])
    defparam i15924_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n58946), .I0(n2614), 
            .I1(VCC_net), .CO(n58947));
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n58945), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n58945), .I0(n2615), 
            .I1(VCC_net), .CO(n58946));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5716), .I3(n58300), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n58944), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15927_3_lut (.I0(\data_in_frame[4] [6]), .I1(rx_data[6]), .I2(n66150), 
            .I3(GND_net), .O(n30139));   // verilog/coms.v(130[12] 305[6])
    defparam i15927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16389_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n23023), .I3(GND_net), .O(n30601));   // verilog/coms.v(130[12] 305[6])
    defparam i16389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16053_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n67037), 
            .I3(GND_net), .O(n30265));   // verilog/coms.v(130[12] 305[6])
    defparam i16053_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n58507));
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(n78284), .I1(n1422), 
            .I2(VCC_net), .I3(n58506), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n58944), .I0(n2616), 
            .I1(VCC_net), .CO(n58945));
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n58943), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15568_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n66998), .I3(GND_net), .O(n29780));   // verilog/coms.v(130[12] 305[6])
    defparam i15568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15565_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n66998), .I3(GND_net), .O(n29777));   // verilog/coms.v(130[12] 305[6])
    defparam i15565_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n58943), .I0(n2617), 
            .I1(VCC_net), .CO(n58944));
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n58942), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61819_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[0] [1]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n65360));   // verilog/coms.v(94[13:20])
    defparam i61819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5720));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15558_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n66998), .I3(GND_net), .O(n29770));   // verilog/coms.v(130[12] 305[6])
    defparam i15558_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5719));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15555_3_lut (.I0(\data_in_frame[20] [1]), .I1(rx_data[1]), 
            .I2(n66998), .I3(GND_net), .O(n29767));   // verilog/coms.v(130[12] 305[6])
    defparam i15555_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n58300), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5716), .CO(n58301));
    SB_LUT4 i15552_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n66998), .I3(GND_net), .O(n29764));   // verilog/coms.v(130[12] 305[6])
    defparam i15552_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5715), .I3(n58299), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n58942), .I0(n2618), 
            .I1(VCC_net), .CO(n58943));
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n58505), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5776));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n58505), .I0(n1423), 
            .I1(VCC_net), .CO(n58506));
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n58941), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n58504), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n58941), .I0(n2619), 
            .I1(VCC_net), .CO(n58942));
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5787));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n58940), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5785));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5779));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5778));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5777));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5765));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5767));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15931_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n66150), 
            .I3(GND_net), .O(n30143));   // verilog/coms.v(130[12] 305[6])
    defparam i15931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31279_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n45359));
    defparam i31279_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5715));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62449_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78284));
    defparam i62449_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n85), .I2(\FRAME_MATCHER.i [4]), 
            .I3(n66982), .O(n61));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5762));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5716));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5771));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5769));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i27429_4_lut (.I0(n61), .I1(n76), .I2(rx_data[6]), .I3(\data_in_frame[17] [6]), 
            .O(n41560));   // verilog/coms.v(94[13:20])
    defparam i27429_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i62132_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77967));
    defparam i62132_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i27430_3_lut (.I0(n41560), .I1(\data_in_frame[17] [6]), .I2(reset), 
            .I3(GND_net), .O(n30616));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1706_3_lut (.I0(n2511), .I1(n2578), 
            .I2(n2544), .I3(GND_net), .O(n2610));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5768));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1779 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n70277));
    defparam i1_2_lut_adj_1779.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n927), .I1(n70277), .I2(n928), .I3(n45359), 
            .O(n960));
    defparam i1_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5763));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16405_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n23023), .I3(GND_net), .O(n30617));   // verilog/coms.v(130[12] 305[6])
    defparam i16405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16050_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n67037), 
            .I3(GND_net), .O(n30262));   // verilog/coms.v(130[12] 305[6])
    defparam i16050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5773));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59289_4_lut (.I0(n11_adj_5768), .I1(n9_adj_5769), .I2(n7_adj_5771), 
            .I3(n5_adj_5773), .O(n75124));
    defparam i59289_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16047_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n67037), 
            .I3(GND_net), .O(n30259));   // verilog/coms.v(130[12] 305[6])
    defparam i16047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16044_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n67037), 
            .I3(GND_net), .O(n30256));   // verilog/coms.v(130[12] 305[6])
    defparam i16044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16041_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n67037), 
            .I3(GND_net), .O(n30253));   // verilog/coms.v(130[12] 305[6])
    defparam i16041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5770), .I1(current_limit[9]), 
            .I2(n19_adj_5762), .I3(GND_net), .O(n16_adj_5764));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5774));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i60837_3_lut (.I0(n4_adj_5774), .I1(current_limit[5]), .I2(n11_adj_5768), 
            .I3(GND_net), .O(n76672));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i60837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60838_3_lut (.I0(n76672), .I1(current_limit[6]), .I2(n13_adj_5767), 
            .I3(GND_net), .O(n76673));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i60838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59250_4_lut (.I0(n17_adj_5763), .I1(n15_adj_5765), .I2(n13_adj_5767), 
            .I3(n75124), .O(n75085));
    defparam i59250_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16038_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n67037), 
            .I3(GND_net), .O(n30250));   // verilog/coms.v(130[12] 305[6])
    defparam i16038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i61047_4_lut (.I0(n16_adj_5764), .I1(n6_adj_5772), .I2(n19_adj_5762), 
            .I3(n75073), .O(n76882));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61047_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59932_3_lut (.I0(n76673), .I1(current_limit[7]), .I2(n15_adj_5765), 
            .I3(GND_net), .O(n75767));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i59932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61570_4_lut (.I0(n75767), .I1(n76882), .I2(n19_adj_5762), 
            .I3(n75085), .O(n77405));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61570_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16035_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n67037), 
            .I3(GND_net), .O(n30247));   // verilog/coms.v(130[12] 305[6])
    defparam i16035_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i61571_3_lut (.I0(n77405), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n22_adj_5761));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i61571_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n58940), .I0(n2620), 
            .I1(VCC_net), .CO(n58941));
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n58939), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16418_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n23023), .I3(GND_net), .O(n30630));   // verilog/coms.v(130[12] 305[6])
    defparam i16418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n58939), .I0(n2621), 
            .I1(VCC_net), .CO(n58940));
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n65920));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1780 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n65921));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1780.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5717));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n58938), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n58299), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5715), .CO(n58300));
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n58938), .I0(n2622), 
            .I1(VCC_net), .CO(n58939));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1781 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n65922));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1781.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n58937), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n58937), .I0(n2623), 
            .I1(VCC_net), .CO(n58938));
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n58936), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1782 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n65923));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1782.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n58936), .I0(n2624), 
            .I1(VCC_net), .CO(n58937));
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n58935), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n58935), .I0(n2625), 
            .I1(VCC_net), .CO(n58936));
    SB_CARRY add_151_12 (.CI(n58146), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n58147));
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n58504), .I0(n1424), 
            .I1(VCC_net), .CO(n58505));
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n58503), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5714), .I3(n58298), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n58934), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n58934), .I0(n2626), 
            .I1(VCC_net), .CO(n58935));
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n58933), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1783 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n65924));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1783.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51118_3_lut (.I0(n4_adj_5750), .I1(n7756), .I2(n66893), .I3(GND_net), 
            .O(n66896));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62869 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n78741));
    defparam byte_transmit_counter_0__bdd_4_lut_62869.LUT_INIT = 16'he4aa;
    SB_LUT4 n78741_bdd_4_lut (.I0(n78741), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71888));
    defparam n78741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51119_3_lut (.I0(encoder0_position[28]), .I1(n66896), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62855 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n78729));
    defparam byte_transmit_counter_0__bdd_4_lut_62855.LUT_INIT = 16'he4aa;
    SB_LUT4 n78729_bdd_4_lut (.I0(n78729), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71912));
    defparam n78729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n58933), .I0(n2627), 
            .I1(VCC_net), .CO(n58934));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1784 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n65925));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1784.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1785 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n65926));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1785.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5850));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31209_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n45289));
    defparam i31209_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5783));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5782));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n58932), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n58932), .I0(n2628), 
            .I1(VCC_net), .CO(n58933));
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5781));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1786 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n65927));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1786.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n58931), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1787 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n65928));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1787.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1788 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n65929));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1788.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28128), 
            .D(n1236), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1789 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n66009));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1789.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1790 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n65862));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1790.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1791 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n66008));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1791.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5713));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5757));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1792 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n65859));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1792.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n65930));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1793.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1794 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n65931));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1794.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1795 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n65932));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1795.LUT_INIT = 16'h2300;
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28128), 
            .D(n1235), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28128), 
            .D(n1234), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5759));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1796 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n65933));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1796.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n58931), .I0(n2629), 
            .I1(GND_net), .CO(n58932));
    SB_LUT4 mux_3812_i6_3_lut (.I0(encoder0_position[5]), .I1(n27), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1797 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n65934));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1797.LUT_INIT = 16'h2300;
    SB_LUT4 i59210_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5757), .I3(n5_adj_5759), 
            .O(n75045));
    defparam i59210_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8_adj_5755));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28128), 
            .D(n1233), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7_adj_5757), 
            .I3(GND_net), .O(n6_adj_5758));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5755), .I1(n301), .I2(n19_adj_5713), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1798 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n65935));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1798.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1799 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n65936));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1799.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1800 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n65937));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1800.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n6_adj_5966));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i2_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1801 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n65938));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1801.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1802 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n65939));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1802.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_adj_1803 (.I0(duty[15]), .I1(duty[22]), .I2(n294), 
            .I3(GND_net), .O(n5_adj_5967));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i1_3_lut_adj_1803.LUT_INIT = 16'h7e7e;
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n58930), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28128), 
            .D(n1232), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28128), 
            .D(n1231), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28128), 
            .D(n1230), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i3_4_lut_adj_1804 (.I0(duty[16]), .I1(n5_adj_5967), .I2(n294), 
            .I3(n6_adj_5966), .O(n10_adj_5970));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i3_4_lut_adj_1804.LUT_INIT = 16'hffde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1805 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n65857));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1805.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1806 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n65940));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1806.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1807 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n65941));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1807.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n305), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1808 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n66007));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1808.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n66006));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n66005));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1811 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n66004));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1811.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n74445), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_5760));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1812 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n66002));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1812.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n65858));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n66001));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n58503), .I0(n1425), 
            .I1(VCC_net), .CO(n58504));
    SB_CARRY add_151_5 (.CI(n58139), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n58140));
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n58502), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n58930), .I0(n2630), 
            .I1(GND_net), .CO(n58931));
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n58929), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n12));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n58502), .I0(n1426), 
            .I1(VCC_net), .CO(n58503));
    SB_LUT4 i59204_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n75045), 
            .O(n75039));
    defparam i59204_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n58501), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61556_4_lut (.I0(n16), .I1(n6_adj_5758), .I2(n19_adj_5713), 
            .I3(n75037), .O(n77391));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61556_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5850), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i61045_4_lut (.I0(n12), .I1(n4_adj_5760), .I2(n15), .I3(n75043), 
            .O(n76880));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61045_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n58929), .I0(n2631), 
            .I1(VCC_net), .CO(n58930));
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n58928), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5955));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n58928), .I0(n2632), 
            .I1(GND_net), .CO(n58929));
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n58501), .I0(n1427), 
            .I1(VCC_net), .CO(n58502));
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n58500), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n58927), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n58927), .I0(n2633), 
            .I1(VCC_net), .CO(n58928));
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n58927));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n58298), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5714), .CO(n58299));
    SB_LUT4 i61695_4_lut (.I0(n76880), .I1(n77391), .I2(n19_adj_5713), 
            .I3(n75039), .O(n77530));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61695_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(GND_net), .I1(n2511), 
            .I2(VCC_net), .I3(n58926), .O(n2578)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n58925), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18), .I3(n58297), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61696_3_lut (.I0(n77530), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n77531));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61696_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61645_3_lut (.I0(n77531), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n77480));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61645_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n58297), .I0(encoder0_position_scaled[7]), 
            .I1(n18), .CO(n58298));
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n1029), .I1(n45289), .I2(n1030), .I3(n1031), 
            .O(n67725));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n58500), .I0(n1428), 
            .I1(VCC_net), .CO(n58501));
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n58499), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n58925), .I0(n2512), 
            .I1(VCC_net), .CO(n58926));
    SB_LUT4 i20506_3_lut (.I0(n67037), .I1(rx_data[0]), .I2(\data_in_frame[9] [0]), 
            .I3(GND_net), .O(n30664));   // verilog/coms.v(94[13:20])
    defparam i20506_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_3812_i7_3_lut (.I0(encoder0_position[6]), .I1(n26), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5806));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5733), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5807));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3812_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5730), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21115_3_lut_4_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4938));
    defparam i21115_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_3812_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5737), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5808));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5827));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5828));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5829));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(duty[20]), .I1(n10_adj_5970), .I2(duty[19]), 
            .I3(n294), .O(n12_adj_5968));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i5_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 mux_3812_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5746), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n934));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5855));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5855), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(duty[17]), .I1(duty[13]), .I2(n294), .I3(duty[21]), 
            .O(n11_adj_5969));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i4_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1816 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5813));
    defparam i1_2_lut_adj_1816.LUT_INIT = 16'heeee;
    SB_LUT4 i16453_3_lut (.I0(current[11]), .I1(data_adj_6039[11]), .I2(n28097), 
            .I3(GND_net), .O(n30665));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16453_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16454_3_lut (.I0(current[10]), .I1(data_adj_6039[10]), .I2(n28097), 
            .I3(GND_net), .O(n30666));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16454_3_lut.LUT_INIT = 16'hcaca;
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n58924), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16455_3_lut (.I0(current[9]), .I1(data_adj_6039[9]), .I2(n28097), 
            .I3(GND_net), .O(n30667));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16456_3_lut (.I0(current[8]), .I1(data_adj_6039[8]), .I2(n28097), 
            .I3(GND_net), .O(n30668));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16457_3_lut (.I0(current[7]), .I1(data_adj_6039[7]), .I2(n28097), 
            .I3(GND_net), .O(n30669));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61081_3_lut (.I0(n77480), .I1(n298), .I2(duty[12]), .I3(GND_net), 
            .O(n76916));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61081_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61082_4_lut (.I0(n76916), .I1(n294), .I2(n11_adj_5969), .I3(n12_adj_5968), 
            .O(n76917));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i61082_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n58924), .I0(n2513), 
            .I1(VCC_net), .CO(n58925));
    SB_LUT4 i16458_3_lut (.I0(current[6]), .I1(data_adj_6039[6]), .I2(n28097), 
            .I3(GND_net), .O(n30670));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51354_4_lut (.I0(n260), .I1(duty[23]), .I2(n294), .I3(n76917), 
            .O(n11847));
    defparam i51354_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i60202_3_lut (.I0(n15_adj_5781), .I1(n13_adj_5782), .I2(n11_adj_5783), 
            .I3(GND_net), .O(n76037));
    defparam i60202_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i16459_3_lut (.I0(current[5]), .I1(data_adj_6039[5]), .I2(n28097), 
            .I3(GND_net), .O(n30671));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16460_3_lut (.I0(current[4]), .I1(data_adj_6039[4]), .I2(n28097), 
            .I3(GND_net), .O(n30672));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n58923), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n58923), .I0(n2514), 
            .I1(VCC_net), .CO(n58924));
    SB_LUT4 i16461_3_lut (.I0(current[3]), .I1(data_adj_6039[3]), .I2(n28097), 
            .I3(GND_net), .O(n30673));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n58922), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n58499), .I0(n1429), 
            .I1(GND_net), .CO(n58500));
    SB_LUT4 i16462_3_lut (.I0(current[2]), .I1(data_adj_6039[2]), .I2(n28097), 
            .I3(GND_net), .O(n30674));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16463_3_lut (.I0(current[1]), .I1(data_adj_6039[1]), .I2(n28097), 
            .I3(GND_net), .O(n30675));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16464_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n23023), .I3(GND_net), .O(n30676));   // verilog/coms.v(130[12] 305[6])
    defparam i16464_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n58922), .I0(n2515), 
            .I1(VCC_net), .CO(n58923));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n58921), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n58921), .I0(n2516), 
            .I1(VCC_net), .CO(n58922));
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n58920), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n58498), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n58920), .I0(n2517), 
            .I1(VCC_net), .CO(n58921));
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n58919), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i60069_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n76037), .O(n75904));
    defparam i60069_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i59194_4_lut (.I0(n21_adj_5777), .I1(n19_adj_5778), .I2(n17_adj_5779), 
            .I3(n9_adj_5785), .O(n75029));
    defparam i59194_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n58919), .I0(n2518), 
            .I1(VCC_net), .CO(n58920));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n58918), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n58918), .I0(n2519), 
            .I1(VCC_net), .CO(n58919));
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n58917), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n58498), .I0(n1430), 
            .I1(GND_net), .CO(n58499));
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n58497), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n58917), .I0(n2520), 
            .I1(VCC_net), .CO(n58918));
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n58497), .I0(n1431), 
            .I1(VCC_net), .CO(n58498));
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n58496), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n58916), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n58296), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60208_4_lut (.I0(n9_adj_5785), .I1(n7_adj_5787), .I2(current[2]), 
            .I3(duty[2]), .O(n76043));
    defparam i60208_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i60771_4_lut (.I0(n15_adj_5781), .I1(n13_adj_5782), .I2(n11_adj_5783), 
            .I3(n76043), .O(n76606));
    defparam i60771_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n58916), .I0(n2521), 
            .I1(VCC_net), .CO(n58917));
    SB_LUT4 i16244_3_lut_4_lut_4_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(reset), .I3(n76), .O(n30456));   // verilog/coms.v(130[12] 305[6])
    defparam i16244_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n58915), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n58496), .I0(n1432), 
            .I1(GND_net), .CO(n58497));
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n58915), .I0(n2522), 
            .I1(VCC_net), .CO(n58916));
    SB_LUT4 i60763_4_lut (.I0(n21_adj_5777), .I1(n19_adj_5778), .I2(n17_adj_5779), 
            .I3(n76606), .O(n76598));
    defparam i60763_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n58914), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61394_4_lut (.I0(current[15]), .I1(n23_adj_5776), .I2(duty[12]), 
            .I3(n76598), .O(n77229));
    defparam i61394_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i11_3_lut_4_lut_4_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(reset), .I3(n76), .O(n65244));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_4_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i60073_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n77229), .O(n75908));
    defparam i60073_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5789));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i59908_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5781), .O(n75743));
    defparam i59908_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5775));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i60827_3_lut (.I0(n4_adj_5789), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n76662));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i60827_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n58914), .I0(n2523), 
            .I1(VCC_net), .CO(n58915));
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n58495), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n58913), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n58913), .I0(n2524), 
            .I1(VCC_net), .CO(n58914));
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n58912), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n58912), .I0(n2525), 
            .I1(VCC_net), .CO(n58913));
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n58495), .I0(n1433), 
            .I1(VCC_net), .CO(n58496));
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(reset), .I1(n41543), .I2(n8_adj_5752), 
            .I3(GND_net), .O(n28715));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i59055_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n75904), .O(n74890));
    defparam i59055_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n58911), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(n15_adj_5791), .I1(n23186), .I2(dti), 
            .I3(GND_net), .O(n28025));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_1817 (.I0(reset), .I1(n41543), .I2(n8_adj_5846), 
            .I3(GND_net), .O(n28711));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_1817.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_3_lut_adj_1818 (.I0(reset), .I1(n41543), .I2(n45146), 
            .I3(GND_net), .O(n28701));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_3_lut_adj_1818.LUT_INIT = 16'h4040;
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n58911), .I0(n2526), 
            .I1(VCC_net), .CO(n58912));
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n58910), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n58910), .I0(n2527), 
            .I1(VCC_net), .CO(n58911));
    SB_LUT4 LessThan_11_i35_rep_232_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n79293));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_232_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16484_3_lut (.I0(baudrate[15]), .I1(data_adj_6032[7]), .I2(n28271), 
            .I3(GND_net), .O(n30696));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n58909), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n58909), .I0(n2528), 
            .I1(VCC_net), .CO(n58910));
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n58495));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n58908), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n58908), .I0(n2529), 
            .I1(GND_net), .CO(n58909));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n58296), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n58297));
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5813), .I2(delay_counter[10]), 
            .I3(n25769), .O(n69083));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1819 (.I0(n69083), .I1(n25771), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n69169));
    defparam i2_4_lut_adj_1819.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5923));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i16486_3_lut (.I0(baudrate[14]), .I1(data_adj_6032[6]), .I2(n28271), 
            .I3(GND_net), .O(n30698));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16487_3_lut (.I0(baudrate[13]), .I1(data_adj_6032[5]), .I2(n28271), 
            .I3(GND_net), .O(n30699));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16488_3_lut (.I0(baudrate[12]), .I1(data_adj_6032[4]), .I2(n28271), 
            .I3(GND_net), .O(n30700));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16489_3_lut (.I0(baudrate[11]), .I1(data_adj_6032[3]), .I2(n28271), 
            .I3(GND_net), .O(n30701));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16490_3_lut (.I0(baudrate[10]), .I1(data_adj_6032[2]), .I2(n28271), 
            .I3(GND_net), .O(n30702));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62478_4_lut (.I0(n1026), .I1(n67725), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i62478_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16491_3_lut (.I0(baudrate[9]), .I1(data_adj_6032[1]), .I2(n28271), 
            .I3(GND_net), .O(n30703));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61602_3_lut (.I0(n30_adj_5775), .I1(n10_adj_5784), .I2(n75743), 
            .I3(GND_net), .O(n77437));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59938_4_lut (.I0(n76662), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n75773));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i59938_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i60823_3_lut (.I0(n6_adj_5788), .I1(duty[10]), .I2(n21_adj_5777), 
            .I3(GND_net), .O(n76658));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i60823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60824_3_lut (.I0(n76658), .I1(duty[11]), .I2(n23_adj_5776), 
            .I3(GND_net), .O(n76659));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i60824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60745_4_lut (.I0(current[15]), .I1(n23_adj_5776), .I2(duty[12]), 
            .I3(n75029), .O(n76580));
    defparam i60745_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5786), .I1(duty[9]), .I2(n19_adj_5778), 
            .I3(GND_net), .O(n16_adj_5780));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n58907), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n58907), .I0(n2530), 
            .I1(GND_net), .CO(n58908));
    SB_LUT4 i59940_3_lut (.I0(n76659), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n75775));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i59940_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_4_lut_adj_1820 (.I0(delay_counter[22]), .I1(n69169), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5924));
    defparam i2_4_lut_adj_1820.LUT_INIT = 16'ha8a0;
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n58906), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n58906), .I0(n2531), 
            .I1(VCC_net), .CO(n58907));
    SB_LUT4 i30593_4_lut (.I0(n7_adj_5924), .I1(delay_counter[31]), .I2(n25774), 
            .I3(n8_adj_5923), .O(n1319));   // verilog/TinyFPGA_B.v(380[14:38])
    defparam i30593_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i61091_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n75908), .O(n76926));
    defparam i61091_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i2_3_lut_adj_1821 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25771));
    defparam i2_3_lut_adj_1821.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n78268), .I1(n1323), 
            .I2(VCC_net), .I3(n58494), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i61754_4_lut (.I0(n75773), .I1(n77437), .I2(n79293), .I3(n74890), 
            .O(n77589));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61754_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i5_4_lut_adj_1822 (.I0(delay_counter[24]), .I1(delay_counter[27]), 
            .I2(delay_counter[28]), .I3(delay_counter[29]), .O(n12_adj_5920));
    defparam i5_4_lut_adj_1822.LUT_INIT = 16'hfffe;
    SB_LUT4 i61049_3_lut (.I0(n75775), .I1(n16_adj_5780), .I2(n76580), 
            .I3(GND_net), .O(n76884));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n58905), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n58905), .I0(n2532), 
            .I1(GND_net), .CO(n58906));
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n58493), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16492_3_lut (.I0(baudrate[8]), .I1(data_adj_6032[0]), .I2(n28271), 
            .I3(GND_net), .O(n30704));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61802_4_lut (.I0(n76884), .I1(n77589), .I2(n79293), .I3(n76926), 
            .O(n77637));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61802_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61795_4_lut (.I0(n77637), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n77630));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i61795_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i1_4_lut_adj_1823 (.I0(n77630), .I1(current[15]), .I2(duty[21]), 
            .I3(duty[20]), .O(n5_adj_5918));
    defparam i1_4_lut_adj_1823.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n5_adj_5918), .I1(duty[23]), .I2(n51), .I3(duty[22]), 
            .O(n11849));
    defparam i7_4_lut.LUT_INIT = 16'h3332;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n58493), .I0(n1324), 
            .I1(VCC_net), .CO(n58494));
    SB_LUT4 i6_4_lut (.I0(delay_counter[26]), .I1(n12_adj_5920), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n25774));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n58904), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1824 (.I0(delay_counter[3]), .I1(delay_counter[8]), 
            .I2(delay_counter[7]), .I3(GND_net), .O(n69122));
    defparam i2_3_lut_adj_1824.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1825 (.I0(delay_counter[1]), .I1(n69122), .I2(delay_counter[2]), 
            .I3(delay_counter[6]), .O(n12_adj_5940));
    defparam i5_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1826 (.I0(delay_counter[0]), .I1(n12_adj_5940), 
            .I2(delay_counter[5]), .I3(delay_counter[4]), .O(n25769));
    defparam i6_4_lut_adj_1826.LUT_INIT = 16'hfffe;
    SB_LUT4 i4978_4_lut (.I0(n25769), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5868));
    defparam i4978_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1827 (.I0(n24_adj_5868), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n68999));
    defparam i2_4_lut_adj_1827.LUT_INIT = 16'hc800;
    SB_LUT4 i31283_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n45363));
    defparam i31283_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(delay_counter[22]), .I1(delay_counter[21]), 
            .I2(n25774), .I3(delay_counter[23]), .O(n4_adj_5747));
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1829 (.I0(n68999), .I1(delay_counter[18]), .I2(n25771), 
            .I3(GND_net), .O(n68987));
    defparam i2_3_lut_adj_1829.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n58904), .I0(n2533), 
            .I1(VCC_net), .CO(n58905));
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n58492), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n58904));
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n58492), .I0(n1325), 
            .I1(VCC_net), .CO(n58493));
    SB_LUT4 i2_4_lut_adj_1830 (.I0(n68987), .I1(n4_adj_5747), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n62));
    defparam i2_4_lut_adj_1830.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n58491), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n59414), .O(n38_adj_5936)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2038_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n59413), .O(n39_adj_5937)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n58491), .I0(n1326), 
            .I1(VCC_net), .CO(n58492));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n58490), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n58490), .I0(n1327), 
            .I1(VCC_net), .CO(n58491));
    SB_LUT4 i56072_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71907));
    defparam i56072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16501_3_lut (.I0(ID[7]), .I1(data_adj_6032[7]), .I2(n68385), 
            .I3(GND_net), .O(n30713));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16502_3_lut (.I0(ID[6]), .I1(data_adj_6032[6]), .I2(n68385), 
            .I3(GND_net), .O(n30714));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16502_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i56073_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71908));
    defparam i56073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55920_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71755));
    defparam i55920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55919_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71754));
    defparam i55919_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2038_add_4_8 (.CI(n59413), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n59414));
    SB_LUT4 dti_counter_2038_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n59412), .O(n40_adj_5938)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_7 (.CI(n59412), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n59413));
    SB_LUT4 dti_counter_2038_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n59411), .O(n41_adj_5939)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_6 (.CI(n59411), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n59412));
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30588_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(366[12:35])
    defparam i30588_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 dti_counter_2038_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n59410), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n58489), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_5 (.CI(n59410), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n59411));
    SB_LUT4 dti_counter_2038_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n59409), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_4 (.CI(n59409), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n59410));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n58295), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n58489), .I0(n1328), 
            .I1(VCC_net), .CO(n58490));
    SB_LUT4 i16503_3_lut (.I0(ID[5]), .I1(data_adj_6032[5]), .I2(n68385), 
            .I3(GND_net), .O(n30715));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16503_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut (.I0(n11849), .I1(current[15]), .I2(duty[15]), 
            .I3(n11847), .O(n79029));
    defparam n11849_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 dti_counter_2038_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n59408), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_3 (.CI(n59408), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n59409));
    SB_LUT4 i16504_3_lut (.I0(ID[4]), .I1(data_adj_6032[4]), .I2(n68385), 
            .I3(GND_net), .O(n30716));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2038_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n58488), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16505_3_lut (.I0(ID[3]), .I1(data_adj_6032[3]), .I2(n68385), 
            .I3(GND_net), .O(n30717));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16505_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2038_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n59408));
    SB_LUT4 n79029_bdd_4_lut (.I0(n79029), .I1(duty[12]), .I2(n4916), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[12]));
    defparam n79029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1831 (.I0(n37336), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_1831.LUT_INIT = 16'h8888;
    SB_LUT4 i16506_3_lut (.I0(ID[2]), .I1(data_adj_6032[2]), .I2(n68385), 
            .I3(GND_net), .O(n30718));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16506_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n58488), .I0(n1329), 
            .I1(GND_net), .CO(n58489));
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n58487), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16507_3_lut (.I0(ID[1]), .I1(data_adj_6032[1]), .I2(n68385), 
            .I3(GND_net), .O(n30719));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16507_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n58487), .I0(n1330), 
            .I1(GND_net), .CO(n58488));
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n58486), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n58486), .I0(n1331), 
            .I1(VCC_net), .CO(n58487));
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [7]), .O(n66680));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n58295), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n58296));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n58294), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n58294), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n58295));
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n44439), .O(n64350));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hb1f1;
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n58485), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n58485), .I0(n1332), 
            .I1(GND_net), .CO(n58486));
    SB_LUT4 i1_2_lut_adj_1832 (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_5845), 
            .I2(GND_net), .I3(GND_net), .O(n85));
    defparam i1_2_lut_adj_1832.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n58484), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n58484), .I0(n1333), 
            .I1(VCC_net), .CO(n58485));
    SB_LUT4 n11849_bdd_4_lut_63098 (.I0(n11849), .I1(current[11]), .I2(duty[14]), 
            .I3(n11847), .O(n79023));
    defparam n11849_bdd_4_lut_63098.LUT_INIT = 16'he4aa;
    SB_LUT4 n79023_bdd_4_lut (.I0(n79023), .I1(duty[11]), .I2(n4917), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[11]));
    defparam n79023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5859), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63093 (.I0(n11849), .I1(current[10]), .I2(duty[13]), 
            .I3(n11847), .O(n79017));
    defparam n11849_bdd_4_lut_63093.LUT_INIT = 16'he4aa;
    SB_LUT4 i16520_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n23023), .I3(GND_net), .O(n30732));   // verilog/coms.v(130[12] 305[6])
    defparam i16520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1833 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n70001));
    defparam i1_3_lut_adj_1833.LUT_INIT = 16'hfefe;
    SB_LUT4 i61844_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77679));
    defparam i61844_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n58293), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62195_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78030));
    defparam i62195_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1834 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n70281));
    defparam i1_2_lut_adj_1834.LUT_INIT = 16'h8888;
    SB_LUT4 i62417_4_lut (.I0(n70281), .I1(n1125), .I2(n70001), .I3(n45363), 
            .O(n1158));
    defparam i62417_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n79017_bdd_4_lut (.I0(n79017), .I1(duty[10]), .I2(n4918), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[10]));
    defparam n79017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n58484));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n58293), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n58294));
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(n78264), .I1(n1224_adj_5848), 
            .I2(VCC_net), .I3(n58483), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5849), 
            .I2(VCC_net), .I3(n58482), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n58482), .I0(n1225_adj_5849), 
            .I1(VCC_net), .CO(n58483));
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5850), 
            .I2(VCC_net), .I3(n58481), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62485_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78320));
    defparam i62485_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31205_3_lut (.I0(n937), .I1(n1232_adj_5856), .I2(n1233_adj_5857), 
            .I3(GND_net), .O(n45285));
    defparam i31205_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1835 (.I0(n1226_adj_5850), .I1(n1227_adj_5851), 
            .I2(n1228_adj_5852), .I3(GND_net), .O(n70343));
    defparam i1_3_lut_adj_1835.LUT_INIT = 16'hfefe;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n28128), 
            .D(n1229), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n28128), 
            .D(n1228), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i61901_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77736));
    defparam i61901_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n1229_adj_5853), .I1(n45285), .I2(n1230_adj_5854), 
            .I3(n1231_adj_5855), .O(n67722));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'ha080;
    SB_LUT4 i62432_4_lut (.I0(n1225_adj_5849), .I1(n1224_adj_5848), .I2(n67722), 
            .I3(n70343), .O(n1257));
    defparam i62432_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5854));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6653_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6653_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i31201_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n45281));
    defparam i31201_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n70265));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(n1329), .I1(n45281), .I2(n1330), .I3(n1331), 
            .O(n67720));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'ha080;
    SB_LUT4 mux_1677_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n11912));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62448_4_lut (.I0(n67720), .I1(n1323), .I2(n1324), .I3(n70265), 
            .O(n1356));
    defparam i62448_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5854), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31211_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n45291));
    defparam i31211_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1839 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n70329));
    defparam i1_2_lut_adj_1839.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n1429), .I1(n45291), .I2(n1430), .I3(n1431), 
            .O(n67733));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n70329), 
            .O(n70335));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1677_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12490));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62465_4_lut (.I0(n1423), .I1(n1422), .I2(n70335), .I3(n67733), 
            .O(n1455));
    defparam i62465_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31213_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n45293));
    defparam i31213_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1842 (.I0(n1525), .I1(n1528), .I2(n1527), .I3(GND_net), 
            .O(n70321));
    defparam i1_3_lut_adj_1842.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1843 (.I0(n1529), .I1(n70321), .I2(n45293), .I3(n1530), 
            .O(n70323));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'heccc;
    SB_LUT4 i1_3_lut_adj_1844 (.I0(n1522), .I1(n1524), .I2(n1526), .I3(GND_net), 
            .O(n70257));
    defparam i1_3_lut_adj_1844.LUT_INIT = 16'hfefe;
    SB_LUT4 i62393_4_lut (.I0(n70257), .I1(n1521), .I2(n70323), .I3(n1523), 
            .O(n1554));
    defparam i62393_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31215_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n45295));
    defparam i31215_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1845 (.I0(\data_in_frame[18] [7]), .I1(n28654), 
            .I2(n28711), .I3(rx_data[7]), .O(n65160));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1845.LUT_INIT = 16'h3a0a;
    SB_LUT4 i16526_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n28711), .I3(GND_net), .O(n30738));   // verilog/coms.v(130[12] 305[6])
    defparam i16526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15520_3_lut (.I0(\data_in_frame[18] [6]), .I1(rx_data[6]), 
            .I2(n28711), .I3(GND_net), .O(n29732));   // verilog/coms.v(130[12] 305[6])
    defparam i15520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1677_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12488));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15517_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n28711), .I3(GND_net), .O(n29729));   // verilog/coms.v(130[12] 305[6])
    defparam i15517_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i6_4_lut_adj_1846 (.I0(ID[5]), .I1(ID[4]), .I2(ID[2]), .I3(ID[6]), 
            .O(n14_adj_5961));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i6_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n28128), 
            .D(n1227), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 mux_1677_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n12486));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i4_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n58481), .I0(n1226_adj_5850), 
            .I1(VCC_net), .CO(n58482));
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n70361));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n1629), .I1(n45295), .I2(n1630), .I3(n1631), 
            .O(n67741));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1849 (.I0(ID[0]), .I1(ID[1]), .I2(ID[7]), .I3(ID[3]), 
            .O(n13_adj_5962));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i5_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i30365_4_lut (.I0(n13_adj_5962), .I1(n33), .I2(n14_adj_5961), 
            .I3(n34), .O(n44439));
    defparam i30365_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i12_4_lut_adj_1850 (.I0(\data_in_frame[18] [4]), .I1(n28654), 
            .I2(n28711), .I3(rx_data[4]), .O(n65164));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1850.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_1677_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12484));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i5_3_lut.LUT_INIT = 16'h3535;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1851 (.I0(n1623), .I1(n67741), .I2(n1624), .I3(n70361), 
            .O(n70367));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62213_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n70367), 
            .O(n1653));
    defparam i62213_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1852 (.I0(n1725), .I1(n1728), .I2(n1727), .I3(n1726), 
            .O(n70207));
    defparam i1_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i31217_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n45297));
    defparam i31217_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1853 (.I0(n1723), .I1(n1724), .I2(n70207), .I3(GND_net), 
            .O(n70211));
    defparam i1_3_lut_adj_1853.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1854 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n70373));
    defparam i1_2_lut_adj_1854.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1677_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12482));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12480));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12478));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12476));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i61941_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77776));
    defparam i61941_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12474));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12472));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16534_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n21152), .I3(n4_adj_5971), .O(n30746));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16534_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 mux_1677_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12470));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12468));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i59097_3_lut (.I0(state_7__N_4110[0]), .I1(n11_adj_5794), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n74657));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i59097_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 mux_1677_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12466));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12464));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12462));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12460));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12458));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12456));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16_4_lut (.I0(state_adj_6068[0]), .I1(n74657), .I2(n6705), 
            .I3(n44499), .O(n8_adj_5974));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut.LUT_INIT = 16'h3afa;
    SB_LUT4 i62535_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78370));
    defparam i62535_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12454));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14964_4_lut (.I0(n28128), .I1(n1319), .I2(n74462), .I3(n44534), 
            .O(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i14964_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16537_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[0]), 
            .I2(n10_adj_5953), .I3(n25888), .O(n30749));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16537_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i62105_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77940));
    defparam i62105_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1677_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12452));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i61989_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77824));
    defparam i61989_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29445_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[11]));
    defparam i29445_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_4_lut_adj_1855 (.I0(\data_in_frame[18] [3]), .I1(n28654), 
            .I2(n28711), .I3(rx_data[3]), .O(n65168));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1855.LUT_INIT = 16'h3a0a;
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n69276));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n66892));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16544_3_lut (.I0(n67079), .I1(r_Bit_Index[0]), .I2(n28238), 
            .I3(GND_net), .O(n30756));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16544_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 mux_1677_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12450));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i62043_1_lut (.I0(n45345), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77878));
    defparam i62043_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5944));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5943));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5946));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5941));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5860), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33_adj_5947));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n3228), .I1(n29_adj_5946), .I2(n3295), 
            .I3(n3237), .O(n70005));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5942));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n19_adj_5942), .I1(n70005), .I2(n33_adj_5947), 
            .I3(n13_adj_5941), .O(n70011));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n3217), .I1(n70011), .I2(n3284), .I3(n3237), 
            .O(n70013));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6651_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6651_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n3216), .I1(n70013), .I2(n3283), .I3(n3237), 
            .O(n70015));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n3215), .I1(n70015), .I2(n3282), .I3(n3237), 
            .O(n70017));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n3213), .I1(n70017), .I2(n3280), .I3(n3237), 
            .O(n70019));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n3212), .I1(n70019), .I2(n3279), .I3(n3237), 
            .O(n70021));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(n3211), .I1(n70021), .I2(n3278), .I3(n3237), 
            .O(n70023));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'heefc;
    SB_LUT4 n11849_bdd_4_lut_63088 (.I0(n11849), .I1(current[9]), .I2(duty[12]), 
            .I3(n11847), .O(n78999));
    defparam n11849_bdd_4_lut_63088.LUT_INIT = 16'he4aa;
    SB_LUT4 n78999_bdd_4_lut (.I0(n78999), .I1(duty[9]), .I2(n4919), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n78999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(n3210), .I1(n70023), .I2(n3277), .I3(n3237), 
            .O(n70025));
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1865 (.I0(n3209), .I1(n70025), .I2(n3276), .I3(n3237), 
            .O(n70027));
    defparam i1_4_lut_adj_1865.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5945));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1866 (.I0(n3231), .I1(n74442), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5922));
    defparam i16_4_lut_adj_1866.LUT_INIT = 16'hac0c;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59254_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n74589));
    defparam i59254_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(n3222), .I1(n23_adj_5944), .I2(n3289), 
            .I3(n3237), .O(n70303));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n3220), .I1(n21_adj_5943), .I2(n3287), 
            .I3(n3237), .O(n70301));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1869 (.I0(n74589), .I1(n5_adj_5922), .I2(n74590), 
            .I3(n3237), .O(n62242));
    defparam i1_4_lut_adj_1869.LUT_INIT = 16'h88c0;
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1870 (.I0(n3227), .I1(n25_adj_5945), .I2(n3294), 
            .I3(n3237), .O(n70305));
    defparam i1_4_lut_adj_1870.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1871 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69681), .O(n69687));
    defparam i1_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1872 (.I0(n70305), .I1(n62242), .I2(n70301), 
            .I3(n70303), .O(n70311));
    defparam i1_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1873 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69687), .O(n69693));
    defparam i1_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1874 (.I0(n70373), .I1(n1722), .I2(n70211), .I3(n45297), 
            .O(n70215));
    defparam i1_4_lut_adj_1874.LUT_INIT = 16'hfefc;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62504_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n70215), 
            .O(n1752));
    defparam i62504_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1875 (.I0(n1825), .I1(n1826), .I2(n1827), .I3(n1828), 
            .O(n70381));
    defparam i1_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i31219_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n45299));
    defparam i31219_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1876 (.I0(n1823), .I1(n1824), .I2(n70381), .I3(GND_net), 
            .O(n70385));
    defparam i1_3_lut_adj_1876.LUT_INIT = 16'hfefe;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1877 (.I0(n1829), .I1(n45299), .I2(n1830), .I3(n1831), 
            .O(n67779));
    defparam i1_4_lut_adj_1877.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1878 (.I0(n1821), .I1(n1822), .I2(n67779), .I3(n70385), 
            .O(n70391));
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i62555_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n70391), 
            .O(n1851));
    defparam i62555_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5861), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_adj_1879 (.I0(n1926), .I1(n1925), .I2(GND_net), .I3(GND_net), 
            .O(n70075));
    defparam i1_2_lut_adj_1879.LUT_INIT = 16'heeee;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1880 (.I0(n70311), .I1(n3218), .I2(n3285), .I3(n3237), 
            .O(n70313));
    defparam i1_4_lut_adj_1880.LUT_INIT = 16'heefa;
    SB_LUT4 i16548_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n69693), 
            .I3(n27_adj_5865), .O(n30760));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16548_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1881 (.I0(n3214), .I1(n70313), .I2(n3281), .I3(n3237), 
            .O(n70315));
    defparam i1_4_lut_adj_1881.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1882 (.I0(n3207), .I1(n70315), .I2(n3274), .I3(n3237), 
            .O(n70317));
    defparam i1_4_lut_adj_1882.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1883 (.I0(n3208), .I1(n70027), .I2(n3275), .I3(n3237), 
            .O(n70029));
    defparam i1_4_lut_adj_1883.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n28128), 
            .D(n1226), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n28128), 
            .D(n1225), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_4_lut_adj_1884 (.I0(n70317), .I1(n3206), .I2(n3273), .I3(n3237), 
            .O(n68824));
    defparam i1_4_lut_adj_1884.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61_adj_5948));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62046_4_lut (.I0(n61_adj_5948), .I1(n71361), .I2(n68824), 
            .I3(n70029), .O(n45345));
    defparam i62046_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12448));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16549_3_lut (.I0(\data_in_frame[0] [0]), .I1(rx_data[0]), .I2(n7_adj_5975), 
            .I3(GND_net), .O(n30761));   // verilog/coms.v(130[12] 305[6])
    defparam i16549_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n28128), 
            .D(n1224), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i16553_4_lut (.I0(CS_MISO_c), .I1(data_adj_6039[0]), .I2(n11_adj_5799), 
            .I3(state_7__N_4319), .O(n30765));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16553_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5851), 
            .I2(VCC_net), .I3(n58480), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n28128), 
            .D(n1223), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n28128), 
            .D(n1222), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n28128), 
            .D(n1221), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n28128), 
            .D(n1220), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n28128), 
            .D(n1219), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_3_lut_adj_1885 (.I0(n1928), .I1(n1924), .I2(n1927), .I3(GND_net), 
            .O(n70077));
    defparam i1_3_lut_adj_1885.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n58480), .I0(n1227_adj_5851), 
            .I1(VCC_net), .CO(n58481));
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n28128), 
            .D(n1218), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n28128), 
            .D(n1217), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n28128), 
            .D(n1216), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n28128), 
            .D(n1215), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n28128), 
            .D(n1214), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n28128), 
            .D(n1213), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n28128), 
            .D(n1212), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n28128), 
            .D(n1211), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n28128), 
            .D(n1210), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n28128), 
            .D(n1209), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n28128), 
            .D(n1208), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR dti_counter_2038__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n28172), 
            .D(n44), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n28172), 
            .D(n43), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n28172), 
            .D(n42), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n28172), 
            .D(n41_adj_5939), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n28172), 
            .D(n40_adj_5938), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n28172), 
            .D(n39_adj_5937), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n28172), 
            .D(n38_adj_5936), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6655_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6655_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i12_4_lut_adj_1886 (.I0(\data_in_frame[18] [2]), .I1(n28654), 
            .I2(n28711), .I3(rx_data[2]), .O(n65172));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1886.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5734), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63073 (.I0(n11849), .I1(current[8]), .I2(duty[11]), 
            .I3(n11847), .O(n78993));
    defparam n11849_bdd_4_lut_63073.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n78993_bdd_4_lut (.I0(n78993), .I1(duty[8]), .I2(n4920), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n78993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1887 (.I0(n3223), .I1(n3225), .I2(GND_net), .I3(GND_net), 
            .O(n70663));
    defparam i1_2_lut_adj_1887.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1888 (.I0(n3221), .I1(n3218), .I2(n3228), .I3(n3224), 
            .O(n70675));
    defparam i1_4_lut_adj_1888.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1889 (.I0(n3217), .I1(n3227), .I2(n3222), .I3(n3226), 
            .O(n70679));
    defparam i1_4_lut_adj_1889.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1890 (.I0(n3219), .I1(n70675), .I2(n70663), .I3(n3220), 
            .O(n70681));
    defparam i1_4_lut_adj_1890.LUT_INIT = 16'hfffe;
    SB_LUT4 i31156_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n45233));
    defparam i31156_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5852), 
            .I2(VCC_net), .I3(n58479), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n58479), .I0(n1228_adj_5852), 
            .I1(VCC_net), .CO(n58480));
    SB_LUT4 i1_4_lut_adj_1891 (.I0(n3215), .I1(n70681), .I2(n3216), .I3(n70679), 
            .O(n70687));
    defparam i1_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1892 (.I0(n3229), .I1(n45233), .I2(n3230), .I3(n3231), 
            .O(n67871));
    defparam i1_4_lut_adj_1892.LUT_INIT = 16'ha080;
    SB_LUT4 n11849_bdd_4_lut_63068 (.I0(n11849), .I1(current[7]), .I2(duty[10]), 
            .I3(n11847), .O(n78981));
    defparam n11849_bdd_4_lut_63068.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1893 (.I0(n3213), .I1(n3214), .I2(n67871), .I3(n70687), 
            .O(n70693));
    defparam i1_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 n78981_bdd_4_lut (.I0(n78981), .I1(duty[7]), .I2(n4921), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n78981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1894 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n70693), 
            .O(n70699));
    defparam i1_4_lut_adj_1894.LUT_INIT = 16'hfffe;
    SB_LUT4 i31138_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n45215));
    defparam i31138_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5853), 
            .I2(GND_net), .I3(n58478), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n58478), .I0(n1229_adj_5853), 
            .I1(GND_net), .CO(n58479));
    SB_LUT4 i1_4_lut_adj_1895 (.I0(n1922), .I1(n1923), .I2(n70077), .I3(n70075), 
            .O(n70083));
    defparam i1_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1896 (.I0(n1929), .I1(n45215), .I2(n1930), .I3(n1931), 
            .O(n67763));
    defparam i1_4_lut_adj_1896.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1897 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n70699), 
            .O(n70705));
    defparam i1_4_lut_adj_1897.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(n1920), .I1(n67763), .I2(n1921), .I3(n70083), 
            .O(n70089));
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62042_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n70089), 
            .O(n1950));
    defparam i62042_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i62020_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n70705), 
            .O(n3237));
    defparam i62020_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31235_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n45315));
    defparam i31235_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1899 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n70427));
    defparam i1_2_lut_adj_1899.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(n2025), .I1(n70427), .I2(n2024), .I3(n2028), 
            .O(n70431));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(n2029), .I1(n45315), .I2(n2030), .I3(n2031), 
            .O(n67800));
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'ha080;
    SB_DFFESR dti_counter_2038__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n28172), 
            .D(n45), .R(n29436));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5854), 
            .I2(GND_net), .I3(n58477), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1902 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n70431), 
            .O(n70437));
    defparam i1_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n58477), .I0(n1230_adj_5854), 
            .I1(GND_net), .CO(n58478));
    SB_LUT4 i15825_3_lut_4_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30037));   // verilog/coms.v(130[12] 305[6])
    defparam i15825_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n11849_bdd_4_lut_63058 (.I0(n11849), .I1(current[6]), .I2(duty[9]), 
            .I3(n11847), .O(n78969));
    defparam n11849_bdd_4_lut_63058.LUT_INIT = 16'he4aa;
    SB_LUT4 n78969_bdd_4_lut (.I0(n78969), .I1(duty[6]), .I2(n4922), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n78969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1903 (.I0(n2019), .I1(n2020), .I2(n70437), .I3(n67800), 
            .O(n70443));
    defparam i1_4_lut_adj_1903.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62296_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n70443), 
            .O(n2049));
    defparam i62296_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1904 (.I0(n2125), .I1(n2127), .I2(GND_net), .I3(GND_net), 
            .O(n70221));
    defparam i1_2_lut_adj_1904.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31303_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n45383));
    defparam i31303_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63048 (.I0(n11849), .I1(current[5]), .I2(duty[8]), 
            .I3(n11847), .O(n78963));
    defparam n11849_bdd_4_lut_63048.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1905 (.I0(n2122), .I1(n2126), .I2(n70221), .I3(n2128), 
            .O(n70227));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1906 (.I0(n2129), .I1(n70227), .I2(n45383), .I3(n2130), 
            .O(n70229));
    defparam i1_4_lut_adj_1906.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15824_3_lut_4_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30036));   // verilog/coms.v(130[12] 305[6])
    defparam i15824_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_1907 (.I0(n2118), .I1(n2119), .I2(n70229), .I3(n2120), 
            .O(n70235));
    defparam i1_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5855), 
            .I2(VCC_net), .I3(n58476), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1908 (.I0(n2121), .I1(n2117), .I2(n2123), .I3(n2124), 
            .O(n68961));
    defparam i1_4_lut_adj_1908.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62320_4_lut (.I0(n68961), .I1(n2115), .I2(n2116), .I3(n70235), 
            .O(n2148));
    defparam i62320_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3812_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5738), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n58476), .I0(n1231_adj_5855), 
            .I1(VCC_net), .CO(n58477));
    SB_LUT4 i31233_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n45313));
    defparam i31233_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 n78963_bdd_4_lut (.I0(n78963), .I1(duty[5]), .I2(n4923), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n78963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6657_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6657_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1909 (.I0(n2224), .I1(n2225), .I2(n2226), .I3(n2227), 
            .O(n70407));
    defparam i1_4_lut_adj_1909.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1910 (.I0(n2229), .I1(n45313), .I2(n2230), .I3(n2231), 
            .O(n67807));
    defparam i1_4_lut_adj_1910.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1911 (.I0(n2221), .I1(n2220), .I2(n2223), .I3(n2228), 
            .O(n68995));
    defparam i1_4_lut_adj_1911.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(n68995), .I1(n67807), .I2(n2222), .I3(n70407), 
            .O(n70413));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1913 (.I0(n2217), .I1(n2218), .I2(n70413), .I3(n2219), 
            .O(n70419));
    defparam i1_4_lut_adj_1913.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62273_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n70419), 
            .O(n2247));
    defparam i62273_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5856), 
            .I2(GND_net), .I3(n58475), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31229_3_lut (.I0(n948), .I1(n2332), .I2(n2333), .I3(GND_net), 
            .O(n45309));
    defparam i31229_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1914 (.I0(n2321), .I1(n2322), .I2(n2324), .I3(GND_net), 
            .O(n70243));
    defparam i1_3_lut_adj_1914.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63043 (.I0(n11849), .I1(current[4]), .I2(duty[7]), 
            .I3(n11847), .O(n78957));
    defparam n11849_bdd_4_lut_63043.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1915 (.I0(n2326), .I1(n2325), .I2(n2328), .I3(GND_net), 
            .O(n70291));
    defparam i1_3_lut_adj_1915.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n58475), .I0(n1232_adj_5856), 
            .I1(GND_net), .CO(n58476));
    SB_LUT4 i1_2_lut_adj_1916 (.I0(n8_adj_5846), .I1(n41543), .I2(GND_net), 
            .I3(GND_net), .O(n28654));
    defparam i1_2_lut_adj_1916.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5857), 
            .I2(VCC_net), .I3(n58474), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n58474), .I0(n1233_adj_5857), 
            .I1(VCC_net), .CO(n58475));
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n58474));
    SB_LUT4 i12_4_lut_adj_1917 (.I0(\data_in_frame[18] [1]), .I1(n28654), 
            .I2(n28711), .I3(rx_data[1]), .O(n65176));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1917.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n78239), .I1(n1125), 
            .I2(VCC_net), .I3(n58473), .O(n1224_adj_5848)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n58472), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31247_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n45327));
    defparam i31247_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1918 (.I0(n3125), .I1(n3123), .I2(n3122), .I3(n3127), 
            .O(n70135));
    defparam i1_4_lut_adj_1918.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1919 (.I0(n3124), .I1(n3128), .I2(n3121), .I3(n3120), 
            .O(n70137));
    defparam i1_4_lut_adj_1919.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1920 (.I0(n70137), .I1(n70135), .I2(n3119), .I3(n3126), 
            .O(n70141));
    defparam i1_4_lut_adj_1920.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1921 (.I0(n3129), .I1(n45327), .I2(n3130), .I3(n3131), 
            .O(n67825));
    defparam i1_4_lut_adj_1921.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n58472), .I0(n1126), 
            .I1(VCC_net), .CO(n58473));
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n58471), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1922 (.I0(n3116), .I1(n3117), .I2(n70141), .I3(n3118), 
            .O(n70147));
    defparam i1_4_lut_adj_1922.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1923 (.I0(n3114), .I1(n3115), .I2(n70147), .I3(n67825), 
            .O(n70153));
    defparam i1_4_lut_adj_1923.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1924 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n70153), 
            .O(n70159));
    defparam i1_4_lut_adj_1924.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1925 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n70159), 
            .O(n70165));
    defparam i1_4_lut_adj_1925.LUT_INIT = 16'hfffe;
    SB_LUT4 i61974_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n70165), 
            .O(n3138));
    defparam i61974_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15822_3_lut_4_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30034));   // verilog/coms.v(130[12] 305[6])
    defparam i15822_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15821_3_lut_4_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30033));   // verilog/coms.v(130[12] 305[6])
    defparam i15821_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n58471), .I0(n1127), 
            .I1(VCC_net), .CO(n58472));
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n58470), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15820_3_lut_4_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30032));   // verilog/coms.v(130[12] 305[6])
    defparam i15820_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15819_3_lut_4_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30031));   // verilog/coms.v(130[12] 305[6])
    defparam i15819_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15818_3_lut_4_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30030));   // verilog/coms.v(130[12] 305[6])
    defparam i15818_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n58470), .I0(n1128), 
            .I1(VCC_net), .CO(n58471));
    SB_LUT4 i59638_4_lut (.I0(data_ready), .I1(n6901), .I2(n24_adj_5957), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n74606));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i59638_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59594_2_lut (.I0(n24_adj_5957), .I1(n6901), .I2(GND_net), 
            .I3(GND_net), .O(n74609));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i59594_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n74609), .I1(n74606), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5963), .O(n64260));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n58469), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n78957_bdd_4_lut (.I0(n78957), .I1(duty[4]), .I2(n4924), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n78957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n64260));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i1_4_lut_adj_1926 (.I0(n3027), .I1(n3022), .I2(n3026), .I3(n3019), 
            .O(n70589));
    defparam i1_4_lut_adj_1926.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1927 (.I0(n3021), .I1(n3020), .I2(n3024), .I3(n3023), 
            .O(n70587));
    defparam i1_4_lut_adj_1927.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1928 (.I0(n70589), .I1(n3028), .I2(n3018), .I3(n3025), 
            .O(n70591));
    defparam i1_4_lut_adj_1928.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n77940), .I1(n2412), 
            .I2(VCC_net), .I3(n58872), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n58469), .I0(n1129), 
            .I1(GND_net), .CO(n58470));
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30746));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n58468), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n58871), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n58468), .I0(n1130), 
            .I1(GND_net), .CO(n58469));
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n58467), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31309_4_lut (.I0(n955), .I1(n3031), .I2(n3032), .I3(n3033), 
            .O(n45389));
    defparam i31309_4_lut.LUT_INIT = 16'hfcec;
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n58871), .I0(n2413), 
            .I1(VCC_net), .CO(n58872));
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n58467), .I0(n1131), 
            .I1(VCC_net), .CO(n58468));
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n58466), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n58870), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n58466), .I0(n1132), 
            .I1(GND_net), .CO(n58467));
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n58465), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1929 (.I0(n3016), .I1(n70591), .I2(n3017), .I3(n70587), 
            .O(n70597));
    defparam i1_4_lut_adj_1929.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n58870), .I0(n2414), 
            .I1(VCC_net), .CO(n58871));
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n58465), .I0(n1133), 
            .I1(VCC_net), .CO(n58466));
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n58869), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n58465));
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n58464), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1930 (.I0(n3029), .I1(n3030), .I2(GND_net), .I3(GND_net), 
            .O(n70721));
    defparam i1_2_lut_adj_1930.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1931 (.I0(n3015), .I1(n70721), .I2(n70597), .I3(n45389), 
            .O(n70601));
    defparam i1_4_lut_adj_1931.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1932 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n70601), 
            .O(n70607));
    defparam i1_4_lut_adj_1932.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1933 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n70607), 
            .O(n70613));
    defparam i1_4_lut_adj_1933.LUT_INIT = 16'hfffe;
    SB_LUT4 i61933_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n70613), 
            .O(n3039));
    defparam i61933_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1907_3_lut (.I0(n2808), .I1(n2875), 
            .I2(n2841), .I3(GND_net), .O(n2907));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15817_3_lut_4_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30029));   // verilog/coms.v(130[12] 305[6])
    defparam i15817_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n58869), .I0(n2415), 
            .I1(VCC_net), .CO(n58870));
    SB_LUT4 i51122_3_lut (.I0(n6_adj_5749), .I1(n7758), .I2(n66893), .I3(GND_net), 
            .O(n66900));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51123_3_lut (.I0(encoder0_position[26]), .I1(n66900), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n58463), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5852));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n58463), .I0(n1027), 
            .I1(VCC_net), .CO(n58464));
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n58868), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n58462), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n58462), .I0(n1028), 
            .I1(VCC_net), .CO(n58463));
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n58868), .I0(n2416), 
            .I1(VCC_net), .CO(n58869));
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n58461), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5852), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819_adj_5867), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n58867), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n58867), .I0(n2417), 
            .I1(VCC_net), .CO(n58868));
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62404_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78239));
    defparam i62404_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n58461), .I0(n1029), 
            .I1(GND_net), .CO(n58462));
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n58866), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n58460), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n58460), .I0(n1030), 
            .I1(GND_net), .CO(n58461));
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n58459), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62505_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78340));
    defparam i62505_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n58866), .I0(n2418), 
            .I1(VCC_net), .CO(n58867));
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n58459), .I0(n1031), 
            .I1(VCC_net), .CO(n58460));
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n58458), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n58865), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n58458), .I0(n1032), 
            .I1(GND_net), .CO(n58459));
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n58457), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n58865), .I0(n2419), 
            .I1(VCC_net), .CO(n58866));
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n58457), .I0(n1033), 
            .I1(VCC_net), .CO(n58458));
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n58864), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n58457));
    SB_LUT4 i31243_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n45323));
    defparam i31243_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n58456), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1934 (.I0(n2928), .I1(n2923), .I2(n2921), .I3(n2927), 
            .O(n70101));
    defparam i1_4_lut_adj_1934.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1935 (.I0(n2922), .I1(n2920), .I2(n2926), .I3(GND_net), 
            .O(n70555));
    defparam i1_3_lut_adj_1935.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1936 (.I0(n2929), .I1(n45323), .I2(n2930), .I3(n2931), 
            .O(n67816));
    defparam i1_4_lut_adj_1936.LUT_INIT = 16'ha080;
    SB_LUT4 i15816_3_lut_4_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30028));   // verilog/coms.v(130[12] 305[6])
    defparam i15816_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_3_lut_adj_1937 (.I0(n70101), .I1(n2924), .I2(n2925), .I3(GND_net), 
            .O(n70103));
    defparam i1_3_lut_adj_1937.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1938 (.I0(n2917), .I1(n2918), .I2(n2919), .I3(n70555), 
            .O(n70561));
    defparam i1_4_lut_adj_1938.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1939 (.I0(n2916), .I1(n70561), .I2(n70103), .I3(n67816), 
            .O(n70107));
    defparam i1_4_lut_adj_1939.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1940 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n70107), 
            .O(n70113));
    defparam i1_4_lut_adj_1940.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1941 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n70113), 
            .O(n70119));
    defparam i1_4_lut_adj_1941.LUT_INIT = 16'hfffe;
    SB_LUT4 i61875_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n70119), 
            .O(n2940));
    defparam i61875_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i62583_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78418));
    defparam i62583_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62188_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78023));
    defparam i62188_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n58864), .I0(n2420), 
            .I1(VCC_net), .CO(n58865));
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n58455), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62236_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78071));
    defparam i62236_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n58455), .I0(n928), 
            .I1(VCC_net), .CO(n58456));
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n58863), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n58454), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62270_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78105));
    defparam i62270_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n58454), .I0(n929), 
            .I1(GND_net), .CO(n58455));
    SB_LUT4 i62293_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78128));
    defparam i62293_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n58863), .I0(n2421), 
            .I1(VCC_net), .CO(n58864));
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n58453), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n58453), .I0(n930), 
            .I1(GND_net), .CO(n58454));
    SB_LUT4 i62039_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n77874));
    defparam i62039_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n58862), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n58452), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n58452), .I0(n931), 
            .I1(VCC_net), .CO(n58453));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5830));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n58862), .I0(n2422), 
            .I1(VCC_net), .CO(n58863));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n58451), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n58451), .I0(n932), 
            .I1(GND_net), .CO(n58452));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n58861), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62390_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78225));
    defparam i62390_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n58450), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62429_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78264));
    defparam i62429_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51120_3_lut (.I0(n5), .I1(n7757), .I2(n66893), .I3(GND_net), 
            .O(n66898));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51120_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n58450), .I0(n933), 
            .I1(VCC_net), .CO(n58451));
    SB_LUT4 i51121_3_lut (.I0(encoder0_position[27]), .I1(n66898), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51121_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n58861), .I0(n2423), 
            .I1(VCC_net), .CO(n58862));
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n58450));
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n58860), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n58449), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n58448), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i62475_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n78310));
    defparam i62475_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5917));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n58448), .I0(n829), 
            .I1(GND_net), .CO(n58449));
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5916));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5915));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n58860), .I0(n2424), 
            .I1(VCC_net), .CO(n58861));
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n58859), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n58859), .I0(n2425), 
            .I1(VCC_net), .CO(n58860));
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n58447), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n58447), .I0(n830), 
            .I1(GND_net), .CO(n58448));
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n58858), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n58292), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n58858), .I0(n2426), 
            .I1(VCC_net), .CO(n58859));
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n58446), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n58857), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n58292), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n58293));
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n58857), .I0(n2427), 
            .I1(VCC_net), .CO(n58858));
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n58856), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n58856), .I0(n2428), 
            .I1(VCC_net), .CO(n58857));
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n58855), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5914));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5913));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5912));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5911));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n58446), .I0(n831), 
            .I1(VCC_net), .CO(n58447));
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1942 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66166));
    defparam i1_2_lut_adj_1942.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n58855), .I0(n2429), 
            .I1(GND_net), .CO(n58856));
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n58854), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n58445), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n58445), .I0(n832), 
            .I1(GND_net), .CO(n58446));
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n58854), .I0(n2430), 
            .I1(GND_net), .CO(n58855));
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n58444), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n58444), .I0(n833), 
            .I1(VCC_net), .CO(n58445));
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5851));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n58853), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n58444));
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n58853), .I0(n2431), 
            .I1(VCC_net), .CO(n58854));
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5851), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n58852), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2584_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n58443), 
            .O(n7754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2584_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n58442), 
            .O(n7755)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n58852), .I0(n2432), 
            .I1(GND_net), .CO(n58853));
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n58851), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_6 (.CI(n58442), .I0(n622), .I1(GND_net), .CO(n58443));
    SB_LUT4 add_2584_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n58441), 
            .O(n7756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n58851), .I0(n2433), 
            .I1(VCC_net), .CO(n58852));
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n58851));
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15815_3_lut_4_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30027));   // verilog/coms.v(130[12] 305[6])
    defparam i15815_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_2584_5 (.CI(n58441), .I0(n623), .I1(VCC_net), .CO(n58442));
    SB_LUT4 add_2584_4_lut (.I0(GND_net), .I1(n291_adj_5812), .I2(GND_net), 
            .I3(n58440), .O(n7757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_4 (.CI(n58440), .I0(n291_adj_5812), .I1(GND_net), 
            .CO(n58441));
    SB_LUT4 add_2584_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n58439), 
            .O(n7758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_3 (.CI(n58439), .I0(n625), .I1(VCC_net), .CO(n58440));
    SB_LUT4 add_2584_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2584_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2584_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n58439));
    SB_LUT4 n11849_bdd_4_lut_63038 (.I0(n11849), .I1(current[3]), .I2(duty[6]), 
            .I3(n11847), .O(n78951));
    defparam n11849_bdd_4_lut_63038.LUT_INIT = 16'he4aa;
    SB_LUT4 n78951_bdd_4_lut (.I0(n78951), .I1(duty[3]), .I2(n4925), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n78951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63033 (.I0(n11849), .I1(current[2]), .I2(duty[5]), 
            .I3(n11847), .O(n78945));
    defparam n11849_bdd_4_lut_63033.LUT_INIT = 16'he4aa;
    SB_LUT4 n78945_bdd_4_lut (.I0(n78945), .I1(duty[2]), .I2(n4926), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n78945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15814_3_lut_4_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30026));   // verilog/coms.v(130[12] 305[6])
    defparam i15814_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n11849_bdd_4_lut_63028 (.I0(n11849), .I1(current[1]), .I2(duty[4]), 
            .I3(n11847), .O(n78939));
    defparam n11849_bdd_4_lut_63028.LUT_INIT = 16'he4aa;
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n64350));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i15813_3_lut_4_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30025));   // verilog/coms.v(130[12] 305[6])
    defparam i15813_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15812_3_lut_4_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30024));   // verilog/coms.v(130[12] 305[6])
    defparam i15812_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n78939_bdd_4_lut (.I0(n78939), .I1(duty[1]), .I2(n4927), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n78939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5910));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5909));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5908));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5907));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5906));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15811_3_lut_4_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30023));   // verilog/coms.v(130[12] 305[6])
    defparam i15811_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n11849_bdd_4_lut_63023 (.I0(n11849), .I1(current[0]), .I2(duty[3]), 
            .I3(n11847), .O(n78933));
    defparam n11849_bdd_4_lut_63023.LUT_INIT = 16'he4aa;
    SB_LUT4 i15810_3_lut_4_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30022));   // verilog/coms.v(130[12] 305[6])
    defparam i15810_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15809_3_lut_4_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30021));   // verilog/coms.v(130[12] 305[6])
    defparam i15809_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n78071), .I1(n2313), 
            .I2(VCC_net), .I3(n58809), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n58808), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n58808), .I0(n2314), 
            .I1(VCC_net), .CO(n58809));
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n58807), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n58807), .I0(n2315), 
            .I1(VCC_net), .CO(n58808));
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n58806), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n78933_bdd_4_lut (.I0(n78933), .I1(duty[0]), .I2(n4928), .I3(n11847), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n78933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n58806), .I0(n2316), 
            .I1(VCC_net), .CO(n58807));
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n58805), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n58805), .I0(n2317), 
            .I1(VCC_net), .CO(n58806));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n66000));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15808_3_lut_4_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30020));   // verilog/coms.v(130[12] 305[6])
    defparam i15808_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n58804), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n58804), .I0(n2318), 
            .I1(VCC_net), .CO(n58805));
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n58803), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n58803), .I0(n2319), 
            .I1(VCC_net), .CO(n58804));
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n58802), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n58802), .I0(n2320), 
            .I1(VCC_net), .CO(n58803));
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n58801), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n58801), .I0(n2321), 
            .I1(VCC_net), .CO(n58802));
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n58800), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5831));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n58800), .I0(n2322), 
            .I1(VCC_net), .CO(n58801));
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n58799), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n58799), .I0(n2323), 
            .I1(VCC_net), .CO(n58800));
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n58798), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n58798), .I0(n2324), 
            .I1(VCC_net), .CO(n58799));
    SB_LUT4 i15807_3_lut_4_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30019));   // verilog/coms.v(130[12] 305[6])
    defparam i15807_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15806_3_lut_4_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30018));   // verilog/coms.v(130[12] 305[6])
    defparam i15806_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n65999));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n58797), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n58797), .I0(n2325), 
            .I1(VCC_net), .CO(n58798));
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n58796), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n58796), .I0(n2326), 
            .I1(VCC_net), .CO(n58797));
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n58795), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n58795), .I0(n2327), 
            .I1(VCC_net), .CO(n58796));
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n58794), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n65854));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n58794), .I0(n2328), 
            .I1(VCC_net), .CO(n58795));
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n58793), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n58793), .I0(n2329), 
            .I1(GND_net), .CO(n58794));
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n58792), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n58792), .I0(n2330), 
            .I1(GND_net), .CO(n58793));
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n58791), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n58791), .I0(n2331), 
            .I1(VCC_net), .CO(n58792));
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n58790), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n58790), .I0(n2332), 
            .I1(GND_net), .CO(n58791));
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n58789), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n58789), .I0(n2333), 
            .I1(VCC_net), .CO(n58790));
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5905));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n58789));
    SB_LUT4 i15798_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n30010));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5904));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n65998));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n65997));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5903));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1948 (.I0(control_mode[1]), .I1(n35278), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15_adj_5825));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1948.LUT_INIT = 16'hfdfd;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n58291), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n58291), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n58292));
    SB_LUT4 i15793_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n30005));   // verilog/coms.v(130[12] 305[6])
    defparam i15793_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5902));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n58395), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n66003));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n65996));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5901));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n66040));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5900));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(n78105), .I1(n2214), 
            .I2(VCC_net), .I3(n58769), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n58768), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5899));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n58768), .I0(n2215), 
            .I1(VCC_net), .CO(n58769));
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n58767), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n58767), .I0(n2216), 
            .I1(VCC_net), .CO(n58768));
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n58766), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n58394), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n58394), .I0(GND_net), .I1(n2), 
            .CO(n58395));
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n58766), .I0(n2217), 
            .I1(VCC_net), .CO(n58767));
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n58765), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n58765), .I0(n2218), 
            .I1(VCC_net), .CO(n58766));
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n58764), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5718), 
            .I3(n58393), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5898));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5897));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n58145), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n58393), .I0(GND_net), .I1(n14_adj_5718), 
            .CO(n58394));
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n58764), .I0(n2219), 
            .I1(VCC_net), .CO(n58765));
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28128), 
            .D(n1239), .R(n29176));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n58763), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n58763), .I0(n2220), 
            .I1(VCC_net), .CO(n58764));
    SB_LUT4 i1_4_lut_adj_1952 (.I0(n2329), .I1(n45309), .I2(n2330), .I3(n2331), 
            .O(n67787));
    defparam i1_4_lut_adj_1952.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5896));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1953 (.I0(n2319), .I1(n70291), .I2(n2323), .I3(n2327), 
            .O(n70295));
    defparam i1_4_lut_adj_1953.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n58762), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5895));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n58762), .I0(n2221), 
            .I1(VCC_net), .CO(n58763));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5719), 
            .I3(n58392), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n58392), .I0(GND_net), .I1(n15_adj_5719), 
            .CO(n58393));
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n58761), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n58761), .I0(n2222), 
            .I1(VCC_net), .CO(n58762));
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n58760), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n58760), .I0(n2223), 
            .I1(VCC_net), .CO(n58761));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5720), 
            .I3(n58391), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n58391), .I0(GND_net), .I1(n16_adj_5720), 
            .CO(n58392));
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n58759), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n58759), .I0(n2224), 
            .I1(VCC_net), .CO(n58760));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5894));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n58758), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n58758), .I0(n2225), 
            .I1(VCC_net), .CO(n58759));
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n58757), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n58757), .I0(n2226), 
            .I1(VCC_net), .CO(n58758));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n58756), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n58756), .I0(n2227), 
            .I1(VCC_net), .CO(n58757));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n65995));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n58755), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n58755), .I0(n2228), 
            .I1(VCC_net), .CO(n58756));
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n58754), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n28049), .D(GHC_N_391), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n28049), .D(GHB_N_377), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n28049), .D(GHA_N_355), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5976), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n58754), .I0(n2229), 
            .I1(GND_net), .CO(n58755));
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n28049), .D(GLA_N_372), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n58753), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n28049), .D(GLB_N_386), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n28049), .D(GLC_N_400), 
            .R(n29153));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n58753), .I0(n2230), 
            .I1(GND_net), .CO(n58754));
    GND i1 (.Y(GND_net));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n65994));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5721), 
            .I3(n58390), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n58390), .I0(GND_net), .I1(n17_adj_5721), 
            .CO(n58391));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5893));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5892));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n65993));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n58752), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n58752), .I0(n2231), 
            .I1(VCC_net), .CO(n58753));
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n58751), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n65992));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n58751), .I0(n2232), 
            .I1(GND_net), .CO(n58752));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5722), 
            .I3(n58389), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n58750), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n58750), .I0(n2233), 
            .I1(VCC_net), .CO(n58751));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n58389), .I0(GND_net), .I1(n18_adj_5722), 
            .CO(n58390));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25), .CO(n58291));
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5891));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5890));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n58750));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5889));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5723), 
            .I3(n58388), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5888));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5887));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n58388), .I0(GND_net), .I1(n19_adj_5723), 
            .CO(n58389));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5724), 
            .I3(n58387), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n65991));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n65990));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n58387), .I0(GND_net), .I1(n20_adj_5724), 
            .CO(n58388));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5725), 
            .I3(n58386), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n65989));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n58386), .I0(GND_net), .I1(n21_adj_5725), 
            .CO(n58387));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n65855));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n65988));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n65987));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5726), 
            .I3(n58385), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n58385), .I0(GND_net), .I1(n22_adj_5726), 
            .CO(n58386));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n65986));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5727), 
            .I3(n58384), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n58384), .I0(GND_net), .I1(n23_adj_5727), 
            .CO(n58385));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5728), 
            .I3(n58383), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n58383), .I0(GND_net), .I1(n24_adj_5728), 
            .CO(n58384));
    SB_LUT4 i7_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5879));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10_2_lut (.I0(PWMLimit[18]), .I1(setpoint[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n45105), .I1(GND_net), .I2(n25_adj_5729), 
            .I3(VCC_net), .O(n74445)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5873));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5729), 
            .CO(n58383));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n65985));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n58138), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20512_3_lut (.I0(n16_adj_5874), .I1(PWMLimit[8]), .I2(setpoint[8]), 
            .I3(GND_net), .O(n34707));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i20512_3_lut.LUT_INIT = 16'hb2b2;
    SB_CARRY add_151_11 (.CI(n58145), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n58146));
    SB_LUT4 i9_2_lut (.I0(PWMLimit[12]), .I1(setpoint[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5877));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(n78132), .I1(n2115), 
            .I2(VCC_net), .I3(n58723), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n58722), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n58722), .I0(n2116), 
            .I1(VCC_net), .CO(n58723));
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n58721), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n58721), .I0(n2117), 
            .I1(VCC_net), .CO(n58722));
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n58720), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n58720), .I0(n2118), 
            .I1(VCC_net), .CO(n58721));
    SB_LUT4 i7_2_lut_adj_1966 (.I0(PWMLimit[16]), .I1(setpoint[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5878));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i7_2_lut_adj_1966.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n58719), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n58719), .I0(n2119), 
            .I1(VCC_net), .CO(n58720));
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n58718), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n58718), .I0(n2120), 
            .I1(VCC_net), .CO(n58719));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n65984));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n65983));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n58717), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n58717), .I0(n2121), 
            .I1(VCC_net), .CO(n58718));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n58716), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n58716), .I0(n2122), 
            .I1(VCC_net), .CO(n58717));
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n58715), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23733_3_lut (.I0(n20_adj_5875), .I1(PWMLimit[10]), .I2(setpoint[10]), 
            .I3(GND_net), .O(n22_adj_5876));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i23733_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 mux_3812_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5739), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n58715), .I0(n2123), 
            .I1(VCC_net), .CO(n58716));
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n58714), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n58714), .I0(n2124), 
            .I1(VCC_net), .CO(n58715));
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n58713), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n58713), .I0(n2125), 
            .I1(VCC_net), .CO(n58714));
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n58712), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n58712), .I0(n2126), 
            .I1(VCC_net), .CO(n58713));
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n58711), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n58711), .I0(n2127), 
            .I1(VCC_net), .CO(n58712));
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n58710), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n58710), .I0(n2128), 
            .I1(VCC_net), .CO(n58711));
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n58709), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n58709), .I0(n2129), 
            .I1(GND_net), .CO(n58710));
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n58708), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n58708), .I0(n2130), 
            .I1(GND_net), .CO(n58709));
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n58707), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n58707), .I0(n2131), 
            .I1(VCC_net), .CO(n58708));
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n58706), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n58706), .I0(n2132), 
            .I1(GND_net), .CO(n58707));
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n58705), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n58705), .I0(n2133), 
            .I1(VCC_net), .CO(n58706));
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n58705));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n65982));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n65981));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n65980));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n65979));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n65978));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n78128), .I1(n2016), 
            .I2(VCC_net), .I3(n58687), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n58686), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n58686), .I0(n2017), 
            .I1(VCC_net), .CO(n58687));
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n58685), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n58685), .I0(n2018), 
            .I1(VCC_net), .CO(n58686));
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n58684), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n58684), .I0(n2019), 
            .I1(VCC_net), .CO(n58685));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n65977));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n65976));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n58683), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n58683), .I0(n2020), 
            .I1(VCC_net), .CO(n58684));
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n58682), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n58167), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n58682), .I0(n2021), 
            .I1(VCC_net), .CO(n58683));
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n58166), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n65975));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n58681), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n58681), .I0(n2022), 
            .I1(VCC_net), .CO(n58682));
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n58680), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n65871));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n58680), .I0(n2023), 
            .I1(VCC_net), .CO(n58681));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n65973));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n58679), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n58679), .I0(n2024), 
            .I1(VCC_net), .CO(n58680));
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n58678), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n58678), .I0(n2025), 
            .I1(VCC_net), .CO(n58679));
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n58677), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n58677), .I0(n2026), 
            .I1(VCC_net), .CO(n58678));
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n58676), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n58676), .I0(n2027), 
            .I1(VCC_net), .CO(n58677));
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n58675), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n58675), .I0(n2028), 
            .I1(VCC_net), .CO(n58676));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n58674), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n58674), .I0(n2029), 
            .I1(GND_net), .CO(n58675));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n58673), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n58673), .I0(n2030), 
            .I1(GND_net), .CO(n58674));
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n58672), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n58672), .I0(n2031), 
            .I1(VCC_net), .CO(n58673));
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n58671), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n58671), .I0(n2032), 
            .I1(GND_net), .CO(n58672));
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n58670), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n58670), .I0(n2033), 
            .I1(VCC_net), .CO(n58671));
    SB_LUT4 i12_2_lut (.I0(PWMLimit[4]), .I1(n475), .I2(GND_net), .I3(GND_net), 
            .O(n35808));
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n58670));
    SB_CARRY add_151_32 (.CI(n58166), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n58167));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5887), .I3(n59170), .O(n2_adj_5751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5888), .I3(n59169), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n59169), 
            .I0(GND_net), .I1(n3_adj_5888), .CO(n59170));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n65972));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5889), .I3(n59168), .O(n4_adj_5750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n59168), 
            .I0(GND_net), .I1(n4_adj_5889), .CO(n59169));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5890), .I3(n59167), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n59167), 
            .I0(GND_net), .I1(n5_adj_5890), .CO(n59168));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5891), .I3(n59166), .O(n6_adj_5749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n59166), 
            .I0(GND_net), .I1(n6_adj_5891), .CO(n59167));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5892), .I3(n59165), .O(n7_adj_5748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n59165), 
            .I0(GND_net), .I1(n7_adj_5892), .CO(n59166));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5893), .I3(n59164), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n59164), 
            .I0(GND_net), .I1(n8_adj_5893), .CO(n59165));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5894), .I3(n59163), .O(n9_adj_5746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n59163), 
            .I0(GND_net), .I1(n9_adj_5894), .CO(n59164));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5895), .I3(n59162), .O(n10_adj_5745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n59162), 
            .I0(GND_net), .I1(n10_adj_5895), .CO(n59163));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5896), .I3(n59161), .O(n11_adj_5744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n59161), 
            .I0(GND_net), .I1(n11_adj_5896), .CO(n59162));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5897), .I3(n59160), .O(n12_adj_5743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n59160), 
            .I0(GND_net), .I1(n12_adj_5897), .CO(n59161));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5898), .I3(n59159), .O(n13_adj_5742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n59159), 
            .I0(GND_net), .I1(n13_adj_5898), .CO(n59160));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5899), .I3(n59158), .O(n14_adj_5741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n59158), 
            .I0(GND_net), .I1(n14_adj_5899), .CO(n59159));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5900), .I3(n59157), .O(n15_adj_5740)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(n77874), .I1(n1917), 
            .I2(VCC_net), .I3(n58646), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n59157), 
            .I0(GND_net), .I1(n15_adj_5900), .CO(n59158));
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n58645), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5901), .I3(n59156), .O(n16_adj_5739)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n59156), 
            .I0(GND_net), .I1(n16_adj_5901), .CO(n59157));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5902), .I3(n59155), .O(n17_adj_5738)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n58645), .I0(n1918), 
            .I1(VCC_net), .CO(n58646));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n59155), 
            .I0(GND_net), .I1(n17_adj_5902), .CO(n59156));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5903), .I3(n59154), .O(n18_adj_5737)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n58644), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n58644), .I0(n1919), 
            .I1(VCC_net), .CO(n58645));
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n58643), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n58643), .I0(n1920), 
            .I1(VCC_net), .CO(n58644));
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n58642), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n59154), 
            .I0(GND_net), .I1(n18_adj_5903), .CO(n59155));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5904), .I3(n59153), .O(n19_adj_5736)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n58642), .I0(n1921), 
            .I1(VCC_net), .CO(n58643));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n59153), 
            .I0(GND_net), .I1(n19_adj_5904), .CO(n59154));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n58641), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5905), .I3(n59152), .O(n20_adj_5735)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n58641), .I0(n1922), 
            .I1(VCC_net), .CO(n58642));
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n58640), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n59152), 
            .I0(GND_net), .I1(n20_adj_5905), .CO(n59153));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5906), .I3(n59151), .O(n21_adj_5734)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n59151), 
            .I0(GND_net), .I1(n21_adj_5906), .CO(n59152));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5907), .I3(n59150), .O(n22_adj_5733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n58640), .I0(n1923), 
            .I1(VCC_net), .CO(n58641));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n59150), 
            .I0(GND_net), .I1(n22_adj_5907), .CO(n59151));
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n58639), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5908), .I3(n59149), .O(n23_adj_5732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n58639), .I0(n1924), 
            .I1(VCC_net), .CO(n58640));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n59149), 
            .I0(GND_net), .I1(n23_adj_5908), .CO(n59150));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n65971));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5909), .I3(n59148), .O(n24_adj_5731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n59148), 
            .I0(GND_net), .I1(n24_adj_5909), .CO(n59149));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n58638), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n58638), .I0(n1925), 
            .I1(VCC_net), .CO(n58639));
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n58637), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n58637), .I0(n1926), 
            .I1(VCC_net), .CO(n58638));
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n58636), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5910), .I3(n59147), .O(n25_adj_5730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n58636), .I0(n1927), 
            .I1(VCC_net), .CO(n58637));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n59147), 
            .I0(GND_net), .I1(n25_adj_5910), .CO(n59148));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5911), .I3(n59146), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n59146), 
            .I0(GND_net), .I1(n26_adj_5911), .CO(n59147));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5912), .I3(n59145), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n59145), 
            .I0(GND_net), .I1(n27_adj_5912), .CO(n59146));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5913), .I3(n59144), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n59144), 
            .I0(GND_net), .I1(n28_adj_5913), .CO(n59145));
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n58635), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n58635), .I0(n1928), 
            .I1(VCC_net), .CO(n58636));
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n58634), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n58634), .I0(n1929), 
            .I1(GND_net), .CO(n58635));
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n58633), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5914), .I3(n59143), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n59143), 
            .I0(GND_net), .I1(n29_adj_5914), .CO(n59144));
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n58633), .I0(n1930), 
            .I1(GND_net), .CO(n58634));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n58632), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5915), .I3(n59142), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n59142), 
            .I0(GND_net), .I1(n30_adj_5915), .CO(n59143));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n65970));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5916), .I3(n59141), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n58632), .I0(n1931), 
            .I1(VCC_net), .CO(n58633));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n65969));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n65968));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n59141), 
            .I0(GND_net), .I1(n31_adj_5916), .CO(n59142));
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n58631), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n58631), .I0(n1932), 
            .I1(GND_net), .CO(n58632));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5917), .I3(n59140), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n58630), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n58630), .I0(n1933), 
            .I1(VCC_net), .CO(n58631));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n59140), 
            .I0(GND_net), .I1(n32_adj_5917), .CO(n59141));
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n58630));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n59140));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n65967));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 add_2634_25_lut (.I0(n78310), .I1(n2_adj_5887), .I2(n1059), 
            .I3(n59139), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1985 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n65966));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1985.LUT_INIT = 16'h2300;
    SB_LUT4 add_2634_24_lut (.I0(n78239), .I1(n2_adj_5887), .I2(n1158), 
            .I3(n59138), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_24 (.CI(n59138), .I0(n2_adj_5887), .I1(n1158), .CO(n59139));
    SB_LUT4 add_2634_23_lut (.I0(n78264), .I1(n2_adj_5887), .I2(n1257), 
            .I3(n59137), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_23 (.CI(n59137), .I0(n2_adj_5887), .I1(n1257), .CO(n59138));
    SB_LUT4 add_2634_22_lut (.I0(n78268), .I1(n2_adj_5887), .I2(n1356), 
            .I3(n59136), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_22 (.CI(n59136), .I0(n2_adj_5887), .I1(n1356), .CO(n59137));
    SB_LUT4 add_2634_21_lut (.I0(n78284), .I1(n2_adj_5887), .I2(n1455), 
            .I3(n59135), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_21 (.CI(n59135), .I0(n2_adj_5887), .I1(n1455), .CO(n59136));
    SB_LUT4 add_2634_20_lut (.I0(n78225), .I1(n2_adj_5887), .I2(n1554), 
            .I3(n59134), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_20 (.CI(n59134), .I0(n2_adj_5887), .I1(n1554), .CO(n59135));
    SB_LUT4 add_2634_19_lut (.I0(n78030), .I1(n2_adj_5887), .I2(n1653), 
            .I3(n59133), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n65965));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_CARRY add_2634_19 (.CI(n59133), .I0(n2_adj_5887), .I1(n1653), .CO(n59134));
    SB_LUT4 i22001_3_lut (.I0(n24_adj_5886), .I1(PWMLimit[12]), .I2(n467), 
            .I3(GND_net), .O(n36173));
    defparam i22001_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 add_2634_18_lut (.I0(n78320), .I1(n2_adj_5887), .I2(n1752), 
            .I3(n59132), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_18 (.CI(n59132), .I0(n2_adj_5887), .I1(n1752), .CO(n59133));
    SB_LUT4 add_2634_17_lut (.I0(n78370), .I1(n2_adj_5887), .I2(n1851), 
            .I3(n59131), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_17 (.CI(n59131), .I0(n2_adj_5887), .I1(n1851), .CO(n59132));
    SB_LUT4 add_2634_16_lut (.I0(n77874), .I1(n2_adj_5887), .I2(n1950), 
            .I3(n59130), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_16 (.CI(n59130), .I0(n2_adj_5887), .I1(n1950), .CO(n59131));
    SB_LUT4 add_2634_15_lut (.I0(n78128), .I1(n2_adj_5887), .I2(n2049), 
            .I3(n59129), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_15 (.CI(n59129), .I0(n2_adj_5887), .I1(n2049), .CO(n59130));
    SB_LUT4 add_2634_14_lut (.I0(n78132), .I1(n2_adj_5887), .I2(n2148), 
            .I3(n59128), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n65964));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_CARRY add_2634_14 (.CI(n59128), .I0(n2_adj_5887), .I1(n2148), .CO(n59129));
    SB_LUT4 add_2634_13_lut (.I0(n78105), .I1(n2_adj_5887), .I2(n2247), 
            .I3(n59127), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_13 (.CI(n59127), .I0(n2_adj_5887), .I1(n2247), .CO(n59128));
    SB_LUT4 add_2634_12_lut (.I0(n78071), .I1(n2_adj_5887), .I2(n2346), 
            .I3(n59126), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_12 (.CI(n59126), .I0(n2_adj_5887), .I1(n2346), .CO(n59127));
    SB_LUT4 add_2634_11_lut (.I0(n77940), .I1(n2_adj_5887), .I2(n2445), 
            .I3(n59125), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_11 (.CI(n59125), .I0(n2_adj_5887), .I1(n2445), .CO(n59126));
    SB_LUT4 add_2634_10_lut (.I0(n78023), .I1(n2_adj_5887), .I2(n2544), 
            .I3(n59124), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_10 (.CI(n59124), .I0(n2_adj_5887), .I1(n2544), .CO(n59125));
    SB_LUT4 add_2634_9_lut (.I0(n77967), .I1(n2_adj_5887), .I2(n2643), 
            .I3(n59123), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_9 (.CI(n59123), .I0(n2_adj_5887), .I1(n2643), .CO(n59124));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n65963));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 add_2634_8_lut (.I0(n78340), .I1(n2_adj_5887), .I2(n2742), 
            .I3(n59122), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_8 (.CI(n59122), .I0(n2_adj_5887), .I1(n2742), .CO(n59123));
    SB_LUT4 add_1190_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n58259), .O(n4905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2634_7_lut (.I0(n78418), .I1(n2_adj_5887), .I2(n2841), 
            .I3(n59121), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_7 (.CI(n59121), .I0(n2_adj_5887), .I1(n2841), .CO(n59122));
    SB_LUT4 add_2634_6_lut (.I0(n77679), .I1(n2_adj_5887), .I2(n2940), 
            .I3(n59120), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_6 (.CI(n59120), .I0(n2_adj_5887), .I1(n2940), .CO(n59121));
    SB_LUT4 add_2634_5_lut (.I0(n77736), .I1(n2_adj_5887), .I2(n3039), 
            .I3(n59119), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_5 (.CI(n59119), .I0(n2_adj_5887), .I1(n3039), .CO(n59120));
    SB_LUT4 add_2634_4_lut (.I0(n77776), .I1(n2_adj_5887), .I2(n3138), 
            .I3(n59118), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2634_4 (.CI(n59118), .I0(n2_adj_5887), .I1(n3138), .CO(n59119));
    SB_LUT4 add_2634_3_lut (.I0(n77824), .I1(n2_adj_5887), .I2(n3237), 
            .I3(n59117), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1190_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12448), 
            .I3(n58258), .O(n4906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n65962));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_CARRY add_2634_3 (.CI(n59117), .I0(n2_adj_5887), .I1(n3237), .CO(n59118));
    SB_CARRY add_1190_24 (.CI(n58258), .I0(GND_net), .I1(n12448), .CO(n58259));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n58165), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2634_2_lut (.I0(n77878), .I1(n2_adj_5887), .I2(n45345), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2634_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1190_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12450), 
            .I3(n58257), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n58165), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n58166));
    SB_CARRY add_2634_2 (.CI(VCC_net), .I0(n2_adj_5887), .I1(n45345), 
            .CO(n59117));
    SB_CARRY add_1190_23 (.CI(n58257), .I0(GND_net), .I1(n12450), .CO(n58258));
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(n77824), .I1(n3204), 
            .I2(VCC_net), .I3(n59116), .O(n71361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1190_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12452), 
            .I3(n58256), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n58144), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1990 (.I0(\data_out_frame[19] [3]), .I1(n66450), 
            .I2(n66594), .I3(n60646), .O(n60808));
    defparam i1_4_lut_adj_1990.LUT_INIT = 16'h9669;
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n58164), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n59115), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_22 (.CI(n58256), .I0(GND_net), .I1(n12452), .CO(n58257));
    SB_CARRY add_151_30 (.CI(n58164), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n58165));
    SB_CARRY add_151_4 (.CI(n58138), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n58139));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n58163), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15744_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5803), .I2(a_new_adj_6018[1]), 
            .I3(position_31__N_3836_adj_5805), .O(n29956));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n65961));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i15742_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_6055[1]), 
            .I2(r_SM_Main_adj_6055[2]), .I3(n6_adj_5954), .O(n29954));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15742_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n65960));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n59115), .I0(n3205), 
            .I1(VCC_net), .CO(n59116));
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n59114), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n59114), .I0(n3206), 
            .I1(VCC_net), .CO(n59115));
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n59113), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n59113), .I0(n3207), 
            .I1(VCC_net), .CO(n59114));
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n59112), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12454), 
            .I3(n58255), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_10 (.CI(n58144), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n58145));
    SB_CARRY add_151_29 (.CI(n58163), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n58164));
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n59112), .I0(n3208), 
            .I1(VCC_net), .CO(n59113));
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(n78370), .I1(n1818), 
            .I2(VCC_net), .I3(n58614), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1190_21 (.CI(n58255), .I0(GND_net), .I1(n12454), .CO(n58256));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n58162), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n59111), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n59111), .I0(n3209), 
            .I1(VCC_net), .CO(n59112));
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n59110), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n59110), .I0(n3210), 
            .I1(VCC_net), .CO(n59111));
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n59109), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n59109), .I0(n3211), 
            .I1(VCC_net), .CO(n59110));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n59108), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n59108), .I0(n3212), 
            .I1(VCC_net), .CO(n59109));
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n59107), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n58613), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n58613), .I0(n1819), 
            .I1(VCC_net), .CO(n58614));
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n58612), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n59107), .I0(n3213), 
            .I1(VCC_net), .CO(n59108));
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n58612), .I0(n1820), 
            .I1(VCC_net), .CO(n58613));
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n58611), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n59106), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n58611), .I0(n1821), 
            .I1(VCC_net), .CO(n58612));
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n59106), .I0(n3214), 
            .I1(VCC_net), .CO(n59107));
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n58610), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n59105), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n59105), .I0(n3215), 
            .I1(VCC_net), .CO(n59106));
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n58610), .I0(n1822), 
            .I1(VCC_net), .CO(n58611));
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n58609), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12456), 
            .I3(n58254), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n59104), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n58609), .I0(n1823), 
            .I1(VCC_net), .CO(n58610));
    SB_CARRY add_1190_20 (.CI(n58254), .I0(GND_net), .I1(n12456), .CO(n58255));
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n59104), .I0(n3216), 
            .I1(VCC_net), .CO(n59105));
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n58608), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12458), 
            .I3(n58253), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n59103), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n58608), .I0(n1824), 
            .I1(VCC_net), .CO(n58609));
    SB_CARRY add_1190_19 (.CI(n58253), .I0(GND_net), .I1(n12458), .CO(n58254));
    SB_CARRY add_151_28 (.CI(n58162), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n58163));
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n59103), .I0(n3217), 
            .I1(VCC_net), .CO(n59104));
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n58607), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12460), 
            .I3(n58252), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n59102), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n58607), .I0(n1825), 
            .I1(VCC_net), .CO(n58608));
    SB_CARRY add_1190_18 (.CI(n58252), .I0(GND_net), .I1(n12460), .CO(n58253));
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n58143), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n59102), .I0(n3218), 
            .I1(VCC_net), .CO(n59103));
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n58606), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12462), 
            .I3(n58251), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n58161), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_27 (.CI(n58161), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n58162));
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n59101), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n58606), .I0(n1826), 
            .I1(VCC_net), .CO(n58607));
    SB_CARRY add_1190_17 (.CI(n58251), .I0(GND_net), .I1(n12462), .CO(n58252));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n58160), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n58137), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n59101), .I0(n3219), 
            .I1(VCC_net), .CO(n59102));
    SB_LUT4 i1_4_lut_adj_1993 (.I0(n2316), .I1(n2318), .I2(n2320), .I3(n70243), 
            .O(n70249));
    defparam i1_4_lut_adj_1993.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n59100), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n59100), .I0(n3220), 
            .I1(VCC_net), .CO(n59101));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n59099), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n59099), .I0(n3221), 
            .I1(VCC_net), .CO(n59100));
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n59098), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n59098), .I0(n3222), 
            .I1(VCC_net), .CO(n59099));
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n59097), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23467_3_lut_4_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n29942));
    defparam i23467_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n59097), .I0(n3223), 
            .I1(VCC_net), .CO(n59098));
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n58605), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n59096), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12464), 
            .I3(n58250), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n59096), .I0(n3224), 
            .I1(VCC_net), .CO(n59097));
    SB_CARRY add_1190_16 (.CI(n58250), .I0(GND_net), .I1(n12464), .CO(n58251));
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n59095), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n58605), .I0(n1827), 
            .I1(VCC_net), .CO(n58606));
    SB_LUT4 add_1190_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12466), 
            .I3(n58249), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n59095), .I0(n3225), 
            .I1(VCC_net), .CO(n59096));
    SB_CARRY add_1190_15 (.CI(n58249), .I0(GND_net), .I1(n12466), .CO(n58250));
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n59094), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n58604), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n58604), .I0(n1828), 
            .I1(VCC_net), .CO(n58605));
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n58603), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n59094), .I0(n3226), 
            .I1(VCC_net), .CO(n59095));
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n59093), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12468), 
            .I3(n58248), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n59093), .I0(n3227), 
            .I1(VCC_net), .CO(n59094));
    SB_CARRY add_1190_14 (.CI(n58248), .I0(GND_net), .I1(n12468), .CO(n58249));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n59092), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n58603), .I0(n1829), 
            .I1(GND_net), .CO(n58604));
    SB_LUT4 add_1190_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12470), 
            .I3(n58247), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n59092), .I0(n3228), 
            .I1(VCC_net), .CO(n59093));
    SB_CARRY add_1190_13 (.CI(n58247), .I0(GND_net), .I1(n12470), .CO(n58248));
    SB_CARRY add_151_9 (.CI(n58143), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n58144));
    SB_CARRY add_151_26 (.CI(n58160), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n58161));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n59091), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n59091), .I0(n3229), 
            .I1(GND_net), .CO(n59092));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n59090), .O(n74442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n59090), .I0(n3230), 
            .I1(GND_net), .CO(n59091));
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n59089), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n59089), .I0(n3231), 
            .I1(VCC_net), .CO(n59090));
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5919), .I1(n3232), 
            .I2(GND_net), .I3(n59088), .O(n74590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n59088), .I0(n3232), 
            .I1(GND_net), .CO(n59089));
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n59087), .O(n6_adj_5919)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n59087), .I0(n3233), 
            .I1(VCC_net), .CO(n59088));
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n58602), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12472), 
            .I3(n58246), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n59086), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_12 (.CI(n58246), .I0(GND_net), .I1(n12472), .CO(n58247));
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n59086), .I0(n957), 
            .I1(GND_net), .CO(n59087));
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n58602), .I0(n1830), 
            .I1(GND_net), .CO(n58603));
    SB_LUT4 add_1190_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12474), 
            .I3(n58245), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n59086));
    SB_CARRY add_1190_11 (.CI(n58245), .I0(GND_net), .I1(n12474), .CO(n58246));
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n77776), .I1(n3105), 
            .I2(VCC_net), .I3(n59085), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n58601), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12476), 
            .I3(n58244), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n59084), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_10 (.CI(n58244), .I0(GND_net), .I1(n12476), .CO(n58245));
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n59084), .I0(n3106), 
            .I1(VCC_net), .CO(n59085));
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n58601), .I0(n1831), 
            .I1(VCC_net), .CO(n58602));
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n58600), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12478), .I3(n58243), 
            .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n59083), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_9 (.CI(n58243), .I0(GND_net), .I1(n12478), .CO(n58244));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n58159), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n59083), .I0(n3107), 
            .I1(VCC_net), .CO(n59084));
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n59082), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n59082), .I0(n3108), 
            .I1(VCC_net), .CO(n59083));
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n59081), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n59081), .I0(n3109), 
            .I1(VCC_net), .CO(n59082));
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n59080), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n59080), .I0(n3110), 
            .I1(VCC_net), .CO(n59081));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n59079), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n58600), .I0(n1832), 
            .I1(GND_net), .CO(n58601));
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n59079), .I0(n3111), 
            .I1(VCC_net), .CO(n59080));
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n58599), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12480), .I3(n58242), 
            .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n59078), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_8 (.CI(n58242), .I0(GND_net), .I1(n12480), .CO(n58243));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n58142), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_25 (.CI(n58159), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n58160));
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n59078), .I0(n3112), 
            .I1(VCC_net), .CO(n59079));
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n59077), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n58599), .I0(n1833), 
            .I1(VCC_net), .CO(n58600));
    SB_LUT4 add_1190_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12482), .I3(n58241), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_3 (.CI(n58137), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n58138));
    SB_CARRY add_151_8 (.CI(n58142), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n58143));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n58158), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n59077), .I0(n3113), 
            .I1(VCC_net), .CO(n59078));
    SB_CARRY add_1190_7 (.CI(n58241), .I0(GND_net), .I1(n12482), .CO(n58242));
    SB_CARRY add_151_24 (.CI(n58158), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n58159));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n58157), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n58157), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n58158));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n59076), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n59076), .I0(n3114), 
            .I1(VCC_net), .CO(n59077));
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n58599));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n59075), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n59075), .I0(n3115), 
            .I1(VCC_net), .CO(n59076));
    SB_LUT4 add_1190_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12484), .I3(n58240), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n59074), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n59074), .I0(n3116), 
            .I1(VCC_net), .CO(n59075));
    SB_CARRY add_1190_6 (.CI(n58240), .I0(GND_net), .I1(n12484), .CO(n58241));
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n59073), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n59073), .I0(n3117), 
            .I1(VCC_net), .CO(n59074));
    SB_LUT4 add_1190_5_lut (.I0(GND_net), .I1(GND_net), .I2(n12486), .I3(n58239), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_5 (.CI(n58239), .I0(GND_net), .I1(n12486), .CO(n58240));
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n59072), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n59072), .I0(n3118), 
            .I1(VCC_net), .CO(n59073));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n59071), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n59071), .I0(n3119), 
            .I1(VCC_net), .CO(n59072));
    SB_LUT4 add_1190_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12488), .I3(n58238), 
            .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n58156), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_22 (.CI(n58156), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n58157));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n58155), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_21 (.CI(n58155), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n58156));
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n59070), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_4 (.CI(n58238), .I0(GND_net), .I1(n12488), .CO(n58239));
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n59070), .I0(n3120), 
            .I1(VCC_net), .CO(n59071));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n59069), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n59069), .I0(n3121), 
            .I1(VCC_net), .CO(n59070));
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n59068), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n59068), .I0(n3122), 
            .I1(VCC_net), .CO(n59069));
    SB_LUT4 i55932_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71767));
    defparam i55932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15726_3_lut_4_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n29938));   // verilog/coms.v(130[12] 305[6])
    defparam i15726_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i55933_4_lut (.I0(n71767), .I1(n44122), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n71768));
    defparam i55933_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n59067), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i55931_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71766));
    defparam i55931_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n59067), .I0(n3123), 
            .I1(VCC_net), .CO(n59068));
    SB_LUT4 i15725_3_lut_4_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n29937));   // verilog/coms.v(130[12] 305[6])
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n59066), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12490), .I3(n58237), 
            .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n59066), .I0(n3124), 
            .I1(VCC_net), .CO(n59067));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n59065), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n59065), .I0(n3125), 
            .I1(VCC_net), .CO(n59066));
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n59064), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n59064), .I0(n3126), 
            .I1(VCC_net), .CO(n59065));
    SB_CARRY add_1190_3 (.CI(n58237), .I0(GND_net), .I1(n12490), .CO(n58238));
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n59063), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_2_lut (.I0(GND_net), .I1(GND_net), .I2(n11912), .I3(VCC_net), 
            .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n59063), .I0(n3127), 
            .I1(VCC_net), .CO(n59064));
    SB_CARRY add_1190_2 (.CI(VCC_net), .I0(GND_net), .I1(n11912), .CO(n58237));
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n59062), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n59062), .I0(n3128), 
            .I1(VCC_net), .CO(n59063));
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n59061), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n59061), .I0(n3129), 
            .I1(GND_net), .CO(n59062));
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n59060), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15724_3_lut_4_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n29936));   // verilog/coms.v(130[12] 305[6])
    defparam i15724_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n59060), .I0(n3130), 
            .I1(GND_net), .CO(n59061));
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n59059), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n58154), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n59059), .I0(n3131), 
            .I1(VCC_net), .CO(n59060));
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n59058), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n59058), .I0(n3132), 
            .I1(GND_net), .CO(n59059));
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n59057), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_20 (.CI(n58154), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n58155));
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n59057), .I0(n3133), 
            .I1(VCC_net), .CO(n59058));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n58141), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n59057));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n58153), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n77736), .I1(n3006), 
            .I2(VCC_net), .I3(n59056), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n59055), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n59055), .I0(n3007), 
            .I1(VCC_net), .CO(n59056));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n59054), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1994 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66225));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1994.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n59054), .I0(n3008), 
            .I1(VCC_net), .CO(n59055));
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n59053), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n59053), .I0(n3009), 
            .I1(VCC_net), .CO(n59054));
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n59052), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n59052), .I0(n3010), 
            .I1(VCC_net), .CO(n59053));
    SB_LUT4 i1_2_lut_adj_1995 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66270));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1995.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n59051), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n59051), .I0(n3011), 
            .I1(VCC_net), .CO(n59052));
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n59050), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n78320), .I1(n1719), 
            .I2(VCC_net), .I3(n58578), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n59050), .I0(n3012), 
            .I1(VCC_net), .CO(n59051));
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n58577), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n58577), .I0(n1720), 
            .I1(VCC_net), .CO(n58578));
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n59049), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n58576), .O(n1788_adj_5859)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n59049), .I0(n3013), 
            .I1(VCC_net), .CO(n59050));
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n58576), .I0(n1721), 
            .I1(VCC_net), .CO(n58577));
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n59048), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n58575), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n59048), .I0(n3014), 
            .I1(VCC_net), .CO(n59049));
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n58575), .I0(n1722), 
            .I1(VCC_net), .CO(n58576));
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n58574), .O(n1790_adj_5860)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n59047), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n58574), .I0(n1723), 
            .I1(VCC_net), .CO(n58575));
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n58573), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n59047), .I0(n3015), 
            .I1(VCC_net), .CO(n59048));
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n58573), .I0(n1724), 
            .I1(VCC_net), .CO(n58574));
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n58572), .O(n1792_adj_5861)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n59046), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n58572), .I0(n1725), 
            .I1(VCC_net), .CO(n58573));
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n59046), .I0(n3016), 
            .I1(VCC_net), .CO(n59047));
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n58571), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n59045), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n58571), .I0(n1726), 
            .I1(VCC_net), .CO(n58572));
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n59045), .I0(n3017), 
            .I1(VCC_net), .CO(n59046));
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n58570), .O(n1794_adj_5862)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n59044), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n58570), .I0(n1727), 
            .I1(VCC_net), .CO(n58571));
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n59044), .I0(n3018), 
            .I1(VCC_net), .CO(n59045));
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n58569), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_2_lut (.I0(deadband[12]), .I1(n467), .I2(GND_net), .I3(GND_net), 
            .O(n25_adj_5884));
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n59043), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n58569), .I0(n1728), 
            .I1(VCC_net), .CO(n58570));
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n59043), .I0(n3019), 
            .I1(VCC_net), .CO(n59044));
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n58568), .O(n1796_adj_5863)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n59042), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n58568), .I0(n1729), 
            .I1(GND_net), .CO(n58569));
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n58567), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n59042), .I0(n3020), 
            .I1(VCC_net), .CO(n59043));
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n58567), .I0(n1730), 
            .I1(GND_net), .CO(n58568));
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n58566), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n59041), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n58566), .I0(n1731), 
            .I1(VCC_net), .CO(n58567));
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n58565), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n59041), .I0(n3021), 
            .I1(VCC_net), .CO(n59042));
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n58565), .I0(n1732), 
            .I1(GND_net), .CO(n58566));
    SB_LUT4 i1_4_lut_adj_1996 (.I0(n2317), .I1(n2315), .I2(n70295), .I3(n67787), 
            .O(n69022));
    defparam i1_4_lut_adj_1996.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n58564), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n59040), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n58564), .I0(n1733), 
            .I1(VCC_net), .CO(n58565));
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n59040), .I0(n3022), 
            .I1(VCC_net), .CO(n59041));
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n58564));
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n59039), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n59039), .I0(n3023), 
            .I1(VCC_net), .CO(n59040));
    SB_LUT4 i15721_3_lut_4_lut (.I0(deadband[0]), .I1(\data_in_frame[16] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n29933));   // verilog/coms.v(130[12] 305[6])
    defparam i15721_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n59038), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n59038), .I0(n3024), 
            .I1(VCC_net), .CO(n59039));
    SB_LUT4 i6_4_lut_adj_1997 (.I0(n66270), .I1(\data_out_frame[9] [2]), 
            .I2(n66225), .I3(n34_adj_5847), .O(n14_adj_5964));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1997.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n59037), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n59037), .I0(n3025), 
            .I1(VCC_net), .CO(n59038));
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n59036), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n59036), .I0(n3026), 
            .I1(VCC_net), .CO(n59037));
    SB_LUT4 i7_4_lut_adj_1998 (.I0(\data_out_frame[13] [4]), .I1(n14_adj_5964), 
            .I2(n10_adj_5965), .I3(\data_out_frame[4] [7]), .O(n61318));   // verilog/coms.v(100[12:26])
    defparam i7_4_lut_adj_1998.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n59035), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n59035), .I0(n3027), 
            .I1(VCC_net), .CO(n59036));
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n59034), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n59034), .I0(n3028), 
            .I1(VCC_net), .CO(n59035));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n65959));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n59033), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n59033), .I0(n3029), 
            .I1(GND_net), .CO(n59034));
    SB_LUT4 i21623_3_lut (.I0(n8_adj_5882), .I1(deadband[4]), .I2(n475), 
            .I3(GND_net), .O(n10_adj_5883));
    defparam i21623_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n65958));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n59032), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n59032), .I0(n3030), 
            .I1(GND_net), .CO(n59033));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n65957));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_CARRY add_151_7 (.CI(n58141), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n58142));
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n59031), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_19 (.CI(n58153), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n58154));
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(n78030), .I1(n1620), 
            .I2(VCC_net), .I3(n58550), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n59031), .I0(n3031), 
            .I1(VCC_net), .CO(n59032));
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [2]), 
            .O(n10_adj_5965));   // verilog/coms.v(100[12:26])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n59030), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n58549), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n58549), .I0(n1621), 
            .I1(VCC_net), .CO(n58550));
    SB_LUT4 i1_2_lut_3_lut_adj_2002 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(n66388), .I3(GND_net), .O(n26732));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_2002.LUT_INIT = 16'h9696;
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n59030), .I0(n3032), 
            .I1(GND_net), .CO(n59031));
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n58548), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n59029), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n58548), .I0(n1622), 
            .I1(VCC_net), .CO(n58549));
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n59029), .I0(n3033), 
            .I1(VCC_net), .CO(n59030));
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n58547), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n65956));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n58547), .I0(n1623), 
            .I1(VCC_net), .CO(n58548));
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n59029));
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n58546), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(n77679), .I1(n2907), 
            .I2(VCC_net), .I3(n59028), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n58546), .I0(n1624), 
            .I1(VCC_net), .CO(n58547));
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n59027), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n59027), .I0(n2908), 
            .I1(VCC_net), .CO(n59028));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n65955));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n58545), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n59026), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n58545), .I0(n1625), 
            .I1(VCC_net), .CO(n58546));
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n59026), .I0(n2909), 
            .I1(VCC_net), .CO(n59027));
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n58544), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n58140), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n58544), .I0(n1626), 
            .I1(VCC_net), .CO(n58545));
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n58543), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n59025), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n58543), .I0(n1627), 
            .I1(VCC_net), .CO(n58544));
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n58152), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_18 (.CI(n58152), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n58153));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n58151), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n58542), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n65954));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n58542), .I0(n1628), 
            .I1(VCC_net), .CO(n58543));
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n58541), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n59025), .I0(n2910), 
            .I1(VCC_net), .CO(n59026));
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n58541), .I0(n1629), 
            .I1(GND_net), .CO(n58542));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n65953));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n58540), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n59024), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n58540), .I0(n1630), 
            .I1(GND_net), .CO(n58541));
    SB_CARRY add_151_17 (.CI(n58151), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n58152));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n58150), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n58539), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n65952));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n59024), .I0(n2911), 
            .I1(VCC_net), .CO(n59025));
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n58539), .I0(n1631), 
            .I1(VCC_net), .CO(n58540));
    SB_CARRY add_151_16 (.CI(n58150), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n58151));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n58149), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n58149), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n58150));
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n58538), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n59023), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n58538), .I0(n1632), 
            .I1(GND_net), .CO(n58539));
    SB_CARRY add_151_6 (.CI(n58140), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n58141));
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n58537), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n59023), .I0(n2912), 
            .I1(VCC_net), .CO(n59024));
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n58537), .I0(n1633), 
            .I1(VCC_net), .CO(n58538));
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n59022), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n58537));
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n58137));
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n58148), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n65951));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n59022), .I0(n2913), 
            .I1(VCC_net), .CO(n59023));
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n59021), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n59021), .I0(n2914), 
            .I1(VCC_net), .CO(n59022));
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n59020), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n59020), .I0(n2915), 
            .I1(VCC_net), .CO(n59021));
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n59019), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n59019), .I0(n2916), 
            .I1(VCC_net), .CO(n59020));
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n59018), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n59018), .I0(n2917), 
            .I1(VCC_net), .CO(n59019));
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n59017), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n59017), .I0(n2918), 
            .I1(VCC_net), .CO(n59018));
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n59016), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n59016), .I0(n2919), 
            .I1(VCC_net), .CO(n59017));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n59015), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n65950));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n59015), .I0(n2920), 
            .I1(VCC_net), .CO(n59016));
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n59014), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n65949));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n59014), .I0(n2921), 
            .I1(VCC_net), .CO(n59015));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n59013), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n59013), .I0(n2922), 
            .I1(VCC_net), .CO(n59014));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n59012), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n59012), .I0(n2923), 
            .I1(VCC_net), .CO(n59013));
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n59011), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n65948));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n59011), .I0(n2924), 
            .I1(VCC_net), .CO(n59012));
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n59010), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n65947));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n65946));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n65945));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n65944));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2016 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69697), .O(n69703));
    defparam i1_4_lut_adj_2016.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2017 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69703), .O(n69709));
    defparam i1_4_lut_adj_2017.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2018 (.I0(n66388), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n66240));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_2018.LUT_INIT = 16'h9696;
    SB_LUT4 i15692_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n69709), 
            .I3(n27_adj_5865), .O(n29904));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15692_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2019 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69601), .O(n69607));
    defparam i1_4_lut_adj_2019.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2020 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69607), .O(n69613));
    defparam i1_4_lut_adj_2020.LUT_INIT = 16'hfffe;
    SB_LUT4 i15696_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n69613), 
            .I3(n27_adj_5865), .O(n29908));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15696_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2021 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n65853));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2021.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n65943));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2023 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69617), .O(n69623));
    defparam i1_4_lut_adj_2023.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2024 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69623), .O(n69629));
    defparam i1_4_lut_adj_2024.LUT_INIT = 16'hfffe;
    SB_LUT4 i15700_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n69629), 
            .I3(n27_adj_5865), .O(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15700_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2025 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69633), .O(n69639));
    defparam i1_4_lut_adj_2025.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2026 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69639), .O(n69645));
    defparam i1_4_lut_adj_2026.LUT_INIT = 16'hfffe;
    SB_LUT4 i15701_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n69645), 
            .I3(n27_adj_5865), .O(n29913));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15701_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2027 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n65856));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2027.LUT_INIT = 16'h2300;
    SB_LUT4 i62239_4_lut (.I0(n2314), .I1(n2313), .I2(n69022), .I3(n70249), 
            .O(n2346));
    defparam i62239_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_2028 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69665), .O(n69671));
    defparam i1_4_lut_adj_2028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2029 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69671), .O(n69677));
    defparam i1_4_lut_adj_2029.LUT_INIT = 16'hfffe;
    SB_LUT4 i15720_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n69677), 
            .I3(n27_adj_5865), .O(n29932));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15720_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_2030 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69649), .O(n69655));
    defparam i1_4_lut_adj_2030.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n65942));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2032 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69655), .O(n69661));
    defparam i1_4_lut_adj_2032.LUT_INIT = 16'hfffe;
    SB_LUT4 i15722_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n69661), 
            .I3(n27_adj_5865), .O(n29934));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15722_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2033 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n65861));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2033.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2034 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69585), .O(n69591));
    defparam i1_4_lut_adj_2034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2035 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69591), .O(n69597));
    defparam i1_4_lut_adj_2035.LUT_INIT = 16'hfffe;
    SB_LUT4 i15723_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n69597), 
            .I3(n27_adj_5865), .O(n29935));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15723_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15727_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n23023), .I3(GND_net), .O(n29939));   // verilog/coms.v(130[12] 305[6])
    defparam i15727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15731_3_lut (.I0(ID[0]), .I1(data_adj_6032[0]), .I2(n68385), 
            .I3(GND_net), .O(n29943));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15733_3_lut (.I0(current[0]), .I1(data_adj_6039[0]), .I2(n28097), 
            .I3(GND_net), .O(n29945));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15735_3_lut (.I0(CS_c), .I1(state_adj_6041[0]), .I2(state_adj_6041[1]), 
            .I3(GND_net), .O(n29947));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15735_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i6_4_lut_adj_2036 (.I0(n66644), .I1(\data_out_frame[13] [1]), 
            .I2(n67902), .I3(n66463), .O(n15_adj_5959));
    defparam i6_4_lut_adj_2036.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5959), .I1(n34_adj_5847), .I2(n14_adj_5960), 
            .I3(n27004), .O(n68798));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i62625_4_lut (.I0(n15_adj_5798), .I1(clk_out), .I2(state_adj_6041[0]), 
            .I3(state_adj_6041[1]), .O(n9_adj_5973));   // verilog/tli4970.v(35[10] 68[6])
    defparam i62625_4_lut.LUT_INIT = 16'hc8fc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2037 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n65865));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2037.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2038 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n65866));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2038.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2039 (.I0(n23_adj_5866), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5218), .I3(r_SM_Main_adj_6055[0]), .O(n69459));
    defparam i1_4_lut_adj_2039.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_2040 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5865), 
            .I2(n29_adj_5864), .I3(n69459), .O(n67642));
    defparam i1_4_lut_adj_2040.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15745_3_lut (.I0(b_prev_adj_5803), .I1(b_new_adj_6019[1]), 
            .I2(debounce_cnt_N_3833_adj_5804), .I3(GND_net), .O(n29957));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15745_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2041 (.I0(n2426), .I1(n2427), .I2(n2424), .I3(n2428), 
            .O(n70463));
    defparam i1_4_lut_adj_2041.LUT_INIT = 16'hfffe;
    SB_LUT4 i15746_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[1]), 
            .I2(n10_adj_5953), .I3(n25930), .O(n29958));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15746_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n65867));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 i15747_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[2]), 
            .I2(n4_adj_5792), .I3(n25888), .O(n29959));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15747_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15751_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[3]), 
            .I2(n4_adj_5792), .I3(n25930), .O(n29963));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15752_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[4]), 
            .I2(n4_adj_5793), .I3(n25888), .O(n29964));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15752_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_adj_2043 (.I0(n2425), .I1(n2422), .I2(n2423), .I3(GND_net), 
            .O(n70461));
    defparam i1_3_lut_adj_2043.LUT_INIT = 16'hfefe;
    SB_LUT4 i15753_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[5]), 
            .I2(n4_adj_5793), .I3(n25930), .O(n29965));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n65868));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n65869));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n65872));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_2047 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[4] [6]), .O(n26478));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_2047.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15754_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3163), .I3(GND_net), 
            .O(n29966));   // verilog/neopixel.v(34[12] 113[6])
    defparam i15754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15755_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[6]), 
            .I2(n44644), .I3(n25888), .O(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15755_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2048 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n65875));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2048.LUT_INIT = 16'h2300;
    SB_LUT4 mux_3812_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5736), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15756_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_6032[7]), 
            .I2(n44644), .I3(n25930), .O(n29968));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15756_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7583_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n21152));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i7583_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8841_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i8841_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51114_3_lut (.I0(n4_adj_5971), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n66892));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i51114_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2049 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n29286));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2049.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2050 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n65876));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2050.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n65877));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_2052 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n69276));
    defparam i3_4_lut_adj_2052.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n65878));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15772_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29984));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2054 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n65879));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2054.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n65880));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1178_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5933));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59172_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n75007));   // verilog/uart_rx.v(119[17:57])
    defparam i59172_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i2_3_lut_4_lut_adj_2056 (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5963));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i2_3_lut_4_lut_adj_2056.LUT_INIT = 16'h080c;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n44439), .O(n24_adj_5957));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i31227_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n45307));
    defparam i31227_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n65874));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2058 (.I0(n2420), .I1(n2421), .I2(n70461), .I3(n70463), 
            .O(n70469));
    defparam i1_4_lut_adj_2058.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n65881));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2060 (.I0(n2429), .I1(n45307), .I2(n2430), .I3(n2431), 
            .O(n67822));
    defparam i1_4_lut_adj_2060.LUT_INIT = 16'ha080;
    SB_LUT4 i30206_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n23023), .I3(GND_net), .O(n29988));
    defparam i30206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15777_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n23023), .I3(GND_net), .O(n29989));   // verilog/coms.v(130[12] 305[6])
    defparam i15777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2061 (.I0(n2418), .I1(n2419), .I2(n67822), .I3(n70469), 
            .O(n70475));
    defparam i1_4_lut_adj_2061.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5809));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16558_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30770));   // verilog/coms.v(130[12] 305[6])
    defparam i16558_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2062 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n70475), 
            .O(n70481));
    defparam i1_4_lut_adj_2062.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n65882));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i62131_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n70481), 
            .O(n2445));
    defparam i62131_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2064 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n65883));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2064.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n65884));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2066 (.I0(n2528), .I1(n2523), .I2(n2527), .I3(GND_net), 
            .O(n70175));
    defparam i1_3_lut_adj_2066.LUT_INIT = 16'hfefe;
    SB_LUT4 i51116_3_lut (.I0(n3), .I1(n7755), .I2(n66893), .I3(GND_net), 
            .O(n66894));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31297_4_lut (.I0(n950), .I1(n2531), .I2(n2532), .I3(n2533), 
            .O(n45377));
    defparam i31297_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i51117_3_lut (.I0(encoder0_position[29]), .I1(n66894), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2067 (.I0(n2518), .I1(n2525), .I2(n2521), .I3(n2522), 
            .O(n70189));
    defparam i1_4_lut_adj_2067.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n65885));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n65886));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2070 (.I0(n70189), .I1(n2529), .I2(n45377), .I3(n2530), 
            .O(n70191));
    defparam i1_4_lut_adj_2070.LUT_INIT = 16'heaaa;
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2071 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n70191), 
            .O(n70197));
    defparam i1_4_lut_adj_2071.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2072 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n65887));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2072.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n65888));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    SB_LUT4 i16554_3_lut_4_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30766));   // verilog/coms.v(130[12] 305[6])
    defparam i16554_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2074 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n65889));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2074.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2075 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n65890));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2075.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2076 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n65891));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2076.LUT_INIT = 16'h2300;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n28115), .O(n61786));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2077 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n65892));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2077.LUT_INIT = 16'h2300;
    SB_LUT4 i59181_3_lut_4_lut (.I0(r_Clock_Count_adj_6056[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_6056[2]), .O(n75016));   // verilog/uart_tx.v(117[17:57])
    defparam i59181_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1181_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_6056[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5926));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i11_2_lut (.I0(pwm_setpoint[19]), .I1(pwm_counter[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/pwm.v(11[19:30])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_2_lut_adj_2078 (.I0(pwm_setpoint[20]), .I1(pwm_counter[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(11[19:30])
    defparam i10_2_lut_adj_2078.LUT_INIT = 16'h6666;
    SB_LUT4 i61896_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n44439), .I3(GND_net), .O(n28128));
    defparam i61896_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i1_4_lut_adj_2079 (.I0(n2520), .I1(n70175), .I2(n2524), .I3(n2526), 
            .O(n70179));
    defparam i1_4_lut_adj_2079.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2080 (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n70197), 
            .O(n69064));
    defparam i1_4_lut_adj_2080.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5849));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62191_4_lut (.I0(n2517), .I1(n69064), .I2(n2519), .I3(n70179), 
            .O(n2544));
    defparam i62191_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i59013_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n74462));
    defparam i59013_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5849), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2081 (.I0(n2626), .I1(n2628), .I2(GND_net), .I3(GND_net), 
            .O(n70519));
    defparam i1_2_lut_adj_2081.LUT_INIT = 16'heeee;
    SB_LUT4 i59275_2_lut (.I0(n78900), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74617));
    defparam i59275_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i30460_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n44439), .I3(GND_net), .O(n44534));
    defparam i30460_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2082 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n65893));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2082.LUT_INIT = 16'h2300;
    SB_LUT4 i23197_3_lut_4_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30053));
    defparam i23197_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15778_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n23023), .I3(GND_net), .O(n29990));   // verilog/coms.v(130[12] 305[6])
    defparam i15778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55856_3_lut (.I0(n4908), .I1(duty[20]), .I2(n11849), .I3(GND_net), 
            .O(n71691));
    defparam i55856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55858_3_lut (.I0(n71691), .I1(n71686), .I2(n11847), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i55858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55853_3_lut (.I0(n4907), .I1(duty[21]), .I2(n11849), .I3(GND_net), 
            .O(n71688));
    defparam i55853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16523_3_lut_4_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30735));   // verilog/coms.v(130[12] 305[6])
    defparam i16523_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i55855_3_lut (.I0(n71688), .I1(n71686), .I2(n11847), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i55855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55851_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11849), 
            .I3(GND_net), .O(n71686));
    defparam i55851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55850_3_lut (.I0(n4906), .I1(duty[22]), .I2(n11849), .I3(GND_net), 
            .O(n71685));
    defparam i55850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20507_3_lut_4_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30734));
    defparam i20507_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i55852_3_lut (.I0(n71685), .I1(n71686), .I2(n11847), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i55852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7290_3_lut (.I0(n4905), .I1(current[15]), .I2(n11847), .I3(GND_net), 
            .O(n21156));
    defparam i7290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7291_3_lut (.I0(n21156), .I1(duty[23]), .I2(n11849), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5718));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2083 (.I0(n2622), .I1(n2625), .I2(n2623), .I3(n2624), 
            .O(n70527));
    defparam i1_4_lut_adj_2083.LUT_INIT = 16'hfffe;
    SB_LUT4 i15779_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n23023), .I3(GND_net), .O(n29991));   // verilog/coms.v(130[12] 305[6])
    defparam i15779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15780_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n23023), .I3(GND_net), .O(n29992));   // verilog/coms.v(130[12] 305[6])
    defparam i15780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15840_3_lut_4_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30052));   // verilog/coms.v(130[12] 305[6])
    defparam i15840_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15839_3_lut_4_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30051));   // verilog/coms.v(130[12] 305[6])
    defparam i15839_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22999_3_lut_4_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30050));
    defparam i22999_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16519_3_lut_4_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30731));   // verilog/coms.v(130[12] 305[6])
    defparam i16519_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i30205_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n23023), .I3(GND_net), .O(n29993));
    defparam i30205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23725_3_lut_4_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30730));
    defparam i23725_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i23462_3_lut (.I0(n32_adj_5871), .I1(pwm_counter[16]), .I2(pwm_setpoint[16]), 
            .I3(GND_net), .O(n34_adj_5872));   // verilog/pwm.v(11[19:30])
    defparam i23462_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30196_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n23023), .I3(GND_net), .O(n29994));
    defparam i30196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15783_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n23023), .I3(GND_net), .O(n29995));   // verilog/coms.v(130[12] 305[6])
    defparam i15783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15784_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n23023), .I3(GND_net), .O(n29996));   // verilog/coms.v(130[12] 305[6])
    defparam i15784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15785_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n23023), .I3(GND_net), .O(n29997));   // verilog/coms.v(130[12] 305[6])
    defparam i15785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15786_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n23023), .I3(GND_net), .O(n29998));   // verilog/coms.v(130[12] 305[6])
    defparam i15786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5740), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15787_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n23023), .I3(GND_net), .O(n29999));   // verilog/coms.v(130[12] 305[6])
    defparam i15787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15788_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n23023), .I3(GND_net), .O(n30000));   // verilog/coms.v(130[12] 305[6])
    defparam i15788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16516_3_lut_4_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30728));   // verilog/coms.v(130[12] 305[6])
    defparam i16516_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2084 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n65894));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2084.LUT_INIT = 16'h2300;
    SB_LUT4 i16513_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(reset), .I3(n76), .O(n30725));   // verilog/coms.v(130[12] 305[6])
    defparam i16513_3_lut_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2085 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n65895));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2085.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2086 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n65896));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2086.LUT_INIT = 16'h2300;
    SB_LUT4 i15837_3_lut_4_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30049));   // verilog/coms.v(130[12] 305[6])
    defparam i15837_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15836_3_lut_4_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30048));   // verilog/coms.v(130[12] 305[6])
    defparam i15836_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(n76), .I2(GND_net), .I3(GND_net), 
            .O(n28713));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i59151_2_lut (.I0(n78804), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74616));
    defparam i59151_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15835_3_lut_4_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30047));   // verilog/coms.v(130[12] 305[6])
    defparam i15835_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2087 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n65897));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2087.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5810));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5811));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16511_3_lut_4_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30723));   // verilog/coms.v(130[12] 305[6])
    defparam i16511_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i30352_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i30352_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2088 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n65898));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2088.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2089 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n65899));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2089.LUT_INIT = 16'h2300;
    SB_LUT4 i30473_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i30473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16509_3_lut_4_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30721));   // verilog/coms.v(130[12] 305[6])
    defparam i16509_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_243_i22_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i24_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16508_3_lut_4_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30720));   // verilog/coms.v(130[12] 305[6])
    defparam i16508_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2090 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n65900));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2090.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_2091 (.I0(n35278), .I1(control_mode[0]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5766));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_2091.LUT_INIT = 16'heeee;
    SB_LUT4 mux_243_i1_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[0]), .I3(encoder0_position_scaled[0]), 
            .O(motor_state[0]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2092 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n65901));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2092.LUT_INIT = 16'h2300;
    SB_LUT4 i15789_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n23023), .I3(GND_net), .O(n30001));   // verilog/coms.v(130[12] 305[6])
    defparam i15789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15794_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n30006));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i9_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[8]), .I3(encoder0_position_scaled[8]), 
            .O(motor_state[8]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i23_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i19_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2093 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n65902));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2093.LUT_INIT = 16'h2300;
    SB_LUT4 mux_243_i10_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i21_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5754), .I3(n15_adj_5825), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5788));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_243_i20_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2094 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n65903));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2094.LUT_INIT = 16'h2300;
    SB_LUT4 mux_243_i18_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i17_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i16485_3_lut_4_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30697));   // verilog/coms.v(130[12] 305[6])
    defparam i16485_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1779(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .n30010(n30010), 
            .n1742(n1742), .n30006(n30006), .a_prev(a_prev), .n29984(n29984), 
            .b_prev(b_prev), .position_31__N_3836(position_31__N_3836), 
            .n1744(n1744), .\encoder0_position[30] (encoder0_position[30]), 
            .\encoder0_position[29] (encoder0_position[29]), .\encoder0_position[28] (encoder0_position[28]), 
            .\encoder0_position[27] (encoder0_position[27]), .\encoder0_position[26] (encoder0_position[26]), 
            .\encoder0_position[25] (encoder0_position[25]), .\encoder0_position[24] (encoder0_position[24]), 
            .\encoder0_position[23] (encoder0_position[23]), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), .GND_net(GND_net), 
            .VCC_net(VCC_net), .debounce_cnt_N_3833(debounce_cnt_N_3833)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5784));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15799_3_lut (.I0(a_prev_adj_5802), .I1(a_new_adj_6018[1]), 
            .I2(debounce_cnt_N_3833_adj_5804), .I3(GND_net), .O(n30011));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2095 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n65904));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2095.LUT_INIT = 16'h2300;
    SB_LUT4 mux_243_i8_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[7]), .I3(encoder0_position_scaled[7]), 
            .O(motor_state[7]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5786));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_243_i16_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i6_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[5]), .I3(encoder0_position_scaled[5]), 
            .O(motor_state[5]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16467_3_lut_4_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30679));   // verilog/coms.v(130[12] 305[6])
    defparam i16467_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_243_i15_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i13_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i7_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[6]), .I3(encoder0_position_scaled[6]), 
            .O(motor_state[6]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i14_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i11_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i5_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[4]), .I3(encoder0_position_scaled[4]), 
            .O(motor_state[4]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i16465_3_lut_4_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30677));   // verilog/coms.v(130[12] 305[6])
    defparam i16465_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2096 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n65905));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2096.LUT_INIT = 16'h2300;
    SB_LUT4 mux_243_i12_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i4_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[3]), .I3(encoder0_position_scaled[3]), 
            .O(motor_state[3]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i2_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[1]), .I3(encoder0_position_scaled[1]), 
            .O(motor_state[1]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i3_3_lut_4_lut (.I0(control_mode[1]), .I1(n25_adj_5766), 
            .I2(motor_state_23__N_91[2]), .I3(encoder0_position_scaled[2]), 
            .O(motor_state[2]));   // verilog/coms.v(130[12] 305[6])
    defparam mux_243_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30363_3_lut_4_lut (.I0(n35278), .I1(control_mode[0]), .I2(control_update), 
            .I3(control_mode[1]), .O(n28074));   // verilog/coms.v(130[12] 305[6])
    defparam i30363_3_lut_4_lut.LUT_INIT = 16'hb0f0;
    SB_LUT4 i1_4_lut_adj_2097 (.I0(n2627), .I1(n70519), .I2(n2620), .I3(n2621), 
            .O(n70529));
    defparam i1_4_lut_adj_2097.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31223_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n45303));
    defparam i31223_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_2098 (.I0(n35278), .I1(control_mode[0]), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_5754));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_2098.LUT_INIT = 16'hfbfb;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n71810), .I3(n71808), .O(n7_adj_5952));   // verilog/coms.v(105[12:33])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16451_3_lut_4_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30663));   // verilog/coms.v(130[12] 305[6])
    defparam i16451_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n71789), .I3(n71787), .O(n7_adj_5951));   // verilog/coms.v(105[12:33])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n71786), .I3(n71784), .O(n7_adj_5950));   // verilog/coms.v(105[12:33])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2099 (.I0(n2618), .I1(n70529), .I2(n2619), .I3(n70527), 
            .O(n70535));
    defparam i1_4_lut_adj_2099.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n71771), .I3(n71769), .O(n7_adj_5796));   // verilog/coms.v(105[12:33])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n71768), .I3(n71766), .O(n7_adj_5949));   // verilog/coms.v(105[12:33])
    defparam i10_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2100 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n65906));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2100.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2101 (.I0(n2629), .I1(n45303), .I2(n2630), .I3(n2631), 
            .O(n67837));
    defparam i1_4_lut_adj_2101.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2102 (.I0(n2616), .I1(n2617), .I2(n67837), .I3(n70535), 
            .O(n70541));
    defparam i1_4_lut_adj_2102.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2103 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n65907));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2103.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2104 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n65908));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2104.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2105 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n65909));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2105.LUT_INIT = 16'h2300;
    SB_LUT4 i59208_2_lut_4_lut (.I0(duty[6]), .I1(n304), .I2(duty[5]), 
            .I3(n305), .O(n75043));
    defparam i59208_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i59202_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n75037));
    defparam i59202_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2106 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n70541), 
            .O(n70547));
    defparam i1_4_lut_adj_2106.LUT_INIT = 16'hfffe;
    SB_LUT4 i62160_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n70547), 
            .O(n2643));
    defparam i62160_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2107 (.I0(n2723), .I1(n2724), .I2(n2727), .I3(n2728), 
            .O(n70043));
    defparam i1_4_lut_adj_2107.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2108 (.I0(n2721), .I1(n2725), .I2(n2726), .I3(n2722), 
            .O(n70045));
    defparam i1_4_lut_adj_2108.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_2109 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n70913));
    defparam i1_2_lut_adj_2109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_2110 (.I0(n66555), .I1(\data_in_frame[12] [4]), 
            .I2(n70913), .I3(\data_in_frame[17] [5]), .O(n70919));
    defparam i1_4_lut_adj_2110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2111 (.I0(n66660), .I1(n66842), .I2(n70919), 
            .I3(n66244), .O(n70925));
    defparam i1_4_lut_adj_2111.LUT_INIT = 16'h6996;
    SB_LUT4 mux_3812_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5741), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2112 (.I0(n27201), .I1(n66788), .I2(n66590), 
            .I3(n70925), .O(n61349));
    defparam i1_4_lut_adj_2112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2113 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n65910));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2113.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2114 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n29249));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2114.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31293_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n45373));
    defparam i31293_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16419_3_lut_4_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30631));   // verilog/coms.v(130[12] 305[6])
    defparam i16419_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16417_3_lut_4_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30629));   // verilog/coms.v(130[12] 305[6])
    defparam i16417_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_2115 (.I0(\data_in_frame[14] [5]), .I1(n26873), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5756));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_2115.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_2116 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [4]), 
            .I2(n27241), .I3(n6_adj_5756), .O(n60656));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_2116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_2117 (.I0(n2719), .I1(n2720), .I2(n70045), .I3(n70043), 
            .O(n70051));
    defparam i1_4_lut_adj_2117.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_2_lut (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5753));   // verilog/coms.v(99[12:25])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16416_3_lut_4_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30628));   // verilog/coms.v(130[12] 305[6])
    defparam i16416_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2118 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n65911));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2118.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2119 (.I0(n2729), .I1(n2730), .I2(GND_net), .I3(GND_net), 
            .O(n70565));
    defparam i1_2_lut_adj_2119.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16412_3_lut_4_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30624));   // verilog/coms.v(130[12] 305[6])
    defparam i16412_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2120 (.I0(n2718), .I1(n70565), .I2(n70051), .I3(n45373), 
            .O(n70055));
    defparam i1_4_lut_adj_2120.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16410_3_lut_4_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30622));   // verilog/coms.v(130[12] 305[6])
    defparam i16410_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_adj_2121 (.I0(hall1), .I1(hall2), .I2(n21152), 
            .I3(GND_net), .O(n4_adj_5971));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_2121.LUT_INIT = 16'hf2f2;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5772));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59238_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n75073));
    defparam i59238_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_2122 (.I0(n2715), .I1(n2716), .I2(n2717), .I3(n70055), 
            .O(n70061));
    defparam i1_4_lut_adj_2122.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5770));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2123 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n65912));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2123.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2124 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n70061), 
            .O(n70067));
    defparam i1_4_lut_adj_2124.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i62534_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n70067), 
            .O(n2742));
    defparam i62534_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2125 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n65913));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2125.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15834_3_lut_4_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30046));   // verilog/coms.v(130[12] 305[6])
    defparam i15834_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2126 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n65914));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2126.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i21_3_lut (.I0(encoder0_position[20]), .I1(n12_adj_5743), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n937));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15833_3_lut_4_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30045));   // verilog/coms.v(130[12] 305[6])
    defparam i15833_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15832_3_lut_4_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30044));   // verilog/coms.v(130[12] 305[6])
    defparam i15832_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15831_3_lut_4_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30043));   // verilog/coms.v(130[12] 305[6])
    defparam i15831_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15830_3_lut_4_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30042));   // verilog/coms.v(130[12] 305[6])
    defparam i15830_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15829_3_lut_4_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30041));   // verilog/coms.v(130[12] 305[6])
    defparam i15829_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15828_3_lut_4_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30040));   // verilog/coms.v(130[12] 305[6])
    defparam i15828_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15827_3_lut_4_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30039));   // verilog/coms.v(130[12] 305[6])
    defparam i15827_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i6661_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6661_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6659_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6659_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2127 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n65873));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2127.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(\data_out_frame[19] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[0]), .O(n78639));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2128 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n66039));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2128.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2129 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n66038));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2129.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2130 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n66037));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2130.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2131 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n66036));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2131.LUT_INIT = 16'h2300;
    SB_LUT4 n78639_bdd_4_lut (.I0(n78639), .I1(\data_out_frame[22] [0]), 
            .I2(\data_out_frame[18] [0]), .I3(byte_transmit_counter[0]), 
            .O(n78642));
    defparam n78639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2132 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n66035));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2132.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2133 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n66034));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2133.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2134 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n65863));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2134.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2135 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n65860));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2135.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2136 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n66033));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2136.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_4_lut_adj_2137 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2819), .O(n25_adj_5956));   // verilog/TinyFPGA_B.v(377[7:11])
    defparam i1_4_lut_4_lut_adj_2137.LUT_INIT = 16'h5450;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5863), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62652_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5976));
    defparam i62652_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_2138 (.I0(\data_in_frame[14] [4]), .I1(n66625), 
            .I2(\data_in_frame[12] [3]), .I3(n61123), .O(n26758));
    defparam i3_4_lut_adj_2138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2139 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n66032));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2139.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2140 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n66031));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2140.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2141 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n65870));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2141.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2142 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n65864));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2142.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2143 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n66030));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2143.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2144 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n66029));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2144.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2145 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n66028));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2145.LUT_INIT = 16'h2300;
    SB_LUT4 i60943_3_lut (.I0(n78768), .I1(n78498), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76778));
    defparam i60943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60944_4_lut (.I0(n76778), .I1(n78834), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n76779));
    defparam i60944_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i55924_3_lut (.I0(n78576), .I1(n76779), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i55924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2146 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n66027));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2146.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31241_3_lut (.I0(n953), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n45321));
    defparam i31241_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1956_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n44439), .O(n6901));   // verilog/TinyFPGA_B.v(362[5] 388[12])
    defparam i1956_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i1_4_lut_adj_2147 (.I0(n2829), .I1(n45321), .I2(n2830), .I3(n2831), 
            .O(n67847));
    defparam i1_4_lut_adj_2147.LUT_INIT = 16'ha080;
    SB_LUT4 mux_3812_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5742), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n938));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2148 (.I0(n2817), .I1(n67847), .I2(n2821), .I3(n2825), 
            .O(n68695));
    defparam i1_4_lut_adj_2148.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2149 (.I0(n2813), .I1(n68695), .I2(n2816), .I3(n2828), 
            .O(n70507));
    defparam i1_4_lut_adj_2149.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2150 (.I0(n2814), .I1(n2812), .I2(n2815), .I3(n2824), 
            .O(n68771));
    defparam i1_4_lut_adj_2150.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2151 (.I0(n2826), .I1(n2822), .I2(n2827), .I3(n2823), 
            .O(n70497));
    defparam i1_4_lut_adj_2151.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2152 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n66026));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2152.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2153 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n66025));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2153.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2154 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n66024));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2154.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2155 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n66023));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2155.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2156 (.I0(n2810), .I1(n68771), .I2(n2811), .I3(n70507), 
            .O(n70513));
    defparam i1_4_lut_adj_2156.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2157 (.I0(n2818), .I1(n70497), .I2(n2819_adj_5867), 
            .I3(n2820), .O(n70501));
    defparam i1_4_lut_adj_2157.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62586_4_lut (.I0(n2808), .I1(n70501), .I2(n70513), .I3(n2809), 
            .O(n2841));
    defparam i62586_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2158 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n66022));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2158.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62761 (.I0(byte_transmit_counter[1]), 
            .I1(n71754), .I2(n71755), .I3(byte_transmit_counter[2]), .O(n78615));
    defparam byte_transmit_counter_1__bdd_4_lut_62761.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n78615_bdd_4_lut (.I0(n78615), .I1(n71908), .I2(n71907), .I3(byte_transmit_counter[2]), 
            .O(n78618));
    defparam n78615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_2159 (.I0(dti_counter[6]), .I1(dti_counter[4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5833));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut_adj_2159.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2160 (.I0(dti_counter[0]), .I1(dti_counter[3]), 
            .I2(n6_adj_5833), .I3(dti_counter[2]), .O(n6_adj_5832));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i1_4_lut_adj_2160.LUT_INIT = 16'hfffe;
    SB_LUT4 i15229_2_lut_3_lut (.I0(n23186), .I1(dti), .I2(n15_adj_5791), 
            .I3(GND_net), .O(n29436));
    defparam i15229_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i4_4_lut_adj_2161 (.I0(dti_counter[1]), .I1(dti_counter[5]), 
            .I2(dti_counter[7]), .I3(n6_adj_5832), .O(n23186));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i4_4_lut_adj_2161.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_2162 (.I0(n23186), .I1(dti), .I2(n15_adj_5791), 
            .I3(GND_net), .O(n28172));
    defparam i1_2_lut_3_lut_adj_2162.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_4_lut_adj_2163 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5972));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2163.LUT_INIT = 16'h7bde;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2164 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n66021));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2164.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2165 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n66020));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2165.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819_adj_5867));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15881_3_lut_4_lut (.I0(deadband[1]), .I1(\data_in_frame[16] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30093));   // verilog/coms.v(130[12] 305[6])
    defparam i15881_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15880_3_lut_4_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30092));   // verilog/coms.v(130[12] 305[6])
    defparam i15880_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_3812_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5744), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n936));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5857));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5857), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.VCC_net(VCC_net), .GND_net(GND_net), .clk16MHz(clk16MHz), 
            .n5(n5_adj_5797), .n5_adj_29(n5_adj_5826), .n5_adj_30(n5_adj_5814), 
            .\state[0] (state_adj_6041[0]), .\state[1] (state_adj_6041[1]), 
            .state_7__N_4319(state_7__N_4319), .n44573(n44573), .clk_out(clk_out), 
            .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .n15(n15_adj_5798), .n30117(n30117), 
            .\data[15] (data_adj_6039[15]), .n30116(n30116), .\data[12] (data_adj_6039[12]), 
            .n30115(n30115), .\data[11] (data_adj_6039[11]), .n30114(n30114), 
            .\data[10] (data_adj_6039[10]), .n30113(n30113), .\data[9] (data_adj_6039[9]), 
            .n30112(n30112), .\data[8] (data_adj_6039[8]), .n30111(n30111), 
            .\data[7] (data_adj_6039[7]), .n30110(n30110), .\data[6] (data_adj_6039[6]), 
            .n30109(n30109), .\data[5] (data_adj_6039[5]), .n30108(n30108), 
            .\data[4] (data_adj_6039[4]), .n30107(n30107), .\data[3] (data_adj_6039[3]), 
            .n30106(n30106), .\data[2] (data_adj_6039[2]), .n30105(n30105), 
            .\data[1] (data_adj_6039[1]), .n25893(n25893), .n11(n11_adj_5799), 
            .n25910(n25910), .n25867(n25867), .n9(n9_adj_5973), .n29947(n29947), 
            .n29945(n29945), .\current[0] (current[0]), .n30765(n30765), 
            .\data[0] (data_adj_6039[0]), .n30675(n30675), .\current[1] (current[1]), 
            .n30674(n30674), .\current[2] (current[2]), .n30673(n30673), 
            .\current[3] (current[3]), .n30672(n30672), .\current[4] (current[4]), 
            .n30671(n30671), .\current[5] (current[5]), .n30670(n30670), 
            .\current[6] (current[6]), .n30669(n30669), .\current[7] (current[7]), 
            .n30668(n30668), .\current[8] (current[8]), .n30667(n30667), 
            .\current[9] (current[9]), .n30666(n30666), .\current[10] (current[10]), 
            .n30665(n30665), .\current[11] (current[11]), .n28097(n28097), 
            .\current[15] (current[15]), .n25883(n25883)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(405[11] 411[4])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2166 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n66019));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2166.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_2167 (.I0(commutation_state[0]), .I1(n4_adj_5972), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5791));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i2_3_lut_adj_2167.LUT_INIT = 16'hdede;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1181_i15_2_lut (.I0(r_Clock_Count_adj_6056[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5931));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i9_2_lut (.I0(r_Clock_Count_adj_6056[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5928));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i13_2_lut (.I0(r_Clock_Count_adj_6056[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5930));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i11_2_lut (.I0(r_Clock_Count_adj_6056[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5929));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2168 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n66018));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2168.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1181_i4_4_lut (.I0(r_Clock_Count_adj_6056[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_6056[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5925));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i60781_3_lut (.I0(n4_adj_5925), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5929), 
            .I3(GND_net), .O(n76616));   // verilog/uart_tx.v(117[17:57])
    defparam i60781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i60782_3_lut (.I0(n76616), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5930), 
            .I3(GND_net), .O(n76617));   // verilog/uart_tx.v(117[17:57])
    defparam i60782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60176_4_lut (.I0(n13_adj_5930), .I1(n11_adj_5929), .I2(n9_adj_5928), 
            .I3(n75016), .O(n76011));
    defparam i60176_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1181_i8_3_lut (.I0(n6_adj_5926), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5928), .I3(GND_net), .O(n8_adj_5927));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5748), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n731));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60056_3_lut (.I0(n76617), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5931), 
            .I3(GND_net), .O(n75891));   // verilog/uart_tx.v(117[17:57])
    defparam i60056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61089_4_lut (.I0(n75891), .I1(n8_adj_5927), .I2(n15_adj_5931), 
            .I3(n76011), .O(n76924));   // verilog/uart_tx.v(117[17:57])
    defparam i61089_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61090_3_lut (.I0(n76924), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_6056[8]), 
            .I3(GND_net), .O(n5218));   // verilog/uart_tx.v(117[17:57])
    defparam i61090_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_2169 (.I0(n23_adj_5866), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5218), .I3(GND_net), .O(n69425));
    defparam i1_3_lut_adj_2169.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_2170 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5865), 
            .I2(n29_adj_5864), .I3(n69425), .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut_adj_2170.LUT_INIT = 16'hfffe;
    SB_LUT4 i51217_2_lut (.I0(r_SM_Main_adj_6055[2]), .I1(r_SM_Main_adj_6055[0]), 
            .I2(GND_net), .I3(GND_net), .O(n67002));
    defparam i51217_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_2171 (.I0(n4_adj_5750), .I1(n5), .I2(n731), .I3(n6_adj_5749), 
            .O(n5_adj_5958));
    defparam i1_4_lut_adj_2171.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_2172 (.I0(n3), .I1(n2_adj_5751), .I2(n5_adj_5958), 
            .I3(GND_net), .O(n66893));
    defparam i1_3_lut_adj_2172.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_2173 (.I0(o_Rx_DV_N_3488[12]), .I1(n5215), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n69006), .O(n69517));
    defparam i1_4_lut_adj_2173.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_2174 (.I0(o_Rx_DV_N_3488[24]), .I1(n29_adj_5864), 
            .I2(n23_adj_5866), .I3(n69517), .O(n69523));
    defparam i1_4_lut_adj_2174.LUT_INIT = 16'hfffe;
    SB_LUT4 i51124_3_lut (.I0(n7_adj_5748), .I1(n7759), .I2(n66893), .I3(GND_net), 
            .O(n66902));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51124_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .n1786(n1786), 
            .GND_net(GND_net), .n1788(n1788), .n1790(n1790), .n1792(n1792), 
            .n1794(n1794), .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .\encoder1_position[3] (encoder1_position[3]), 
            .\encoder1_position[2] (encoder1_position[2]), .\encoder1_position[1] (encoder1_position[1]), 
            .\encoder1_position[0] (encoder1_position[0]), .VCC_net(VCC_net), 
            .n30011(n30011), .a_prev(a_prev_adj_5802), .n29957(n29957), 
            .b_prev(b_prev_adj_5803), .n29956(n29956), .n1784(n1784), 
            .position_31__N_3836(position_31__N_3836_adj_5805), .\a_new[1] (a_new_adj_6018[1]), 
            .\b_new[1] (b_new_adj_6019[1]), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5804)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2175 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n65974));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2175.LUT_INIT = 16'h2300;
    SB_LUT4 i16265_4_lut_4_lut (.I0(n28192), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30477));   // verilog/neopixel.v(34[12] 113[6])
    defparam i16265_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i9_2_lut_adj_2176 (.I0(n291), .I1(n239), .I2(GND_net), .I3(GND_net), 
            .O(n37_adj_5881));
    defparam i9_2_lut_adj_2176.LUT_INIT = 16'h6666;
    SB_LUT4 i15879_3_lut_4_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30091));   // verilog/coms.v(130[12] 305[6])
    defparam i15879_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i51125_3_lut (.I0(encoder0_position[25]), .I1(n66902), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam i51125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21614_3_lut_4_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30090));
    defparam i21614_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15_2_lut (.I0(n299_adj_5795), .I1(n247), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_5880));
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2177 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n66017));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2177.LUT_INIT = 16'h2300;
    SB_LUT4 i15877_3_lut_4_lut (.I0(deadband[5]), .I1(\data_in_frame[16] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30089));   // verilog/coms.v(130[12] 305[6])
    defparam i15877_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2178 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n66016));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2178.LUT_INIT = 16'h2300;
    SB_LUT4 i43992_2_lut_3_lut_4_lut (.I0(n37146), .I1(Ki[0]), .I2(n339), 
            .I3(Ki[1]), .O(n20493));
    defparam i43992_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i43994_2_lut_3_lut_4_lut (.I0(n37146), .I1(Ki[0]), .I2(n339), 
            .I3(Ki[1]), .O(n58049));
    defparam i43994_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15876_3_lut_4_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30088));   // verilog/coms.v(130[12] 305[6])
    defparam i15876_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15875_3_lut_4_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30087));   // verilog/coms.v(130[12] 305[6])
    defparam i15875_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i43829_3_lut_4_lut (.I0(n37336), .I1(Ki[3]), .I2(n4), .I3(n20465), 
            .O(n6));
    defparam i43829_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut (.I0(n37336), .I1(Ki[3]), .I2(n4), .I3(n20465), 
            .O(n20419));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_2179 (.I0(n37336), .I1(Ki[2]), .I2(n57846), 
            .I3(n20466), .O(n20420));
    defparam i1_3_lut_4_lut_adj_2179.LUT_INIT = 16'h8778;
    SB_LUT4 i43821_3_lut_4_lut (.I0(n37336), .I1(Ki[2]), .I2(n57846), 
            .I3(n20466), .O(n4));
    defparam i43821_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i15874_3_lut_4_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30086));   // verilog/coms.v(130[12] 305[6])
    defparam i15874_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15873_3_lut_4_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30085));   // verilog/coms.v(130[12] 305[6])
    defparam i15873_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2180 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n66015));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2180.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_62775 (.I0(byte_transmit_counter[2]), 
            .I1(n71888), .I2(n71912), .I3(byte_transmit_counter[3]), .O(n78573));
    defparam byte_transmit_counter_2__bdd_4_lut_62775.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5853));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i62400_2_lut (.I0(n23186), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i62400_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5853), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15872_3_lut_4_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30084));   // verilog/coms.v(130[12] 305[6])
    defparam i15872_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n78573_bdd_4_lut (.I0(n78573), .I1(n71764), .I2(n71763), .I3(byte_transmit_counter[3]), 
            .O(n78576));
    defparam n78573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15871_3_lut_4_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30083));   // verilog/coms.v(130[12] 305[6])
    defparam i15871_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_63018 (.I0(n11849), .I1(current[15]), .I2(duty[22]), 
            .I3(n11847), .O(n78567));
    defparam n11849_bdd_4_lut_63018.LUT_INIT = 16'he4aa;
    SB_LUT4 i21995_3_lut_4_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30082));
    defparam i21995_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2181 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n66014));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2181.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15869_3_lut_4_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30081));   // verilog/coms.v(130[12] 305[6])
    defparam i15869_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15868_3_lut_4_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30080));   // verilog/coms.v(130[12] 305[6])
    defparam i15868_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n78567_bdd_4_lut (.I0(n78567), .I1(duty[19]), .I2(n4909), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[19]));
    defparam n78567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2182 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n66013));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2182.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15867_3_lut_4_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30079));   // verilog/coms.v(130[12] 305[6])
    defparam i15867_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15866_3_lut_4_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30078));   // verilog/coms.v(130[12] 305[6])
    defparam i15866_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.\data_out_frame[13] ({\data_out_frame[13] }), 
         .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), .setpoint({setpoint}), 
         .VCC_net(VCC_net), .\data_in_frame[8] ({\data_in_frame[8] }), .clk16MHz(clk16MHz), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .GND_net(GND_net), 
         .n2872(n2872), .\data_out_frame[8] ({\data_out_frame[8] }), .n66000(n66000), 
         .n65999(n65999), .byte_transmit_counter({Open_4, Open_5, Open_6, 
         byte_transmit_counter[4:0]}), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n78804(n78804), 
         .\data_out_frame[1][1] (\data_out_frame[1] [1]), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n71810(n71810), .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .n71808(n71808), .rx_data({rx_data}), .n7(n7_adj_5975), .\data_in_frame[2] ({\data_in_frame[2] [7], 
         Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, Open_13}), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_in_frame[16] ({\data_in_frame[16] }), .n28715(n28715), .n65854(n65854), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .Kp_23__N_1748(Kp_23__N_1748), 
         .reset(reset), .n8(n8_adj_5845), .n65998(n65998), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n65997(n65997), .n66003(n66003), .n65996(n65996), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .n66040(n66040), .n65995(n65995), .n65994(n65994), .n65993(n65993), 
         .n65992(n65992), .n65991(n65991), .n65990(n65990), .n65989(n65989), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .n65855(n65855), 
         .n65988(n65988), .n65987(n65987), .n65986(n65986), .n65985(n65985), 
         .n65984(n65984), .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), 
         .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .n65983(n65983), .n65982(n65982), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n65981(n65981), 
         .n65980(n65980), .n65979(n65979), .n65978(n65978), .n65977(n65977), 
         .n65976(n65976), .n65975(n65975), .n65871(n65871), .n65973(n65973), 
         .n65972(n65972), .n65971(n65971), .n65970(n65970), .n65969(n65969), 
         .n65968(n65968), .\data_in_frame[1][0] (\data_in_frame[1] [0]), 
         .encoder0_position({encoder0_position[23:0]}), .n65967(n65967), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .n65966(n65966), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n71801(n71801), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .n71799(n71799), 
         .n78768(n78768), .n65965(n65965), .\data_in_frame[0][0] (\data_in_frame[0] [0]), 
         .\data_in_frame[0][1] (\data_in_frame[0] [1]), .ID({ID}), .\data_in_frame[0][7] (\data_in_frame[0] [7]), 
         .n65964(n65964), .pwm_setpoint({pwm_setpoint}), .\data_in_frame[0][6] (\data_in_frame[0] [6]), 
         .\data_in_frame[0][3] (\data_in_frame[0] [3]), .\data_in_frame[0][5] (\data_in_frame[0] [5]), 
         .n66998(n66998), .\data_in_frame[2][4] (\data_in_frame[2] [4]), 
         .\data_out_frame[1][5] (\data_out_frame[1] [5]), .\data_in_frame[2][6] (\data_in_frame[2] [6]), 
         .n65963(n65963), .n30143(n30143), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[1][6] (\data_in_frame[1] [6]), .\data_in_frame[2][0] (\data_in_frame[2] [0]), 
         .n51(n51), .n30139(n30139), .n22(n22_adj_5761), .\current[11] (current[11]), 
         .n30136(n30136), .n30133(n30133), .\current[15] (current[15]), 
         .n260(n260), .n65728(n65728), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n30130(n30130), .n30127(n30127), .n30124(n30124), .n30121(n30121), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .Kp_23__N_612(Kp_23__N_612), .rx_data_ready(rx_data_ready), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n66982(n66982), .\data_in_frame[18] ({\data_in_frame[18] }), .\data_in_frame[2][3] (\data_in_frame[2] [3]), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n30093(n30093), .deadband({deadband}), .n30092(n30092), .\data_in_frame[2][1] (\data_in_frame[2] [1]), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n30091(n30091), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n30090(n30090), 
         .n30089(n30089), .n30088(n30088), .n30087(n30087), .n30086(n30086), 
         .n30085(n30085), .n30084(n30084), .n30083(n30083), .n30082(n30082), 
         .n30081(n30081), .n30080(n30080), .DE_c(DE_c), .n30079(n30079), 
         .n30078(n30078), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .\data_out_frame[3][4] (\data_out_frame[3] [4]), .n30077(n30077), 
         .n30076(n30076), .n30074(n30074), .n30073(n30073), .n30072(n30072), 
         .n30071(n30071), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n71763(n71763), .n30070(n30070), .IntegralLimit({IntegralLimit}), 
         .n30069(n30069), .n30068(n30068), .n30066(n30066), .n30065(n30065), 
         .n30064(n30064), .n30063(n30063), .n30062(n30062), .n30061(n30061), 
         .n30060(n30060), .n30059(n30059), .n30058(n30058), .n30057(n30057), 
         .n30056(n30056), .n30055(n30055), .n30054(n30054), .n65962(n65962), 
         .n65961(n65961), .n65960(n65960), .n30053(n30053), .n65959(n65959), 
         .n65958(n65958), .n30052(n30052), .n65957(n65957), .n65956(n65956), 
         .n30051(n30051), .n30050(n30050), .n30049(n30049), .n30048(n30048), 
         .n30047(n30047), .\Kp[1] (Kp[1]), .n65955(n65955), .n30046(n30046), 
         .\Kp[2] (Kp[2]), .n30045(n30045), .\Kp[3] (Kp[3]), .n30044(n30044), 
         .\Kp[4] (Kp[4]), .n30043(n30043), .\Kp[5] (Kp[5]), .n30042(n30042), 
         .\Kp[6] (Kp[6]), .n65954(n65954), .n65953(n65953), .n65952(n65952), 
         .n65951(n65951), .n65950(n65950), .n30041(n30041), .\Kp[7] (Kp[7]), 
         .n30040(n30040), .\Kp[8] (Kp[8]), .n30039(n30039), .\Kp[9] (Kp[9]), 
         .n65949(n65949), .n65948(n65948), .\Kp[10] (Kp[10]), .n30037(n30037), 
         .\Kp[11] (Kp[11]), .n30036(n30036), .\Kp[12] (Kp[12]), .n65947(n65947), 
         .n65946(n65946), .n65945(n65945), .\Kp[13] (Kp[13]), .n66594(n66594), 
         .n30034(n30034), .\Kp[14] (Kp[14]), .n30033(n30033), .\Kp[15] (Kp[15]), 
         .n30032(n30032), .\Ki[1] (Ki[1]), .n30031(n30031), .\Ki[2] (Ki[2]), 
         .n30030(n30030), .\Ki[3] (Ki[3]), .n65944(n65944), .n65853(n65853), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .n65943(n65943), .n65856(n65856), 
         .n30029(n30029), .\Ki[4] (Ki[4]), .n30028(n30028), .\Ki[5] (Ki[5]), 
         .n65942(n65942), .n30027(n30027), .\Ki[6] (Ki[6]), .LED_c(LED_c), 
         .n30026(n30026), .\Ki[7] (Ki[7]), .n65861(n65861), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n65865(n65865), .n65866(n65866), .n30025(n30025), .\Ki[8] (Ki[8]), 
         .n30024(n30024), .\Ki[9] (Ki[9]), .n30023(n30023), .\Ki[10] (Ki[10]), 
         .n65867(n65867), .n30022(n30022), .\Ki[11] (Ki[11]), .n65868(n65868), 
         .n65869(n65869), .n65872(n65872), .n30021(n30021), .\Ki[12] (Ki[12]), 
         .n65875(n65875), .n29286(n29286), .n65876(n65876), .n65877(n65877), 
         .n30020(n30020), .\Ki[13] (Ki[13]), .n30019(n30019), .\Ki[14] (Ki[14]), 
         .n30018(n30018), .\Ki[15] (Ki[15]), .n65878(n65878), .n65879(n65879), 
         .n65880(n65880), .n65874(n65874), .n65881(n65881), .n65882(n65882), 
         .n65883(n65883), .n26873(n26873), .n61123(n61123), .n65884(n65884), 
         .n30005(n30005), .n30001(n30001), .neopxl_color({neopxl_color}), 
         .n74616(n74616), .n78618(n78618), .n7_adj_7(n7_adj_5796), .\data_in_frame[10] ({Open_14, 
         Open_15, Open_16, Open_17, \data_in_frame[10] [3], Open_18, 
         Open_19, Open_20}), .n30000(n30000), .n29999(n29999), .n29998(n29998), 
         .n29997(n29997), .n29996(n29996), .n29995(n29995), .n29994(n29994), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .n29993(n29993), .n29992(n29992), 
         .n29991(n29991), .n29990(n29990), .n74617(n74617), .n29989(n29989), 
         .n29988(n29988), .control_mode({Open_21, Open_22, Open_23, 
         Open_24, Open_25, Open_26, control_mode[1], Open_27}), .\control_mode[5] (control_mode[5]), 
         .\control_mode[6] (control_mode[6]), .\control_mode[7] (control_mode[7]), 
         .\current_limit[1] (current_limit[1]), .\current_limit[2] (current_limit[2]), 
         .\current_limit[3] (current_limit[3]), .\current_limit[4] (current_limit[4]), 
         .\current_limit[5] (current_limit[5]), .n29942(n29942), .PWMLimit({PWMLimit}), 
         .\current_limit[0] (current_limit[0]), .\control_mode[0] (control_mode[0]), 
         .n29939(n29939), .n29938(n29938), .\Ki[0] (Ki[0]), .n29937(n29937), 
         .\Kp[0] (Kp[0]), .n29936(n29936), .n29933(n29933), .n65885(n65885), 
         .n65886(n65886), .n65887(n65887), .n65888(n65888), .n65889(n65889), 
         .n65890(n65890), .n65891(n65891), .n65892(n65892), .n65893(n65893), 
         .n65894(n65894), .n65895(n65895), .n65896(n65896), .n65897(n65897), 
         .n65898(n65898), .n65899(n65899), .n65900(n65900), .n65901(n65901), 
         .n65902(n65902), .n65903(n65903), .n65904(n65904), .n65905(n65905), 
         .n65906(n65906), .n65907(n65907), .n65908(n65908), .n65909(n65909), 
         .n7_adj_8(n7_adj_5949), .n26329(n26329), .n8_adj_9(n8_adj_5752), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .\data_in_frame[13] ({Open_28, 
         Open_29, \data_in_frame[13] [5], Open_30, \data_in_frame[13] [3:0]}), 
         .n65910(n65910), .n29249(n29249), .n65911(n65911), .n65912(n65912), 
         .n65913(n65913), .n65914(n65914), .n7_adj_10(n7_adj_5950), .n7_adj_11(n7_adj_5951), 
         .n65873(n65873), .n66039(n66039), .n66038(n66038), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .n66037(n66037), .n66036(n66036), .\current_limit[8] (current_limit[8]), 
         .n66450(n66450), .n66166(n66166), .encoder1_position({encoder1_position[23:0]}), 
         .n69038(n69038), .\current_limit[9] (current_limit[9]), .\current_limit[10] (current_limit[10]), 
         .n65176(n65176), .n30770(n30770), .n65172(n65172), .n30766(n30766), 
         .n30764(n30764), .n30761(n30761), .n65168(n65168), .n65164(n65164), 
         .n29729(n29729), .n29732(n29732), .n30738(n30738), .n65160(n65160), 
         .n30735(n30735), .n30734(n30734), .n30732(n30732), .n30731(n30731), 
         .n30730(n30730), .n30728(n30728), .n30725(n30725), .n30723(n30723), 
         .n30721(n30721), .n30720(n30720), .n30697(n30697), .n30679(n30679), 
         .n30677(n30677), .n30676(n30676), .n30664(n30664), .n30663(n30663), 
         .n66035(n66035), .n30631(n30631), .n30630(n30630), .n30629(n30629), 
         .n30628(n30628), .n30247(n30247), .n30250(n30250), .n30624(n30624), 
         .n30253(n30253), .n30622(n30622), .n30256(n30256), .n30259(n30259), 
         .n30262(n30262), .n30617(n30617), .n30616(n30616), .n66034(n66034), 
         .n29764(n29764), .\data_in_frame[20][0] (\data_in_frame[20] [0]), 
         .n29767(n29767), .\data_in_frame[20][1] (\data_in_frame[20] [1]), 
         .n29770(n29770), .\data_in_frame[20][2] (\data_in_frame[20] [2]), 
         .n65360(n65360), .n29777(n29777), .\data_in_frame[20][3] (\data_in_frame[20] [3]), 
         .n29780(n29780), .\data_in_frame[20][4] (\data_in_frame[20] [4]), 
         .n30265(n30265), .n30601(n30601), .\data_in_frame[10][0] (\data_in_frame[10] [0]), 
         .\data_in_frame[10][5] (\data_in_frame[10] [5]), .\data_in_frame[10][6] (\data_in_frame[10] [6]), 
         .n30591(n30591), .n30587(n30587), .n30586(n30586), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
         .n30583(n30583), .n30294(n30294), .n30298(n30298), .n65336(n65336), 
         .n30304(n30304), .n30308(n30308), .n65318(n65318), .n30314(n30314), 
         .n30318(n30318), .\data_in_frame[13][6] (\data_in_frame[13] [6]), 
         .\data_in_frame[13][7] (\data_in_frame[13] [7]), .\data_in_frame[14] ({Open_31, 
         Open_32, Open_33, Open_34, Open_35, \data_in_frame[14] [2:0]}), 
         .n65863(n65863), .n65860(n65860), .\data_in_frame[14][4] (\data_in_frame[14] [4]), 
         .\data_in_frame[14][5] (\data_in_frame[14] [5]), .\data_in_frame[14][6] (\data_in_frame[14] [6]), 
         .\data_in_frame[14][7] (\data_in_frame[14] [7]), .n65154(n65154), 
         .n30430(n30430), .n65150(n65150), .n65146(n65146), .n65094(n65094), 
         .n65142(n65142), .n65244(n65244), .n30456(n30456), .n65276(n65276), 
         .n65272(n65272), .n65268(n65268), .n30515(n30515), .n66033(n66033), 
         .n29840(n29840), .\data_in_frame[23] ({\data_in_frame[23] }), .n29843(n29843), 
         .n29849(n29849), .n65134(n65134), .n29858(n29858), .n29861(n29861), 
         .n65132(n65132), .n65130(n65130), .n29870(n29870), .n29874(n29874), 
         .n29877(n29877), .n65398(n65398), .n66032(n66032), .n66031(n66031), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n65870(n65870), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n65864(n65864), 
         .n66030(n66030), .n66029(n66029), .n66028(n66028), .n71789(n71789), 
         .n71787(n71787), .n4938(n4938), .n66027(n66027), .n66026(n66026), 
         .n66025(n66025), .n66024(n66024), .n60656(n60656), .n26758(n26758), 
         .n66023(n66023), .n66022(n66022), .n66021(n66021), .n66020(n66020), 
         .n66019(n66019), .n66018(n66018), .n65974(n65974), .n66017(n66017), 
         .n66016(n66016), .n66015(n66015), .n66014(n66014), .n66013(n66013), 
         .n71786(n71786), .n71784(n71784), .n66012(n66012), .n66011(n66011), 
         .n66010(n66010), .n65915(n65915), .n65916(n65916), .\current_limit[6] (current_limit[6]), 
         .n65917(n65917), .n65918(n65918), .n65919(n65919), .n65920(n65920), 
         .n65921(n65921), .n65922(n65922), .n65923(n65923), .n65924(n65924), 
         .n65925(n65925), .n65926(n65926), .n65927(n65927), .n65928(n65928), 
         .n65929(n65929), .n66009(n66009), .n23023(n23023), .n65862(n65862), 
         .n66008(n66008), .n65859(n65859), .n65930(n65930), .n65931(n65931), 
         .n65932(n65932), .n65933(n65933), .n65934(n65934), .n65935(n65935), 
         .n65936(n65936), .n65937(n65937), .n65938(n65938), .n65939(n65939), 
         .n65857(n65857), .n65940(n65940), .n65941(n65941), .n66007(n66007), 
         .n66006(n66006), .\current_limit[7] (current_limit[7]), .n66005(n66005), 
         .n66004(n66004), .n66002(n66002), .\current[3] (current[3]), 
         .n65858(n65858), .\current[2] (current[2]), .n66001(n66001), 
         .\current[1] (current[1]), .\current[0] (current[0]), .n60808(n60808), 
         .n7_adj_12(n7_adj_5952), .n61318(n61318), .n68798(n68798), .n65754(n65754), 
         .n25794(n25794), .n8_adj_13(n8_adj_5846), .n71764(n71764), .n60646(n60646), 
         .n66463(n66463), .n34(n34_adj_5847), .n66240(n66240), .n44122(n44122), 
         .n26732(n26732), .n460(n460), .n39(n39_adj_5885), .n26478(n26478), 
         .\current[10] (current[10]), .n66388(n66388), .\current[9] (current[9]), 
         .\current[8] (current[8]), .displacement({displacement}), .n27004(n27004), 
         .n38(n38), .n486(n486), .n40(n40), .n66644(n66644), .n67902(n67902), 
         .n66992(n66992), .n67037(n67037), .tx_active(tx_active), .\pwm_counter[8] (pwm_counter[8]), 
         .n17(n17_adj_5870), .\pwm_counter[6] (pwm_counter[6]), .n13(n13_adj_5869), 
         .n66680(n66680), .n66842(n66842), .n66625(n66625), .n71771(n71771), 
         .n66244(n66244), .n71769(n71769), .n76(n76), .n78810(n78810), 
         .n78642(n78642), .n22_adj_14(n22_adj_5858), .n35278(n35278), 
         .\current[7] (current[7]), .\current[6] (current[6]), .\current[5] (current[5]), 
         .\current[4] (current[4]), .n78900(n78900), .n66788(n66788), 
         .n68353(n68353), .n66590(n66590), .n61349(n61349), .n66150(n66150), 
         .n6(n6_adj_5753), .n66769(n66769), .n27241(n27241), .n71189(n71189), 
         .n66791(n66791), .n27201(n27201), .n66751(n66751), .n66555(n66555), 
         .n70983(n70983), .n7_adj_15(n7_adj_5790), .n66660(n66660), .n68099(n68099), 
         .n45146(n45146), .n14(n14_adj_5960), .n41543(n41543), .n78834(n78834), 
         .n78498(n78498), .tx_o(tx_o), .r_SM_Main({r_SM_Main_adj_6055}), 
         .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), .n29954(n29954), 
         .r_Clock_Count({r_Clock_Count_adj_6056}), .\tx_data[3] (tx_data[3]), 
         .n67642(n67642), .n6_adj_16(n6_adj_5954), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
         .n27(n27_adj_5865), .n29(n29_adj_5864), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
         .n23(n23_adj_5866), .n5218(n5218), .n67002(n67002), .tx_enable(tx_enable), 
         .baudrate({baudrate}), .n28238(n28238), .n67079(n67079), .\r_SM_Main[2]_adj_17 (r_SM_Main[2]), 
         .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .n33(n33), .n34_adj_18(n34), 
         .n29935(n29935), .n29934(n29934), .n29932(n29932), .n29913(n29913), 
         .n29912(n29912), .n29908(n29908), .n29904(n29904), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), 
         .n5215(n5215), .\r_SM_Main[1]_adj_19 (r_SM_Main[1]), .n28115(n28115), 
         .r_Clock_Count_adj_28({r_Clock_Count}), .n30760(n30760), .n61786(n61786), 
         .n30756(n30756), .\r_Bit_Index[0] (r_Bit_Index[0]), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), 
         .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), 
         .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), 
         .n69006(n69006), .n69649(n69649), .n69585(n69585), .n69665(n69665), 
         .n69633(n69633), .n69601(n69601), .n69617(n69617), .n69697(n69697), 
         .n69681(n69681), .n69523(n69523)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i4_3_lut (.I0(encoder0_position[3]), .I1(n29), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1178_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5935));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_3812_i23_3_lut (.I0(encoder0_position[22]), .I1(n10_adj_5745), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n935));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15865_3_lut_4_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30077));   // verilog/coms.v(130[12] 305[6])
    defparam i15865_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15864_3_lut_4_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30076));   // verilog/coms.v(130[12] 305[6])
    defparam i15864_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n935), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15862_3_lut_4_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30074));   // verilog/coms.v(130[12] 305[6])
    defparam i15862_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 LessThan_1178_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5932));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5856));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15561_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n28074), .I3(GND_net), .O(n29773));   // verilog/motorControl.v(42[14] 73[8])
    defparam i15561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_1178_i8_3_lut (.I0(n6_adj_5933), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5935), .I3(GND_net), .O(n8_adj_5934));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15861_3_lut_4_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30073));   // verilog/coms.v(130[12] 305[6])
    defparam i15861_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5856), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_62717 (.I0(n11849), .I1(current[15]), .I2(duty[21]), 
            .I3(n11847), .O(n78549));
    defparam n11849_bdd_4_lut_62717.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_3812_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5749), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61448_4_lut (.I0(n8_adj_5934), .I1(n4_adj_5932), .I2(n9_adj_5935), 
            .I3(n75007), .O(n77283));   // verilog/uart_rx.v(119[17:57])
    defparam i61448_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_3812_i28_3_lut (.I0(encoder0_position[27]), .I1(n5), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n291_adj_5812));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n78549_bdd_4_lut (.I0(n78549), .I1(duty[18]), .I2(n4910), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[18]));
    defparam n78549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15860_3_lut_4_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30072));   // verilog/coms.v(130[12] 305[6])
    defparam i15860_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i61449_3_lut (.I0(n77283), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n77284));   // verilog/uart_rx.v(119[17:57])
    defparam i61449_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15859_3_lut_4_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30071));   // verilog/coms.v(130[12] 305[6])
    defparam i15859_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i61184_3_lut (.I0(n77284), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n77019));   // verilog/uart_rx.v(119[17:57])
    defparam i61184_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60060_3_lut (.I0(n77019), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5215));   // verilog/uart_rx.v(119[17:57])
    defparam i60060_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_2183 (.I0(n23_adj_5866), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5215), .I3(o_Rx_DV_N_3488[8]), .O(n69383));
    defparam i1_4_lut_adj_2183.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_2184 (.I0(o_Rx_DV_N_3488[24]), .I1(n27_adj_5865), 
            .I2(n29_adj_5864), .I3(n69383), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_2184.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_62703 (.I0(n11849), .I1(current[15]), .I2(duty[20]), 
            .I3(n11847), .O(n78531));
    defparam n11849_bdd_4_lut_62703.LUT_INIT = 16'he4aa;
    SB_LUT4 n78531_bdd_4_lut (.I0(n78531), .I1(duty[17]), .I2(n4911), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[17]));
    defparam n78531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5862), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_62690 (.I0(n11849), .I1(current[15]), .I2(duty[19]), 
            .I3(n11847), .O(n78519));
    defparam n11849_bdd_4_lut_62690.LUT_INIT = 16'he4aa;
    SB_LUT4 n78519_bdd_4_lut (.I0(n78519), .I1(duty[16]), .I2(n4912), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[16]));
    defparam n78519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_62680 (.I0(n11849), .I1(current[15]), .I2(duty[18]), 
            .I3(n11847), .O(n78513));
    defparam n11849_bdd_4_lut_62680.LUT_INIT = 16'he4aa;
    SB_LUT4 n78513_bdd_4_lut (.I0(n78513), .I1(duty[15]), .I2(n4913), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[15]));
    defparam n78513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11849_bdd_4_lut_62675 (.I0(n11849), .I1(current[15]), .I2(duty[17]), 
            .I3(n11847), .O(n78507));
    defparam n11849_bdd_4_lut_62675.LUT_INIT = 16'he4aa;
    SB_LUT4 n78507_bdd_4_lut (.I0(n78507), .I1(duty[14]), .I2(n4914), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[14]));
    defparam n78507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15858_3_lut_4_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30070));   // verilog/coms.v(130[12] 305[6])
    defparam i15858_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15857_3_lut_4_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30069));   // verilog/coms.v(130[12] 305[6])
    defparam i15857_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15856_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30068));   // verilog/coms.v(130[12] 305[6])
    defparam i15856_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2185 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n66012));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2185.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2186 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n66011));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2186.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2187 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n66010));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2187.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_2188 (.I0(state[0]), .I1(bit_ctr[3]), .I2(n44603), 
            .I3(bit_ctr[4]), .O(n4_adj_5977));   // verilog/neopixel.v(34[12] 113[6])
    defparam i1_2_lut_4_lut_adj_2188.LUT_INIT = 16'hd555;
    SB_LUT4 mux_3812_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2189 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n65915));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2189.LUT_INIT = 16'h2300;
    SB_LUT4 i15854_3_lut_4_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30066));   // verilog/coms.v(130[12] 305[6])
    defparam i15854_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3812_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5750), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3812_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam mux_3812_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15853_3_lut_4_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30065));   // verilog/coms.v(130[12] 305[6])
    defparam i15853_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i6167_2_lut (.I0(n2_adj_5751), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i6167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2190 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n65916));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2190.LUT_INIT = 16'h2300;
    SB_LUT4 i15852_3_lut_4_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30064));   // verilog/coms.v(130[12] 305[6])
    defparam i15852_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2191 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n65917));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2191.LUT_INIT = 16'h2300;
    SB_LUT4 i15851_3_lut_4_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30063));   // verilog/coms.v(130[12] 305[6])
    defparam i15851_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15850_3_lut_4_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30062));   // verilog/coms.v(130[12] 305[6])
    defparam i15850_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22720_3_lut_4_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30061));
    defparam i22720_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22676_3_lut_4_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30060));
    defparam i22676_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22677_3_lut_4_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30059));
    defparam i22677_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15846_3_lut_4_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30058));   // verilog/coms.v(130[12] 305[6])
    defparam i15846_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15845_3_lut_4_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30057));   // verilog/coms.v(130[12] 305[6])
    defparam i15845_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15844_3_lut_4_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30056));   // verilog/coms.v(130[12] 305[6])
    defparam i15844_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 n11849_bdd_4_lut_62670 (.I0(n11849), .I1(current[15]), .I2(duty[16]), 
            .I3(n11847), .O(n78489));
    defparam n11849_bdd_4_lut_62670.LUT_INIT = 16'he4aa;
    SB_LUT4 i15843_3_lut_4_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30055));   // verilog/coms.v(130[12] 305[6])
    defparam i15843_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    pwm PWM (.n2872(n2872), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .pwm_counter({Open_36, 
        Open_37, Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
        Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, Open_50, 
        pwm_counter[8], Open_51, pwm_counter[6], Open_52, Open_53, 
        Open_54, Open_55, Open_56, Open_57}), .GND_net(GND_net), .\pwm_counter[16] (pwm_counter[16]), 
        .\pwm_counter[20] (pwm_counter[20]), .\pwm_counter[19] (pwm_counter[19]), 
        .VCC_net(VCC_net), .reset(reset), .\pwm_setpoint[2] (pwm_setpoint[2]), 
        .\pwm_setpoint[3] (pwm_setpoint[3]), .\pwm_setpoint[8] (pwm_setpoint[8]), 
        .\pwm_setpoint[4] (pwm_setpoint[4]), .\pwm_setpoint[6] (pwm_setpoint[6]), 
        .\pwm_setpoint[5] (pwm_setpoint[5]), .\PWMLimit[6] (PWMLimit[6]), 
        .\data_in_frame[10][6] (\data_in_frame[10] [6]), .Kp_23__N_612(Kp_23__N_612), 
        .Kp_23__N_1748(Kp_23__N_1748), .n30764(n30764), .\pwm_setpoint[22] (pwm_setpoint[22]), 
        .\pwm_setpoint[21] (pwm_setpoint[21]), .\pwm_setpoint[12] (pwm_setpoint[12]), 
        .\pwm_setpoint[10] (pwm_setpoint[10]), .\pwm_setpoint[11] (pwm_setpoint[11]), 
        .\pwm_setpoint[9] (pwm_setpoint[9]), .\pwm_setpoint[7] (pwm_setpoint[7]), 
        .n17(n17_adj_5870), .n13(n13_adj_5869), .\pwm_setpoint[1] (pwm_setpoint[1]), 
        .\pwm_setpoint[0] (pwm_setpoint[0]), .\pwm_setpoint[13] (pwm_setpoint[13]), 
        .\pwm_setpoint[14] (pwm_setpoint[14]), .\pwm_setpoint[15] (pwm_setpoint[15]), 
        .n32(n32_adj_5871), .n34(n34_adj_5872), .\pwm_setpoint[20] (pwm_setpoint[20]), 
        .n41(n41), .n39(n39), .\pwm_setpoint[19] (pwm_setpoint[19]), .\pwm_setpoint[23] (pwm_setpoint[23]), 
        .\data_in_frame[12][7] (\data_in_frame[12] [7]), .\data_in_frame[12][0] (\data_in_frame[12] [0]), 
        .\data_in_frame[11][7] (\data_in_frame[11] [7]), .n70983(n70983), 
        .\data_in_frame[10][5] (\data_in_frame[10] [5]), .n71189(n71189), 
        .\pwm_setpoint[18] (pwm_setpoint[18]), .\pwm_setpoint[17] (pwm_setpoint[17]), 
        .n66769(n66769), .\data_in_frame[15][3] (\data_in_frame[15] [3]), 
        .n66751(n66751), .n68353(n68353), .n7(n7_adj_5790), .n69038(n69038), 
        .\data_in_frame[10][7] (\data_in_frame[10] [7]), .\data_in_frame[11][0] (\data_in_frame[11] [0]), 
        .n66791(n66791), .n26329(n26329), .n68099(n68099)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i15842_3_lut_4_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30054));   // verilog/coms.v(130[12] 305[6])
    defparam i15842_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2192 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n65918));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2192.LUT_INIT = 16'h2300;
    SB_LUT4 n78489_bdd_4_lut (.I0(n78489), .I1(duty[13]), .I2(n4915), 
            .I3(n11847), .O(pwm_setpoint_23__N_3[13]));
    defparam n78489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(322[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.enable_slow_N_4213(enable_slow_N_4213), .clk16MHz(clk16MHz), 
           .GND_net(GND_net), .data({data_adj_6032}), .baudrate({baudrate}), 
           .n28271(n28271), .data_ready(data_ready), .n29943(n29943), 
           .ID({ID}), .\state_7__N_3918[0] (state_7__N_3918[0]), .n30719(n30719), 
           .n30718(n30718), .n30717(n30717), .n30716(n30716), .n30715(n30715), 
           .n30714(n30714), .n30713(n30713), .n30704(n30704), .n30703(n30703), 
           .n30702(n30702), .n30701(n30701), .n30700(n30700), .n30699(n30699), 
           .n30698(n30698), .n30696(n30696), .n68385(n68385), .\state_7__N_4110[0] (state_7__N_4110[0]), 
           .\state[0] (state_adj_6068[0]), .scl_enable(scl_enable), .scl(scl), 
           .sda_enable(sda_enable), .sda_out(sda_out), .n11(n11_adj_5794), 
           .n29968(n29968), .n29967(n29967), .n29965(n29965), .n29964(n29964), 
           .n29963(n29963), .n29959(n29959), .n29958(n29958), .n6705(n6705), 
           .n30749(n30749), .n8(n8_adj_5974), .VCC_net(VCC_net), .n44499(n44499), 
           .\state_7__N_4126[3] (state_7__N_4126[3]), .n10(n10_adj_5953), 
           .n4(n4_adj_5792), .n4_adj_6(n4_adj_5793), .n25888(n25888), 
           .n25930(n25930), .n44644(n44644)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(391[10] 403[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2193 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n65919));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2193.LUT_INIT = 16'h2300;
    motorControl control (.PWMLimit({PWMLimit}), .GND_net(GND_net), .\Kp[6] (Kp[6]), 
            .\Kp[4] (Kp[4]), .\Ki[9] (Ki[9]), .n349(n349), .\Ki[10] (Ki[10]), 
            .IntegralLimit({IntegralLimit}), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Kp[7] (Kp[7]), .\Ki[13] (Ki[13]), 
            .\Ki[1] (Ki[1]), .n350(n350), .\Kp[8] (Kp[8]), .\Ki[0] (Ki[0]), 
            .\Kp[2] (Kp[2]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Ki[2] (Ki[2]), 
            .\Kp[3] (Kp[3]), .\Ki[3] (Ki[3]), .\Kp[11] (Kp[11]), .\Kp[5] (Kp[5]), 
            .\Ki[4] (Ki[4]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Kp[15] (Kp[15]), .n284(n284), .n258(n258), .n356(n356), 
            .n357(n357), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .n337(n337), .n313(n313), .\Ki[14] (Ki[14]), 
            .\Ki[15] (Ki[15]), .n339(n339), .n340(n340), .n358(n358), 
            .duty({duty}), .n45105(n45105), .n342(n342), .n343(n343), 
            .n344(n344), .n322(n322), .n348(n348), .n359(n359), .n336(n336), 
            .control_update(control_update), .clk16MHz(clk16MHz), .reset(reset), 
            .n345(n345), .n346(n346), .n347(n347), .VCC_net(VCC_net), 
            .setpoint({setpoint}), .motor_state({motor_state}), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .n239(n239), .n247(n247), .n467(n467), .n6(n6), .n37336(n37336), 
            .n58049(n58049), .n37146(n37146), .n475(n475), .n30514(n30514), 
            .n30513(n30513), .n30512(n30512), .n30511(n30511), .n30510(n30510), 
            .n30509(n30509), .n30508(n30508), .n30507(n30507), .n30506(n30506), 
            .n30505(n30505), .n30503(n30503), .n30501(n30501), .n30500(n30500), 
            .n30499(n30499), .n30498(n30498), .n30497(n30497), .n30496(n30496), 
            .n30495(n30495), .n30494(n30494), .n30493(n30493), .n30488(n30488), 
            .n30487(n30487), .n30479(n30479), .deadband({deadband}), .n29773(n29773), 
            .n460(n460), .n65754(n65754), .n22(n22_adj_5858), .n351(n351), 
            .n38(n38_adj_5921), .\control_mode[5] (control_mode[5]), .\control_mode[0] (control_mode[0]), 
            .\control_mode[1] (control_mode[1]), .\control_mode[6] (control_mode[6]), 
            .\control_mode[7] (control_mode[7]), .n110(n110), .n9(n9_adj_5873), 
            .n16(n16_adj_5874), .n34707(n34707), .n20(n20_adj_5875), .n25(n25_adj_5877), 
            .n33(n33_adj_5878), .n37(n37), .n41(n41_adj_5879), .n22_adj_1(n22_adj_5876), 
            .n486(n486), .n35808(n35808), .n24(n24_adj_5886), .n36173(n36173), 
            .n291(n291), .n25794(n25794), .n352(n352), .n299(n299_adj_5795), 
            .n38_adj_2(n38), .n8(n8_adj_5882), .n25_adj_3(n25_adj_5884), 
            .n10(n10_adj_5883), .n39(n39_adj_5885), .n20419(n20419), .n20420(n20420), 
            .n56(n56), .n40(n40), .n353(n353), .n354(n354), .n20466(n20466), 
            .n355(n355), .n21(n21_adj_5880), .n37_adj_4(n37_adj_5881), 
            .n57846(n57846), .n20493(n20493), .n20465(n20465)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, neopxl_color, \color_bit_N_502[1] , 
            state, GND_net, bit_ctr, n60716, n60685, n7, timer, 
            VCC_net, \bit_ctr[1] , \bit_ctr[3] , n29966, t0, n28192, 
            \bit_ctr[4] , n30582, n30581, n30580, n30579, n30578, 
            n30577, n30576, n30575, n30574, n30553, n30477, n65078, 
            NEOPXL_c, n44603, \color_bit_N_502[2] , n3163, n25404, 
            LED_c) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    input [23:0]neopxl_color;
    output \color_bit_N_502[1] ;
    output [1:0]state;
    input GND_net;
    output [4:0]bit_ctr;
    output n60716;
    output n60685;
    input n7;
    output [10:0]timer;
    input VCC_net;
    output \bit_ctr[1] ;
    output \bit_ctr[3] ;
    input n29966;
    output [10:0]t0;
    output n28192;
    output \bit_ctr[4] ;
    input n30582;
    input n30581;
    input n30580;
    input n30579;
    input n30578;
    input n30577;
    input n30576;
    input n30575;
    input n30574;
    input n30553;
    input n30477;
    input n65078;
    output NEOPXL_c;
    output n44603;
    output \color_bit_N_502[2] ;
    output n3163;
    output n25404;
    input LED_c;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n68307, \neo_pixel_transmitter.done , 
        start_N_507, n65304, start, n78783, n78786, n25906, n74675, 
        n67995, n68, n67111, n68312, n53, n44, one_wire_N_499, 
        n44538, n67008, n66063, n29446, n71854, n71853, n78582, 
        n71855, n71890, n71891, n81, n78612, n73118;
    wire [1:0]state_1__N_451;
    
    wire n25901, n25861, n6, n25904, n67117, n6_adj_5707, n66125, 
        n15, n15_adj_5708, n32, n69308;
    wire [10:0]n49;
    
    wire n59424, n59423, n59422, n59421, n59420, n59419, n59418, 
        n59417, n59416, n71904, n71905, n71902, n71901, n59415;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    wire [31:0]n149;
    
    wire n71838, n71839, n71842, n71841, n29444;
    wire [10:0]n1;
    
    wire n58427, n58426, n58425, n58424, n58423, n58422, n58421, 
        n58420, n58419, n58418, n20528, n28182, n29158, n28196, 
        n68432, n45271, n8_adj_5712, n25788, n7191, n66986, n45097, 
        n22, n25, n74666, n74664, n22988, n78609, n78579;
    
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n68307), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n65304), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 n78783_bdd_4_lut (.I0(n78783), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(\color_bit_N_502[1] ), .O(n78786));
    defparam n78783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59787_3_lut (.I0(n25906), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n74675));
    defparam i59787_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i72_4_lut (.I0(n67995), .I1(n74675), .I2(state[1]), .I3(start), 
            .O(n68));
    defparam i72_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i62644_4_lut (.I0(n67111), .I1(n68), .I2(n68312), .I3(n53), 
            .O(n44));
    defparam i62644_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30464_2_lut (.I0(n25906), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n44538));
    defparam i30464_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(start), .I1(n67008), .I2(state[1]), .I3(n66063), 
            .O(n29446));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i56019_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71854));
    defparam i56019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56018_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71853));
    defparam i56018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56020_4_lut (.I0(n71854), .I1(n78582), .I2(n60716), .I3(n60685), 
            .O(n71855));
    defparam i56020_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i56055_4_lut (.I0(n71855), .I1(n71853), .I2(n60716), .I3(\color_bit_N_502[1] ), 
            .O(n71890));
    defparam i56055_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i56056_3_lut (.I0(n71890), .I1(n78786), .I2(n7), .I3(GND_net), 
            .O(n71891));
    defparam i56056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30367_4_lut (.I0(n71891), .I1(n81), .I2(n78612), .I3(n73118), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i30367_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n25901), .I2(t1[10]), 
            .I3(t1[8]), .O(n25861));
    defparam i3_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut (.I0(n25901), .I1(t1[8]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/neopixel.v(100[14:42])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(t1[10]), .I1(n25904), .I2(t1[2]), .I3(n6), 
            .O(n25906));   // verilog/neopixel.v(100[14:42])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i22_4_lut (.I0(n66063), .I1(n67117), .I2(state[1]), .I3(start), 
            .O(n65304));
    defparam i22_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i61877_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i61877_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(t1[6]), .I1(t1[7]), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5707));   // verilog/neopixel.v(100[14:42])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1749 (.I0(t1[0]), .I1(t1[4]), .I2(GND_net), .I3(GND_net), 
            .O(n66125));
    defparam i1_2_lut_adj_1749.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1750 (.I0(t1[2]), .I1(n25904), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1750.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut (.I0(n15_adj_5708), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n53));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i3_4_lut_adj_1751 (.I0(n25901), .I1(n32), .I2(t1[10]), .I3(t1[8]), 
            .O(n69308));
    defparam i3_4_lut_adj_1751.LUT_INIT = 16'h0004;
    SB_LUT4 i2_3_lut (.I0(state[1]), .I1(n69308), .I2(start), .I3(GND_net), 
            .O(n68307));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 timer_2039_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n59424), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2039_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n59423), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_11 (.CI(n59423), .I0(GND_net), .I1(timer[9]), 
            .CO(n59424));
    SB_LUT4 timer_2039_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n59422), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_10 (.CI(n59422), .I0(GND_net), .I1(timer[8]), 
            .CO(n59423));
    SB_LUT4 timer_2039_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n59421), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_9 (.CI(n59421), .I0(GND_net), .I1(timer[7]), 
            .CO(n59422));
    SB_LUT4 timer_2039_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n59420), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_8 (.CI(n59420), .I0(GND_net), .I1(timer[6]), 
            .CO(n59421));
    SB_LUT4 timer_2039_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n59419), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_7 (.CI(n59419), .I0(GND_net), .I1(timer[5]), 
            .CO(n59420));
    SB_LUT4 timer_2039_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n59418), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_1__I_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY timer_2039_add_4_6 (.CI(n59418), .I0(GND_net), .I1(timer[4]), 
            .CO(n59419));
    SB_LUT4 timer_2039_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n59417), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_5 (.CI(n59417), .I0(GND_net), .I1(timer[3]), 
            .CO(n59418));
    SB_LUT4 timer_2039_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n59416), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_4 (.CI(n59416), .I0(GND_net), .I1(timer[2]), 
            .CO(n59417));
    SB_LUT4 i56069_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71904));
    defparam i56069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56070_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71905));
    defparam i56070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56067_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71902));
    defparam i56067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56066_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n71901));
    defparam i56066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2039_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n59415), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_3 (.CI(n59415), .I0(GND_net), .I1(timer[1]), 
            .CO(n59416));
    SB_LUT4 timer_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n59415));
    SB_LUT4 i2215_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(\bit_ctr[1] ), 
            .I2(bit_ctr[0]), .I3(\bit_ctr[3] ), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2215_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i56003_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n71838));
    defparam i56003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56004_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n71839));
    defparam i56004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56007_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n71842));
    defparam i56007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56006_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n71841));
    defparam i56006_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF timer_2039__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n29966));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n28192), 
            .D(n149[2]), .R(n29444));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(\bit_ctr[3] ), .C(clk16MHz), .E(n28192), 
            .D(n149[3]), .R(n29444));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i4 (.Q(\bit_ctr[4] ), .C(clk16MHz), .E(n28192), 
            .D(n149[4]), .R(n29444));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2039__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n30582));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n30581));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n30580));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n30579));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n30578));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n30577));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n30576));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n30575));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n30574));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n30553));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF bit_ctr_i1 (.Q(\bit_ctr[1] ), .C(clk16MHz), .D(n30477));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n65078));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n58427), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n58426), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n58426), .I0(timer[9]), .I1(n1[9]), 
            .CO(n58427));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n58425), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n58425), .I0(timer[8]), .I1(n1[8]), 
            .CO(n58426));
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n58424), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n58424), .I0(timer[7]), .I1(n1[7]), 
            .CO(n58425));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n58423), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n58423), .I0(timer[6]), .I1(n1[6]), 
            .CO(n58424));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n58422), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n58422), .I0(timer[5]), .I1(n1[5]), 
            .CO(n58423));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n58421), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n58421), .I0(timer[4]), .I1(n1[4]), 
            .CO(n58422));
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n58420), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n58420), .I0(timer[3]), .I1(n1[3]), 
            .CO(n58421));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n58419), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n58419), .I0(timer[2]), .I1(n1[2]), 
            .CO(n58420));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n1[1]), 
            .I3(n58418), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n58418), .I0(timer[1]), .I1(n1[1]), 
            .CO(n58419));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n58418));
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n28182), .D(n20528), 
            .R(n29158));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n28196), .D(state_1__N_451[0]), 
            .S(n29446));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n44), .D(one_wire_N_499), 
            .R(n68432));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i1_2_lut_adj_1752 (.I0(\bit_ctr[3] ), .I1(n44603), .I2(GND_net), 
            .I3(GND_net), .O(n60685));
    defparam i1_2_lut_adj_1752.LUT_INIT = 16'h6666;
    SB_LUT4 i1174_4_lut (.I0(\color_bit_N_502[1] ), .I1(n45271), .I2(n8_adj_5712), 
            .I3(\color_bit_N_502[2] ), .O(n81));   // verilog/neopixel.v(24[26:38])
    defparam i1174_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1753 (.I0(start), .I1(n25861), .I2(GND_net), 
            .I3(GND_net), .O(n25788));
    defparam i1_2_lut_adj_1753.LUT_INIT = 16'h4444;
    SB_LUT4 i2203_2_lut (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n7191));   // verilog/neopixel.v(65[23:32])
    defparam i2203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15233_2_lut (.I0(n28192), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29444));   // verilog/neopixel.v(34[12] 113[6])
    defparam i15233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2208_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(\bit_ctr[1] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2208_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_3_lut_4_lut (.I0(\bit_ctr[3] ), .I1(n44603), .I2(n60716), 
            .I3(bit_ctr[0]), .O(n8_adj_5712));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hff9f;
    SB_LUT4 i51201_2_lut (.I0(t1[10]), .I1(t1[9]), .I2(GND_net), .I3(GND_net), 
            .O(n66986));
    defparam i51201_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51325_4_lut (.I0(t1[8]), .I1(n66986), .I2(n6_adj_5707), .I3(t1[5]), 
            .O(n67111));
    defparam i51325_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31023_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n45097));
    defparam i31023_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i58874_4_lut (.I0(n22), .I1(n25), .I2(n45097), .I3(state[0]), 
            .O(n74666));
    defparam i58874_4_lut.LUT_INIT = 16'h0c0a;
    SB_LUT4 i60091_4_lut (.I0(n74666), .I1(t1[4]), .I2(t1[2]), .I3(n67111), 
            .O(n74664));
    defparam i60091_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i45_3_lut (.I0(n74664), .I1(state[1]), .I2(start), .I3(GND_net), 
            .O(n3163));
    defparam i45_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_4_lut (.I0(n15_adj_5708), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(n15), .O(n32));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h14d7;
    SB_LUT4 i3_3_lut_4_lut_adj_1754 (.I0(t1[9]), .I1(t1[6]), .I2(t1[7]), 
            .I3(t1[5]), .O(n25901));   // verilog/neopixel.v(100[14:42])
    defparam i3_3_lut_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(t1[1]), .I1(t1[0]), .I2(t1[4]), .I3(t1[3]), 
            .O(n25904));   // verilog/neopixel.v(60[15:45])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46_3_lut_4_lut_3_lut (.I0(t1[3]), .I1(t1[1]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n25));
    defparam i46_3_lut_4_lut_3_lut.LUT_INIT = 16'h1818;
    SB_LUT4 i47_3_lut_4_lut_3_lut (.I0(t1[3]), .I1(t1[1]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n22));
    defparam i47_3_lut_4_lut_3_lut.LUT_INIT = 16'h8181;
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6672_3_lut_4_lut (.I0(bit_ctr[0]), .I1(start), .I2(n25861), 
            .I3(n22988), .O(n20528));   // verilog/neopixel.v(35[4] 112[11])
    defparam i6672_3_lut_4_lut.LUT_INIT = 16'haa9a;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_1__I_0_103_Mux_0_i1_3_lut_4_lut (.I0(n15_adj_5708), .I1(t1[2]), 
            .I2(n25904), .I3(state[0]), .O(n22988));   // verilog/neopixel.v(35[4] 112[11])
    defparam state_1__I_0_103_Mux_0_i1_3_lut_4_lut.LUT_INIT = 16'hf3aa;
    SB_LUT4 i57283_2_lut_3_lut (.I0(n60716), .I1(\bit_ctr[3] ), .I2(n44603), 
            .I3(GND_net), .O(n73118));   // verilog/neopixel.v(24[26:38])
    defparam i57283_2_lut_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51223_2_lut_3_lut (.I0(n25906), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n67008));
    defparam i51223_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1755 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(t1[2]), .I3(n25904), .O(n68312));
    defparam i2_3_lut_4_lut_adj_1755.LUT_INIT = 16'h0080;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(\bit_ctr[1] ), .O(n78783));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_4_lut_4_lut_adj_1756 (.I0(n25404), .I1(state[1]), .I2(n44538), 
            .I3(state[0]), .O(n28196));
    defparam i1_4_lut_4_lut_adj_1756.LUT_INIT = 16'hee2e;
    SB_LUT4 i1_2_lut_3_lut (.I0(n25404), .I1(state[1]), .I2(n28182), .I3(GND_net), 
            .O(n28192));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n28182));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h20ff;
    SB_LUT4 i14946_2_lut_4_lut (.I0(state[0]), .I1(n81), .I2(LED_c), .I3(state[1]), 
            .O(n29158));   // verilog/neopixel.v(35[4] 112[11])
    defparam i14946_2_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_adj_1757 (.I0(\bit_ctr[3] ), .I1(n44603), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n60716));
    defparam i1_2_lut_3_lut_adj_1757.LUT_INIT = 16'h7878;
    SB_LUT4 i31191_2_lut_3_lut (.I0(\bit_ctr[3] ), .I1(n44603), .I2(\bit_ctr[4] ), 
            .I3(GND_net), .O(n45271));
    defparam i31191_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i30529_2_lut_3_lut (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n44603));
    defparam i30529_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1758 (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), 
            .I2(bit_ctr_c[2]), .I3(GND_net), .O(\color_bit_N_502[2] ));
    defparam i1_2_lut_3_lut_adj_1758.LUT_INIT = 16'h1e1e;
    SB_LUT4 i2222_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n7191), .I2(\bit_ctr[3] ), 
            .I3(\bit_ctr[4] ), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2222_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(\color_bit_N_502[1] ), .I1(n71841), 
            .I2(n71842), .I3(\color_bit_N_502[2] ), .O(n78609));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n78609_bdd_4_lut (.I0(n78609), .I1(n71839), .I2(n71838), .I3(\color_bit_N_502[2] ), 
            .O(n78612));
    defparam n78609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2201_2_lut (.I0(\bit_ctr[1] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(\color_bit_N_502[1] ));   // verilog/neopixel.v(65[23:32])
    defparam i2201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_62751 (.I0(\color_bit_N_502[1] ), 
            .I1(n71901), .I2(n71902), .I3(\color_bit_N_502[2] ), .O(n78579));
    defparam color_bit_N_502_1__bdd_4_lut_62751.LUT_INIT = 16'he4aa;
    SB_LUT4 n78579_bdd_4_lut (.I0(n78579), .I1(n71905), .I2(n71904), .I3(\color_bit_N_502[2] ), 
            .O(n78582));
    defparam n78579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_4_lut_adj_1759 (.I0(t1[1]), .I1(t1[3]), .I2(t1[2]), 
            .I3(n66125), .O(n15_adj_5708));
    defparam i3_3_lut_4_lut_adj_1759.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_1760 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25906), .I3(state[1]), .O(n68432));
    defparam i2_3_lut_4_lut_adj_1760.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_1761 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n67111), .I3(n15), .O(n67995));
    defparam i2_3_lut_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_LUT4 i51331_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25906), .I3(GND_net), .O(n67117));
    defparam i51331_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1762 (.I0(n15_adj_5708), .I1(n15), .I2(state[0]), 
            .I3(n25788), .O(n25404));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut_adj_1762.LUT_INIT = 16'h3500;
    SB_LUT4 i1_2_lut_4_lut_adj_1763 (.I0(n15_adj_5708), .I1(n15), .I2(state[0]), 
            .I3(n25861), .O(n66063));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut_adj_1763.LUT_INIT = 16'h3500;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1779, ENCODER0_A_N_keep, 
            n30010, n1742, n30006, a_prev, n29984, b_prev, position_31__N_3836, 
            n1744, \encoder0_position[30] , \encoder0_position[29] , \encoder0_position[28] , 
            \encoder0_position[27] , \encoder0_position[26] , \encoder0_position[25] , 
            \encoder0_position[24] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , \a_new[1] , \b_new[1] , GND_net, 
            VCC_net, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    input n30010;
    output n1742;
    input n30006;
    output a_prev;
    input n29984;
    output b_prev;
    output position_31__N_3836;
    output n1744;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    output \a_new[1] ;
    output \b_new[1] ;
    input GND_net;
    input VCC_net;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n59580, n59579, n59578, n59577, n59576, 
        n59575, n59574, n59573, n59572, n59571, n59570, n59569, 
        n59568, n59567, n59566, n59565, n59564, n59563, n59562, 
        n59561, n59560, n59559, n59558, n59557, n59556, n59555, 
        n59554, n59553, n59552, n59551, n59550;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1742), .C(n1779), .D(n30010));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n30006));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29984));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1744), .I3(n59580), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[30] ), .I3(n59579), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n59579), .I0(direction_N_3840), 
            .I1(\encoder0_position[30] ), .CO(n59580));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[29] ), .I3(n59578), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n59578), .I0(direction_N_3840), 
            .I1(\encoder0_position[29] ), .CO(n59579));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[28] ), .I3(n59577), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n59577), .I0(direction_N_3840), 
            .I1(\encoder0_position[28] ), .CO(n59578));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[27] ), .I3(n59576), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n59576), .I0(direction_N_3840), 
            .I1(\encoder0_position[27] ), .CO(n59577));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[26] ), .I3(n59575), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n59575), .I0(direction_N_3840), 
            .I1(\encoder0_position[26] ), .CO(n59576));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[25] ), .I3(n59574), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n59574), .I0(direction_N_3840), 
            .I1(\encoder0_position[25] ), .CO(n59575));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[24] ), .I3(n59573), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n59573), .I0(direction_N_3840), 
            .I1(\encoder0_position[24] ), .CO(n59574));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[23] ), .I3(n59572), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n59572), .I0(direction_N_3840), 
            .I1(\encoder0_position[23] ), .CO(n59573));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n59571), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n59571), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n59572));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n59570), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n59570), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n59571));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n59569), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n59569), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n59570));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n59568), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n59568), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n59569));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n59567), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n59567), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n59568));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n59566), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n59566), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n59567));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n59565), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n59565), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n59566));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n59564), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n59564), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n59565));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n59563), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n59563), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n59564));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n59562), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n59562), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n59563));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n59561), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n59561), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n59562));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n59560), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n59560), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n59561));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n59559), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n59559), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n59560));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n59558), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n59558), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n59559));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n59557), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n59557), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n59558));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n59556), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n59556), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n59557));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n59555), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n59555), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n59556));
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n59554), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n59554), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n59555));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n59553), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_6 (.CI(n59553), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n59554));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n59552), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n59552), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n59553));
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n59551), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n59551), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n59552));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n59550), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n59550), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n59551));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n59550));
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (VCC_net, GND_net, clk16MHz, n5, n5_adj_29, n5_adj_30, 
            \state[0] , \state[1] , state_7__N_4319, n44573, clk_out, 
            CS_c, CS_CLK_c, n15, n30117, \data[15] , n30116, \data[12] , 
            n30115, \data[11] , n30114, \data[10] , n30113, \data[9] , 
            n30112, \data[8] , n30111, \data[7] , n30110, \data[6] , 
            n30109, \data[5] , n30108, \data[4] , n30107, \data[3] , 
            n30106, \data[2] , n30105, \data[1] , n25893, n11, n25910, 
            n25867, n9, n29947, n29945, \current[0] , n30765, \data[0] , 
            n30675, \current[1] , n30674, \current[2] , n30673, \current[3] , 
            n30672, \current[4] , n30671, \current[5] , n30670, \current[6] , 
            n30669, \current[7] , n30668, \current[8] , n30667, \current[9] , 
            n30666, \current[10] , n30665, \current[11] , n28097, 
            \current[15] , n25883) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    input clk16MHz;
    output n5;
    output n5_adj_29;
    output n5_adj_30;
    output \state[0] ;
    output \state[1] ;
    output state_7__N_4319;
    output n44573;
    output clk_out;
    output CS_c;
    output CS_CLK_c;
    output n15;
    input n30117;
    output \data[15] ;
    input n30116;
    output \data[12] ;
    input n30115;
    output \data[11] ;
    input n30114;
    output \data[10] ;
    input n30113;
    output \data[9] ;
    input n30112;
    output \data[8] ;
    input n30111;
    output \data[7] ;
    input n30110;
    output \data[6] ;
    input n30109;
    output \data[5] ;
    input n30108;
    output \data[4] ;
    input n30107;
    output \data[3] ;
    input n30106;
    output \data[2] ;
    input n30105;
    output \data[1] ;
    output n25893;
    output n11;
    output n25910;
    output n25867;
    input n9;
    input n29947;
    input n29945;
    output \current[0] ;
    input n30765;
    output \data[0] ;
    input n30675;
    output \current[1] ;
    input n30674;
    output \current[2] ;
    input n30673;
    output \current[3] ;
    input n30672;
    output \current[4] ;
    input n30671;
    output \current[5] ;
    input n30670;
    output \current[6] ;
    input n30669;
    output \current[7] ;
    input n30668;
    output \current[8] ;
    input n30667;
    output \current[9] ;
    input n30666;
    output \current[10] ;
    input n30665;
    output \current[11] ;
    output n28097;
    output \current[15] ;
    output n25883;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n59510, clk_slow_N_4232, n45148, n2, n12493, n28261, n29165, 
        n22860, n28154;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4314;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4233, n22862, n22864, n22866;
    wire [7:0]n37;
    
    wire n29433;
    wire [13:0]n241;
    
    wire n74521, n74522, n74526, n74527, n59542, n59541, n59540, 
        n59539, n59538, n59537, n59536, n59535, n59534, n59533, 
        n59532, n59531, n59530, n59516, n59515, n59514, n59513, 
        n59512, n59511, n4, n8, n12, n10;
    
    SB_CARRY bit_counter_2044_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n59510));
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_29));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_330_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_30));   // verilog/tli4970.v(54[9:26])
    defparam equal_330_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i30499_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n44573));
    defparam i30499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i61938_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n45148));
    defparam i61938_2_lut.LUT_INIT = 16'h1111;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n30117));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n30116));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n30115));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n30114));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n30113));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n30112));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n30111));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n30110));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n30109));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n30108));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n30107));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n30106));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n30105));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n25893));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1747 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n25910));
    defparam i1_2_lut_3_lut_4_lut_adj_1747.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1748 (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n25867));
    defparam i1_2_lut_3_lut_4_lut_adj_1748.LUT_INIT = 16'hffbf;
    SB_LUT4 i2521_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));
    defparam i2521_1_lut.LUT_INIT = 16'h5555;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n28261), .D(n12493), 
            .R(n29165));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29947));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29945));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n28154), 
            .D(n22860));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2048_2049__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNE bit_counter_2044__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n28154), 
            .D(n22862));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n28154), 
            .D(n22864));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n28154), 
            .D(n22866));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n28154), 
            .D(n37[4]), .R(n29433));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n28154), 
            .D(n37[5]), .R(n29433));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n28154), 
            .D(n37[6]), .R(n29433));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n28154), 
            .D(n37[7]), .R(n29433));   // verilog/tli4970.v(55[24:39])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30765));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30675));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30674));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30673));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30672));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30671));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30670));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30669));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30668));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30667));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30666));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30665));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n28097), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n28261), .D(n45148), 
            .S(n29165));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i8936_3_lut (.I0(\state[0] ), .I1(n74521), .I2(\state[1] ), 
            .I3(GND_net), .O(n22866));   // verilog/tli4970.v(55[24:39])
    defparam i8936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8934_3_lut (.I0(\state[0] ), .I1(n74522), .I2(\state[1] ), 
            .I3(GND_net), .O(n22864));   // verilog/tli4970.v(55[24:39])
    defparam i8934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8932_3_lut (.I0(\state[0] ), .I1(n74526), .I2(\state[1] ), 
            .I3(GND_net), .O(n22862));   // verilog/tli4970.v(55[24:39])
    defparam i8932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14096_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28154));
    defparam i14096_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8930_3_lut (.I0(\state[0] ), .I1(n74527), .I2(\state[1] ), 
            .I3(GND_net), .O(n22860));   // verilog/tli4970.v(55[24:39])
    defparam i8930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2050_2051_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n59542), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2050_2051_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n59541), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_3 (.CI(n59541), .I0(GND_net), .I1(counter[1]), 
            .CO(n59542));
    SB_LUT4 counter_2050_2051_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n59541));
    SB_LUT4 delay_counter_2048_2049_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n59540), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2048_2049_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n59539), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_12 (.CI(n59539), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n59540));
    SB_LUT4 delay_counter_2048_2049_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n59538), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_11 (.CI(n59538), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n59539));
    SB_LUT4 delay_counter_2048_2049_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n59537), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_10 (.CI(n59537), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n59538));
    SB_LUT4 delay_counter_2048_2049_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n59536), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_9 (.CI(n59536), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n59537));
    SB_LUT4 delay_counter_2048_2049_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n59535), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_8 (.CI(n59535), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n59536));
    SB_LUT4 delay_counter_2048_2049_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n59534), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_7 (.CI(n59534), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n59535));
    SB_LUT4 delay_counter_2048_2049_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n59533), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_6 (.CI(n59533), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n59534));
    SB_LUT4 delay_counter_2048_2049_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n59532), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_5 (.CI(n59532), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n59533));
    SB_LUT4 delay_counter_2048_2049_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n59531), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_4 (.CI(n59531), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n59532));
    SB_LUT4 delay_counter_2048_2049_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n59530), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_3 (.CI(n59530), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n59531));
    SB_LUT4 delay_counter_2048_2049_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n59530));
    SB_LUT4 bit_counter_2044_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n59516), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2044_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n59515), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_8 (.CI(n59515), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n59516));
    SB_LUT4 bit_counter_2044_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n59514), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_7 (.CI(n59514), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n59515));
    SB_LUT4 bit_counter_2044_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n59513), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_6 (.CI(n59513), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n59514));
    SB_LUT4 bit_counter_2044_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n59512), .O(n74526)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_5 (.CI(n59512), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n59513));
    SB_LUT4 bit_counter_2044_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n59511), .O(n74522)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_4 (.CI(n59511), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n59512));
    SB_LUT4 bit_counter_2044_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n59510), .O(n74521)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_3 (.CI(n59510), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n59511));
    SB_LUT4 bit_counter_2044_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n74527)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15222_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29433));   // verilog/tli4970.v(55[24:39])
    defparam i15222_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i61898_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n28097));
    defparam i61898_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut (.I0(bit_counter[4]), .I1(bit_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(n11), .I1(bit_counter[5]), .I2(bit_counter[7]), 
            .I3(n4), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2180_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2180_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 mux_2153_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n12493));
    defparam mux_2153_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2243_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2243_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n28261));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i14953_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n29165));
    defparam i14953_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n25883));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2179_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2179_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, 
            n1786, GND_net, n1788, n1790, n1792, n1794, n1796, 
            \encoder1_position[25] , \encoder1_position[24] , \encoder1_position[23] , 
            \encoder1_position[22] , \encoder1_position[21] , \encoder1_position[20] , 
            \encoder1_position[19] , \encoder1_position[18] , \encoder1_position[17] , 
            \encoder1_position[16] , \encoder1_position[15] , \encoder1_position[14] , 
            \encoder1_position[13] , \encoder1_position[12] , \encoder1_position[11] , 
            \encoder1_position[10] , \encoder1_position[9] , \encoder1_position[8] , 
            \encoder1_position[7] , \encoder1_position[6] , \encoder1_position[5] , 
            \encoder1_position[4] , \encoder1_position[3] , \encoder1_position[2] , 
            \encoder1_position[1] , \encoder1_position[0] , VCC_net, n30011, 
            a_prev, n29957, b_prev, n29956, n1784, position_31__N_3836, 
            \a_new[1] , \b_new[1] , debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    output n1786;
    input GND_net;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output \encoder1_position[1] ;
    output \encoder1_position[0] ;
    input VCC_net;
    input n30011;
    output a_prev;
    input n29957;
    output b_prev;
    input n29956;
    output n1784;
    output position_31__N_3836;
    output \a_new[1] ;
    output \b_new[1] ;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n59478, n59477, n59476, n59475, n59474, 
        n59473, n59472, n59471, n59470, n59469, n59468, n59467, 
        n59466, n59465, n59464, n59463, n59462, n59461, n59460, 
        n59459, n59458, n59457, n59456, n59455, n59454, n59453, 
        n59452, n59451, n59450, n59449, n59448;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2041_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1786), .I3(n59478), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2041_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1788), .I3(n59477), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_32 (.CI(n59477), .I0(direction_N_3840), 
            .I1(n1788), .CO(n59478));
    SB_LUT4 position_2041_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1790), .I3(n59476), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_31 (.CI(n59476), .I0(direction_N_3840), 
            .I1(n1790), .CO(n59477));
    SB_LUT4 position_2041_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1792), .I3(n59475), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_30 (.CI(n59475), .I0(direction_N_3840), 
            .I1(n1792), .CO(n59476));
    SB_LUT4 position_2041_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1794), .I3(n59474), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_29 (.CI(n59474), .I0(direction_N_3840), 
            .I1(n1794), .CO(n59475));
    SB_LUT4 position_2041_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1796), .I3(n59473), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_28 (.CI(n59473), .I0(direction_N_3840), 
            .I1(n1796), .CO(n59474));
    SB_LUT4 position_2041_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[25] ), .I3(n59472), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_27 (.CI(n59472), .I0(direction_N_3840), 
            .I1(\encoder1_position[25] ), .CO(n59473));
    SB_LUT4 position_2041_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[24] ), .I3(n59471), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_26 (.CI(n59471), .I0(direction_N_3840), 
            .I1(\encoder1_position[24] ), .CO(n59472));
    SB_LUT4 position_2041_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[23] ), .I3(n59470), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_25 (.CI(n59470), .I0(direction_N_3840), 
            .I1(\encoder1_position[23] ), .CO(n59471));
    SB_LUT4 position_2041_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[22] ), .I3(n59469), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_24 (.CI(n59469), .I0(direction_N_3840), 
            .I1(\encoder1_position[22] ), .CO(n59470));
    SB_LUT4 position_2041_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[21] ), .I3(n59468), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_23 (.CI(n59468), .I0(direction_N_3840), 
            .I1(\encoder1_position[21] ), .CO(n59469));
    SB_LUT4 position_2041_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[20] ), .I3(n59467), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_22 (.CI(n59467), .I0(direction_N_3840), 
            .I1(\encoder1_position[20] ), .CO(n59468));
    SB_LUT4 position_2041_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[19] ), .I3(n59466), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_21 (.CI(n59466), .I0(direction_N_3840), 
            .I1(\encoder1_position[19] ), .CO(n59467));
    SB_LUT4 position_2041_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[18] ), .I3(n59465), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_20 (.CI(n59465), .I0(direction_N_3840), 
            .I1(\encoder1_position[18] ), .CO(n59466));
    SB_LUT4 position_2041_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[17] ), .I3(n59464), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_19 (.CI(n59464), .I0(direction_N_3840), 
            .I1(\encoder1_position[17] ), .CO(n59465));
    SB_LUT4 position_2041_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[16] ), .I3(n59463), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_18 (.CI(n59463), .I0(direction_N_3840), 
            .I1(\encoder1_position[16] ), .CO(n59464));
    SB_LUT4 position_2041_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[15] ), .I3(n59462), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_17 (.CI(n59462), .I0(direction_N_3840), 
            .I1(\encoder1_position[15] ), .CO(n59463));
    SB_LUT4 position_2041_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[14] ), .I3(n59461), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_16 (.CI(n59461), .I0(direction_N_3840), 
            .I1(\encoder1_position[14] ), .CO(n59462));
    SB_LUT4 position_2041_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[13] ), .I3(n59460), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_15 (.CI(n59460), .I0(direction_N_3840), 
            .I1(\encoder1_position[13] ), .CO(n59461));
    SB_LUT4 position_2041_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[12] ), .I3(n59459), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_14 (.CI(n59459), .I0(direction_N_3840), 
            .I1(\encoder1_position[12] ), .CO(n59460));
    SB_LUT4 position_2041_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[11] ), .I3(n59458), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_13 (.CI(n59458), .I0(direction_N_3840), 
            .I1(\encoder1_position[11] ), .CO(n59459));
    SB_LUT4 position_2041_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[10] ), .I3(n59457), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_12 (.CI(n59457), .I0(direction_N_3840), 
            .I1(\encoder1_position[10] ), .CO(n59458));
    SB_LUT4 position_2041_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[9] ), .I3(n59456), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_11 (.CI(n59456), .I0(direction_N_3840), 
            .I1(\encoder1_position[9] ), .CO(n59457));
    SB_LUT4 position_2041_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[8] ), .I3(n59455), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_10 (.CI(n59455), .I0(direction_N_3840), 
            .I1(\encoder1_position[8] ), .CO(n59456));
    SB_LUT4 position_2041_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[7] ), .I3(n59454), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_9 (.CI(n59454), .I0(direction_N_3840), 
            .I1(\encoder1_position[7] ), .CO(n59455));
    SB_LUT4 position_2041_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[6] ), .I3(n59453), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_8 (.CI(n59453), .I0(direction_N_3840), 
            .I1(\encoder1_position[6] ), .CO(n59454));
    SB_LUT4 position_2041_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[5] ), .I3(n59452), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_7 (.CI(n59452), .I0(direction_N_3840), 
            .I1(\encoder1_position[5] ), .CO(n59453));
    SB_LUT4 position_2041_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[4] ), .I3(n59451), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_6 (.CI(n59451), .I0(direction_N_3840), 
            .I1(\encoder1_position[4] ), .CO(n59452));
    SB_LUT4 position_2041_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[3] ), .I3(n59450), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_5 (.CI(n59450), .I0(direction_N_3840), 
            .I1(\encoder1_position[3] ), .CO(n59451));
    SB_LUT4 position_2041_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[2] ), .I3(n59449), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_4 (.CI(n59449), .I0(direction_N_3840), 
            .I1(\encoder1_position[2] ), .CO(n59450));
    SB_LUT4 position_2041_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[1] ), .I3(n59448), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_3 (.CI(n59448), .I0(direction_N_3840), 
            .I1(\encoder1_position[1] ), .CO(n59449));
    SB_LUT4 position_2041_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder1_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder1_position[0] ), 
            .CO(n59448));
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1779), .D(n30011));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1779), .D(n29957));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1784), .C(n1779), .D(n29956));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i0 (.Q(\encoder1_position[0] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i1 (.Q(\encoder1_position[1] ), .C(n1779), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1779), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[13] , \FRAME_MATCHER.i_31__N_2509 , setpoint, 
            VCC_net, \data_in_frame[8] , clk16MHz, \data_out_frame[3][3] , 
            GND_net, n2872, \data_out_frame[8] , n66000, n65999, byte_transmit_counter, 
            \data_out_frame[25] , \data_out_frame[24] , n78804, \data_out_frame[1][1] , 
            \data_out_frame[3][1] , \data_out_frame[6] , \data_out_frame[7] , 
            n71810, \data_out_frame[4] , \data_out_frame[5] , n71808, 
            rx_data, n7, \data_in_frame[2] , \data_in_frame[3] , \data_in_frame[6] , 
            \data_in_frame[16] , n28715, n65854, \data_out_frame[14] , 
            \data_out_frame[15] , \data_out_frame[12] , Kp_23__N_1748, 
            reset, n8, n65998, \data_out_frame[1][7] , \data_out_frame[1][6] , 
            \data_in_frame[5] , n65997, n66003, n65996, \data_out_frame[9] , 
            n66040, n65995, n65994, n65993, n65992, n65991, n65990, 
            n65989, \data_out_frame[10] , n65855, n65988, n65987, 
            n65986, n65985, n65984, \FRAME_MATCHER.i[5] , \FRAME_MATCHER.i[4] , 
            \FRAME_MATCHER.i[3] , n65983, n65982, \data_out_frame[11] , 
            n65981, n65980, n65979, n65978, n65977, n65976, n65975, 
            n65871, n65973, n65972, n65971, n65970, n65969, n65968, 
            \data_in_frame[1][0] , encoder0_position, n65967, \data_out_frame[0][2] , 
            n65966, \data_out_frame[18] , \data_out_frame[19] , n71801, 
            \data_out_frame[17] , \data_out_frame[16] , n71799, n78768, 
            n65965, \data_in_frame[0][0] , \data_in_frame[0][1] , ID, 
            \data_in_frame[0][7] , n65964, pwm_setpoint, \data_in_frame[0][6] , 
            \data_in_frame[0][3] , \data_in_frame[0][5] , n66998, \data_in_frame[2][4] , 
            \data_out_frame[1][5] , \data_in_frame[2][6] , n65963, n30143, 
            \data_in_frame[4] , \data_in_frame[1][6] , \data_in_frame[2][0] , 
            n51, n30139, n22, \current[11] , n30136, n30133, \current[15] , 
            n260, n65728, \data_out_frame[1][3] , n30130, n30127, 
            n30124, n30121, \FRAME_MATCHER.state[3] , \data_in_frame[17] , 
            Kp_23__N_612, rx_data_ready, \FRAME_MATCHER.rx_data_ready_prev , 
            n66982, \data_in_frame[18] , \data_in_frame[2][3] , \data_out_frame[23] , 
            \data_out_frame[21] , n30093, deadband, n30092, \data_in_frame[2][1] , 
            \data_out_frame[20] , n30091, \data_out_frame[22] , n30090, 
            n30089, n30088, n30087, n30086, n30085, n30084, n30083, 
            n30082, n30081, n30080, DE_c, n30079, n30078, \data_out_frame[0][4] , 
            \data_out_frame[3][4] , n30077, n30076, n30074, n30073, 
            n30072, n30071, \data_out_frame[0][3] , n71763, n30070, 
            IntegralLimit, n30069, n30068, n30066, n30065, n30064, 
            n30063, n30062, n30061, n30060, n30059, n30058, n30057, 
            n30056, n30055, n30054, n65962, n65961, n65960, n30053, 
            n65959, n65958, n30052, n65957, n65956, n30051, n30050, 
            n30049, n30048, n30047, \Kp[1] , n65955, n30046, \Kp[2] , 
            n30045, \Kp[3] , n30044, \Kp[4] , n30043, \Kp[5] , n30042, 
            \Kp[6] , n65954, n65953, n65952, n65951, n65950, n30041, 
            \Kp[7] , n30040, \Kp[8] , n30039, \Kp[9] , n65949, n65948, 
            \Kp[10] , n30037, \Kp[11] , n30036, \Kp[12] , n65947, 
            n65946, n65945, \Kp[13] , n66594, n30034, \Kp[14] , 
            n30033, \Kp[15] , n30032, \Ki[1] , n30031, \Ki[2] , 
            n30030, \Ki[3] , n65944, n65853, \data_in_frame[12] , 
            n65943, n65856, n30029, \Ki[4] , n30028, \Ki[5] , n65942, 
            n30027, \Ki[6] , LED_c, n30026, \Ki[7] , n65861, \data_in_frame[9] , 
            n65865, n65866, n30025, \Ki[8] , n30024, \Ki[9] , n30023, 
            \Ki[10] , n65867, n30022, \Ki[11] , n65868, n65869, 
            n65872, n30021, \Ki[12] , n65875, n29286, n65876, n65877, 
            n30020, \Ki[13] , n30019, \Ki[14] , n30018, \Ki[15] , 
            n65878, n65879, n65880, n65874, n65881, n65882, n65883, 
            n26873, n61123, n65884, n30005, n30001, neopxl_color, 
            n74616, n78618, n7_adj_7, \data_in_frame[10] , n30000, 
            n29999, n29998, n29997, n29996, n29995, n29994, \data_in_frame[11] , 
            n29993, n29992, n29991, n29990, n74617, n29989, n29988, 
            control_mode, \control_mode[5] , \control_mode[6] , \control_mode[7] , 
            \current_limit[1] , \current_limit[2] , \current_limit[3] , 
            \current_limit[4] , \current_limit[5] , n29942, PWMLimit, 
            \current_limit[0] , \control_mode[0] , n29939, n29938, \Ki[0] , 
            n29937, \Kp[0] , n29936, n29933, n65885, n65886, n65887, 
            n65888, n65889, n65890, n65891, n65892, n65893, n65894, 
            n65895, n65896, n65897, n65898, n65899, n65900, n65901, 
            n65902, n65903, n65904, n65905, n65906, n65907, n65908, 
            n65909, n7_adj_8, n26329, n8_adj_9, \data_in_frame[15] , 
            \data_in_frame[13] , n65910, n29249, n65911, n65912, n65913, 
            n65914, n7_adj_10, n7_adj_11, n65873, n66039, n66038, 
            \data_out_frame[1][0] , n66037, n66036, \current_limit[8] , 
            n66450, n66166, encoder1_position, n69038, \current_limit[9] , 
            \current_limit[10] , n65176, n30770, n65172, n30766, n30764, 
            n30761, n65168, n65164, n29729, n29732, n30738, n65160, 
            n30735, n30734, n30732, n30731, n30730, n30728, n30725, 
            n30723, n30721, n30720, n30697, n30679, n30677, n30676, 
            n30664, n30663, n66035, n30631, n30630, n30629, n30628, 
            n30247, n30250, n30624, n30253, n30622, n30256, n30259, 
            n30262, n30617, n30616, n66034, n29764, \data_in_frame[20][0] , 
            n29767, \data_in_frame[20][1] , n29770, \data_in_frame[20][2] , 
            n65360, n29777, \data_in_frame[20][3] , n29780, \data_in_frame[20][4] , 
            n30265, n30601, \data_in_frame[10][0] , \data_in_frame[10][5] , 
            \data_in_frame[10][6] , n30591, n30587, n30586, \data_in_frame[10][7] , 
            n30583, n30294, n30298, n65336, n30304, n30308, n65318, 
            n30314, n30318, \data_in_frame[13][6] , \data_in_frame[13][7] , 
            \data_in_frame[14] , n65863, n65860, \data_in_frame[14][4] , 
            \data_in_frame[14][5] , \data_in_frame[14][6] , \data_in_frame[14][7] , 
            n65154, n30430, n65150, n65146, n65094, n65142, n65244, 
            n30456, n65276, n65272, n65268, n30515, n66033, n29840, 
            \data_in_frame[23] , n29843, n29849, n65134, n29858, n29861, 
            n65132, n65130, n29870, n29874, n29877, n65398, n66032, 
            n66031, \data_out_frame[3][6] , n65870, \data_out_frame[3][7] , 
            n65864, n66030, n66029, n66028, n71789, n71787, n4938, 
            n66027, n66026, n66025, n66024, n60656, n26758, n66023, 
            n66022, n66021, n66020, n66019, n66018, n65974, n66017, 
            n66016, n66015, n66014, n66013, n71786, n71784, n66012, 
            n66011, n66010, n65915, n65916, \current_limit[6] , n65917, 
            n65918, n65919, n65920, n65921, n65922, n65923, n65924, 
            n65925, n65926, n65927, n65928, n65929, n66009, n23023, 
            n65862, n66008, n65859, n65930, n65931, n65932, n65933, 
            n65934, n65935, n65936, n65937, n65938, n65939, n65857, 
            n65940, n65941, n66007, n66006, \current_limit[7] , n66005, 
            n66004, n66002, \current[3] , n65858, \current[2] , n66001, 
            \current[1] , \current[0] , n60808, n7_adj_12, n61318, 
            n68798, n65754, n25794, n8_adj_13, n71764, n60646, n66463, 
            n34, n66240, n44122, n26732, n460, n39, n26478, \current[10] , 
            n66388, \current[9] , \current[8] , displacement, n27004, 
            n38, n486, n40, n66644, n67902, n66992, n67037, tx_active, 
            \pwm_counter[8] , n17, \pwm_counter[6] , n13, n66680, 
            n66842, n66625, n71771, n66244, n71769, n76, n78810, 
            n78642, n22_adj_14, n35278, \current[7] , \current[6] , 
            \current[5] , \current[4] , n78900, n66788, n68353, n66590, 
            n61349, n66150, n6, n66769, n27241, n71189, n66791, 
            n27201, n66751, n66555, n70983, n7_adj_15, n66660, n68099, 
            n45146, n14, n41543, n78834, n78498, tx_o, r_SM_Main, 
            \r_SM_Main_2__N_3536[1] , n29954, r_Clock_Count, \tx_data[3] , 
            n67642, n6_adj_16, \o_Rx_DV_N_3488[24] , n27, n29, \o_Rx_DV_N_3488[12] , 
            n23, n5218, n67002, tx_enable, baudrate, n28238, n67079, 
            \r_SM_Main[2]_adj_17 , r_Rx_Data, RX_N_2, n33, n34_adj_18, 
            n29935, n29934, n29932, n29913, n29912, n29908, n29904, 
            \o_Rx_DV_N_3488[8] , n5215, \r_SM_Main[1]_adj_19 , n28115, 
            r_Clock_Count_adj_28, n30760, n61786, n30756, \r_Bit_Index[0] , 
            \r_SM_Main_2__N_3446[1] , \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            n69006, n69649, n69585, n69665, n69633, n69601, n69617, 
            n69697, n69681, n69523) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[13] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    output [23:0]setpoint;
    input VCC_net;
    output [7:0]\data_in_frame[8] ;
    input clk16MHz;
    output \data_out_frame[3][3] ;
    input GND_net;
    output n2872;
    output [7:0]\data_out_frame[8] ;
    input n66000;
    input n65999;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    output n78804;
    output \data_out_frame[1][1] ;
    output \data_out_frame[3][1] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output n71810;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output n71808;
    output [7:0]rx_data;
    output n7;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[16] ;
    input n28715;
    input n65854;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output Kp_23__N_1748;
    input reset;
    output n8;
    input n65998;
    output \data_out_frame[1][7] ;
    output \data_out_frame[1][6] ;
    output [7:0]\data_in_frame[5] ;
    input n65997;
    input n66003;
    input n65996;
    output [7:0]\data_out_frame[9] ;
    input n66040;
    input n65995;
    input n65994;
    input n65993;
    input n65992;
    input n65991;
    input n65990;
    input n65989;
    output [7:0]\data_out_frame[10] ;
    input n65855;
    input n65988;
    input n65987;
    input n65986;
    input n65985;
    input n65984;
    output \FRAME_MATCHER.i[5] ;
    output \FRAME_MATCHER.i[4] ;
    output \FRAME_MATCHER.i[3] ;
    input n65983;
    input n65982;
    output [7:0]\data_out_frame[11] ;
    input n65981;
    input n65980;
    input n65979;
    input n65978;
    input n65977;
    input n65976;
    input n65975;
    input n65871;
    input n65973;
    input n65972;
    input n65971;
    input n65970;
    input n65969;
    input n65968;
    output \data_in_frame[1][0] ;
    input [23:0]encoder0_position;
    input n65967;
    output \data_out_frame[0][2] ;
    input n65966;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output n71801;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[16] ;
    output n71799;
    output n78768;
    input n65965;
    output \data_in_frame[0][0] ;
    output \data_in_frame[0][1] ;
    input [7:0]ID;
    output \data_in_frame[0][7] ;
    input n65964;
    input [23:0]pwm_setpoint;
    output \data_in_frame[0][6] ;
    output \data_in_frame[0][3] ;
    output \data_in_frame[0][5] ;
    output n66998;
    output \data_in_frame[2][4] ;
    output \data_out_frame[1][5] ;
    output \data_in_frame[2][6] ;
    input n65963;
    input n30143;
    output [7:0]\data_in_frame[4] ;
    output \data_in_frame[1][6] ;
    output \data_in_frame[2][0] ;
    output n51;
    input n30139;
    input n22;
    input \current[11] ;
    input n30136;
    input n30133;
    input \current[15] ;
    output n260;
    input n65728;
    output \data_out_frame[1][3] ;
    input n30130;
    input n30127;
    input n30124;
    input n30121;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_in_frame[17] ;
    output Kp_23__N_612;
    output rx_data_ready;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output n66982;
    output [7:0]\data_in_frame[18] ;
    output \data_in_frame[2][3] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[21] ;
    input n30093;
    output [23:0]deadband;
    input n30092;
    output \data_in_frame[2][1] ;
    output [7:0]\data_out_frame[20] ;
    input n30091;
    output [7:0]\data_out_frame[22] ;
    input n30090;
    input n30089;
    input n30088;
    input n30087;
    input n30086;
    input n30085;
    input n30084;
    input n30083;
    input n30082;
    input n30081;
    input n30080;
    output DE_c;
    input n30079;
    input n30078;
    output \data_out_frame[0][4] ;
    output \data_out_frame[3][4] ;
    input n30077;
    input n30076;
    input n30074;
    input n30073;
    input n30072;
    input n30071;
    output \data_out_frame[0][3] ;
    output n71763;
    input n30070;
    output [23:0]IntegralLimit;
    input n30069;
    input n30068;
    input n30066;
    input n30065;
    input n30064;
    input n30063;
    input n30062;
    input n30061;
    input n30060;
    input n30059;
    input n30058;
    input n30057;
    input n30056;
    input n30055;
    input n30054;
    input n65962;
    input n65961;
    input n65960;
    input n30053;
    input n65959;
    input n65958;
    input n30052;
    input n65957;
    input n65956;
    input n30051;
    input n30050;
    input n30049;
    input n30048;
    input n30047;
    output \Kp[1] ;
    input n65955;
    input n30046;
    output \Kp[2] ;
    input n30045;
    output \Kp[3] ;
    input n30044;
    output \Kp[4] ;
    input n30043;
    output \Kp[5] ;
    input n30042;
    output \Kp[6] ;
    input n65954;
    input n65953;
    input n65952;
    input n65951;
    input n65950;
    input n30041;
    output \Kp[7] ;
    input n30040;
    output \Kp[8] ;
    input n30039;
    output \Kp[9] ;
    input n65949;
    input n65948;
    output \Kp[10] ;
    input n30037;
    output \Kp[11] ;
    input n30036;
    output \Kp[12] ;
    input n65947;
    input n65946;
    input n65945;
    output \Kp[13] ;
    output n66594;
    input n30034;
    output \Kp[14] ;
    input n30033;
    output \Kp[15] ;
    input n30032;
    output \Ki[1] ;
    input n30031;
    output \Ki[2] ;
    input n30030;
    output \Ki[3] ;
    input n65944;
    input n65853;
    output [7:0]\data_in_frame[12] ;
    input n65943;
    input n65856;
    input n30029;
    output \Ki[4] ;
    input n30028;
    output \Ki[5] ;
    input n65942;
    input n30027;
    output \Ki[6] ;
    output LED_c;
    input n30026;
    output \Ki[7] ;
    input n65861;
    output [7:0]\data_in_frame[9] ;
    input n65865;
    input n65866;
    input n30025;
    output \Ki[8] ;
    input n30024;
    output \Ki[9] ;
    input n30023;
    output \Ki[10] ;
    input n65867;
    input n30022;
    output \Ki[11] ;
    input n65868;
    input n65869;
    input n65872;
    input n30021;
    output \Ki[12] ;
    input n65875;
    input n29286;
    input n65876;
    input n65877;
    input n30020;
    output \Ki[13] ;
    input n30019;
    output \Ki[14] ;
    input n30018;
    output \Ki[15] ;
    input n65878;
    input n65879;
    input n65880;
    input n65874;
    input n65881;
    input n65882;
    input n65883;
    output n26873;
    output n61123;
    input n65884;
    input n30005;
    input n30001;
    output [23:0]neopxl_color;
    input n74616;
    input n78618;
    input n7_adj_7;
    output [7:0]\data_in_frame[10] ;
    input n30000;
    input n29999;
    input n29998;
    input n29997;
    input n29996;
    input n29995;
    input n29994;
    output [7:0]\data_in_frame[11] ;
    input n29993;
    input n29992;
    input n29991;
    input n29990;
    input n74617;
    input n29989;
    input n29988;
    output [7:0]control_mode;
    output \control_mode[5] ;
    output \control_mode[6] ;
    output \control_mode[7] ;
    output \current_limit[1] ;
    output \current_limit[2] ;
    output \current_limit[3] ;
    output \current_limit[4] ;
    output \current_limit[5] ;
    input n29942;
    output [23:0]PWMLimit;
    output \current_limit[0] ;
    output \control_mode[0] ;
    input n29939;
    input n29938;
    output \Ki[0] ;
    input n29937;
    output \Kp[0] ;
    input n29936;
    input n29933;
    input n65885;
    input n65886;
    input n65887;
    input n65888;
    input n65889;
    input n65890;
    input n65891;
    input n65892;
    input n65893;
    input n65894;
    input n65895;
    input n65896;
    input n65897;
    input n65898;
    input n65899;
    input n65900;
    input n65901;
    input n65902;
    input n65903;
    input n65904;
    input n65905;
    input n65906;
    input n65907;
    input n65908;
    input n65909;
    input n7_adj_8;
    output n26329;
    output n8_adj_9;
    output [7:0]\data_in_frame[15] ;
    output [7:0]\data_in_frame[13] ;
    input n65910;
    input n29249;
    input n65911;
    input n65912;
    input n65913;
    input n65914;
    input n7_adj_10;
    input n7_adj_11;
    input n65873;
    input n66039;
    input n66038;
    output \data_out_frame[1][0] ;
    input n66037;
    input n66036;
    output \current_limit[8] ;
    output n66450;
    input n66166;
    input [23:0]encoder1_position;
    output n69038;
    output \current_limit[9] ;
    output \current_limit[10] ;
    input n65176;
    input n30770;
    input n65172;
    input n30766;
    input n30764;
    input n30761;
    input n65168;
    input n65164;
    input n29729;
    input n29732;
    input n30738;
    input n65160;
    input n30735;
    input n30734;
    input n30732;
    input n30731;
    input n30730;
    input n30728;
    input n30725;
    input n30723;
    input n30721;
    input n30720;
    input n30697;
    input n30679;
    input n30677;
    input n30676;
    input n30664;
    input n30663;
    input n66035;
    input n30631;
    input n30630;
    input n30629;
    input n30628;
    input n30247;
    input n30250;
    input n30624;
    input n30253;
    input n30622;
    input n30256;
    input n30259;
    input n30262;
    input n30617;
    input n30616;
    input n66034;
    input n29764;
    output \data_in_frame[20][0] ;
    input n29767;
    output \data_in_frame[20][1] ;
    input n29770;
    output \data_in_frame[20][2] ;
    input n65360;
    input n29777;
    output \data_in_frame[20][3] ;
    input n29780;
    output \data_in_frame[20][4] ;
    input n30265;
    input n30601;
    output \data_in_frame[10][0] ;
    output \data_in_frame[10][5] ;
    output \data_in_frame[10][6] ;
    input n30591;
    input n30587;
    input n30586;
    output \data_in_frame[10][7] ;
    input n30583;
    input n30294;
    input n30298;
    input n65336;
    input n30304;
    input n30308;
    input n65318;
    input n30314;
    input n30318;
    output \data_in_frame[13][6] ;
    output \data_in_frame[13][7] ;
    output [7:0]\data_in_frame[14] ;
    input n65863;
    input n65860;
    output \data_in_frame[14][4] ;
    output \data_in_frame[14][5] ;
    output \data_in_frame[14][6] ;
    output \data_in_frame[14][7] ;
    input n65154;
    input n30430;
    input n65150;
    input n65146;
    input n65094;
    input n65142;
    input n65244;
    input n30456;
    input n65276;
    input n65272;
    input n65268;
    input n30515;
    input n66033;
    input n29840;
    output [7:0]\data_in_frame[23] ;
    input n29843;
    input n29849;
    input n65134;
    input n29858;
    input n29861;
    input n65132;
    input n65130;
    input n29870;
    input n29874;
    input n29877;
    input n65398;
    input n66032;
    input n66031;
    output \data_out_frame[3][6] ;
    input n65870;
    output \data_out_frame[3][7] ;
    input n65864;
    input n66030;
    input n66029;
    input n66028;
    output n71789;
    output n71787;
    input n4938;
    input n66027;
    input n66026;
    input n66025;
    input n66024;
    input n60656;
    input n26758;
    input n66023;
    input n66022;
    input n66021;
    input n66020;
    input n66019;
    input n66018;
    input n65974;
    input n66017;
    input n66016;
    input n66015;
    input n66014;
    input n66013;
    output n71786;
    output n71784;
    input n66012;
    input n66011;
    input n66010;
    input n65915;
    input n65916;
    output \current_limit[6] ;
    input n65917;
    input n65918;
    input n65919;
    input n65920;
    input n65921;
    input n65922;
    input n65923;
    input n65924;
    input n65925;
    input n65926;
    input n65927;
    input n65928;
    input n65929;
    input n66009;
    output n23023;
    input n65862;
    input n66008;
    input n65859;
    input n65930;
    input n65931;
    input n65932;
    input n65933;
    input n65934;
    input n65935;
    input n65936;
    input n65937;
    input n65938;
    input n65939;
    input n65857;
    input n65940;
    input n65941;
    input n66007;
    input n66006;
    output \current_limit[7] ;
    input n66005;
    input n66004;
    input n66002;
    input \current[3] ;
    input n65858;
    input \current[2] ;
    input n66001;
    input \current[1] ;
    input \current[0] ;
    input n60808;
    input n7_adj_12;
    input n61318;
    input n68798;
    input n65754;
    output n25794;
    output n8_adj_13;
    output n71764;
    output n60646;
    output n66463;
    output n34;
    input n66240;
    output n44122;
    input n26732;
    input n460;
    output n39;
    input n26478;
    input \current[10] ;
    output n66388;
    input \current[9] ;
    input \current[8] ;
    input [23:0]displacement;
    output n27004;
    input n38;
    input n486;
    output n40;
    output n66644;
    output n67902;
    output n66992;
    output n67037;
    output tx_active;
    input \pwm_counter[8] ;
    output n17;
    input \pwm_counter[6] ;
    output n13;
    input n66680;
    output n66842;
    output n66625;
    output n71771;
    output n66244;
    output n71769;
    output n76;
    input n78810;
    input n78642;
    output n22_adj_14;
    output n35278;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    output n78900;
    output n66788;
    input n68353;
    output n66590;
    input n61349;
    output n66150;
    input n6;
    output n66769;
    output n27241;
    input n71189;
    input n66791;
    output n27201;
    output n66751;
    output n66555;
    input n70983;
    output n7_adj_15;
    output n66660;
    input n68099;
    output n45146;
    output n14;
    output n41543;
    output n78834;
    output n78498;
    output tx_o;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    input n29954;
    output [8:0]r_Clock_Count;
    input \tx_data[3] ;
    input n67642;
    output n6_adj_16;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n29;
    output \o_Rx_DV_N_3488[12] ;
    output n23;
    input n5218;
    input n67002;
    output tx_enable;
    input [31:0]baudrate;
    output n28238;
    output n67079;
    output \r_SM_Main[2]_adj_17 ;
    output r_Rx_Data;
    input RX_N_2;
    output n33;
    output n34_adj_18;
    input n29935;
    input n29934;
    input n29932;
    input n29913;
    input n29912;
    input n29908;
    input n29904;
    output \o_Rx_DV_N_3488[8] ;
    input n5215;
    output \r_SM_Main[1]_adj_19 ;
    output n28115;
    output [7:0]r_Clock_Count_adj_28;
    input n30760;
    input n61786;
    input n30756;
    output \r_Bit_Index[0] ;
    input \r_SM_Main_2__N_3446[1] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n69006;
    output n69649;
    output n69585;
    output n69665;
    output n69633;
    output n69601;
    output n69617;
    output n69697;
    output n69681;
    input n69523;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2, n30241, n2_adj_5308, n30238, n30235, n28325, n28649;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n59509, n74525, n28327, n59508, n74524, n28329, n59507, 
        n74523, n2_adj_5309, n2_adj_5310, n30232, n28331, n59506, 
        n74520, n28335, n59505, n74517, n28337, n59504, n74509, 
        n28339, n59503, n74487;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n78801, n28398, n71809;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n65402, n65400, n30229, n30226, n30223, n30220, n30217;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n29951, n30213, n30210, n30207, n30204, n30201, n30198, 
        n30195, \FRAME_MATCHER.i_31__N_2507 , n29960, n30191, n30188, 
        n30185, n30182, n30179, n30176, n28341, n59502, n74486, 
        n78795, n2_adj_5311, n28343, n59501, n74469, n30446, n30443, 
        n78798, n28345, n59500, n74468, n28347, n59499, n74467, 
        n28349, n59498, n74465, n28351, n59497, n74463, n28353, 
        n59496, n74448, n28355, n59495, n74447, n28357, n59494, 
        n74446, n28359, n59493, n74440, n30173, n2_adj_5312, n78789, 
        n71834, n28361, n59492, n74439, n2066, n28363, n59491, 
        n74435, n66156;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    
    wire n29886;
    wire [23:0]n4930;
    
    wire n28129, n2_adj_5313, n30170, n28365, n59490, n74434, n28367, 
        n59489, n74433, n2_adj_5314, n2_adj_5315, n28369, n59488, 
        n74430, n28371, n59487, n74427, n28373, n59486, n74422, 
        n30167, n2_adj_5316, n2_adj_5317, n2_adj_5318, n2_adj_5319, 
        n28375, n59485, n74421, n2_adj_5320, n2_adj_5321, n2_adj_5322, 
        n2_adj_5323, n2_adj_5324, n2_adj_5325, n2_adj_5326, n2_adj_5327, 
        n2_adj_5328, n2_adj_5329, n2_adj_5330, n2_adj_5331, n2_adj_5332, 
        n28377, n59484, n74417, n28379, n59483, n74415, n28381, 
        n59482, n74414, n28383, n59481, n74411, n28385, n59480, 
        n74410, n28387, n59479, n74409;
    wire [31:0]n133;
    
    wire n161, n2_adj_5333, n2_adj_5334, n2_adj_5335, n2_adj_5336, 
        n2_adj_5337, n2_adj_5338, n2_adj_5339, n2_adj_5340, n2_adj_5341, 
        n2_adj_5342, n2_adj_5343, n2_adj_5344, n2_adj_5345, n2_adj_5346, 
        n2_adj_5347, n2_adj_5348, n29883, n2_adj_5349, n2_adj_5350, 
        n30164, n74621, n2_adj_5351, n78771, n71800, n78774, n78765, 
        n78828, n74612, n78504, n76680, n2_adj_5352;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(99[12:25])
    
    wire n26750, n12, n30161, n30158, n30155, n30152, n30149, 
        n2_adj_5353, n30146, n78822, n74610, n78738, n78528, n76800, 
        n2_adj_5354, n2_adj_5355, n7_adj_5356, n10, n2_adj_5357, n2_adj_5358, 
        n2_adj_5359, n2_adj_5360, n2_adj_5361, n11;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    
    wire n65224, n29786, n9, n65218, n69189, n2_adj_5362, Kp_23__N_748, 
        n66309, n2_adj_5363, n2_adj_5364, n66267, n66417, Kp_23__N_753, 
        n66359, n2_adj_5365, n2_adj_5366, n27046, n10_adj_5367, n23_c, 
        n27_c, n2_adj_5368, n29978, n26;
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    
    wire n71103, n65, n26188, n29_c, n74457, n22_adj_5369, n31, 
        n71370, n78759, n71867, n78753, n78756, n78747, n78600;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n78735, n78723, n78726, n2_adj_5370, n2_adj_5371, n30118, 
        n66444, n3, n68828, n6_c, n60670, n3_adj_5372, n66546, 
        n3_adj_5373, n66381, n66416, n61341, n3_adj_5374, n3474, 
        n30002, n30007, n30012, n69031, n3_adj_5375, n30095, n66339, 
        n66710, n3_adj_5376, n66348, n66716, n60565, n60666, n66772, 
        n66474, n20, n66413, n26201, n66518, n19, n30015, n60585, 
        n26659, n60698, n21, n25417, n61545, n16, n61568, n61315, 
        n17_c, n60677, n26605, n66797, n66745, n66572, n66845, 
        n10_adj_5377;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    
    wire n66552, n69046, n12_adj_5378, n68518, n61070, n26526, n66707, 
        n5, n82, n66099, n3_adj_5379, n61587, n66515, n3_adj_5380, 
        n61643, n61306, n61603, n66108, tx_transmit_N_3416, \FRAME_MATCHER.i_31__N_2511 , 
        n1, n6_adj_5381, n66131, n27316, n2_adj_5382, n71760, n30075, 
        n1_adj_5383, n71829, n71830, n66672, n66824, n10_adj_5384, 
        n71899, n71898, n71826, n71827, n30067, n25877, n5_adj_5385, 
        n71836, n71835, n71847, n71848, n71857, n71856, n71874, 
        n71875, n71776, n71775, n60757;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n70933, n71913, n66333, n3_adj_5386, n71914, n71917, n71916, 
        n10_adj_5387, n71868, n71869, n6_adj_5388, n2_adj_5389, n2_adj_5390, 
        n2_adj_5391, n2_adj_5392, n2_adj_5393, n71803, n71802, n65839, 
        n65841, n65842, n65843, n65844, n65837, n65845, n65836, 
        n65840, n30038, n65846, n65847, n65848, n2_adj_5394, n65849, 
        n65838, n66276, Kp_23__N_767, n2_adj_5395, n2_adj_5396, n30035, 
        n65850, n65851, n61751, n6_adj_5397, n27157, n70901, n2_adj_5398, 
        n2_adj_5399, n28670, n65378, n65432, n66216, n2_adj_5400, 
        n2_adj_5401, n65434, n66264, n6_adj_5402, n2_adj_5403, n66689, 
        Kp_23__N_772, Kp_23__N_872, LED_N_3408, LED_N_3407, n27768, 
        \FRAME_MATCHER.i_31__N_2513 , n29209, n2_adj_5404, n3_adj_5405, 
        n5_adj_5406, n24043, n24272, n66763, n66719, n2_adj_5407, 
        n2_adj_5408, n66352, n2_adj_5409, n2_adj_5410, n2_adj_5411, 
        n2_adj_5412, n2_adj_5413, n2_adj_5414, n2_adj_5415, n2_adj_5416, 
        n2_adj_5417, n2_adj_5418, n25456, n66549, n2_adj_5419, n2_adj_5420, 
        n2_adj_5421, n2_adj_5422, n2_adj_5423, n26416, n61589, n2_adj_5424;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n30632;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n29949, n26424, n30662, n76856, n79011, n71295, n68582, 
        n3_adj_5426, n30661, n30660, n68633, n66863, n66584, n66698, 
        n26685, n26957, Kp_23__N_974, n30659, n30658, n30657, n30656;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n30655, n24039, n6_adj_5427, n76854, n79005, n30653, n61765, 
        n3_adj_5428, n30652, n30651, n29987, n53030;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(246[14:26])
    
    wire n29985, n29983, n29982, n29981, n29977, n29974, n29973, 
        n29972, n29971, n29970, n29941, n29940, Kp_23__N_993, n66312, 
        n66695, n71181, n66739, n10_adj_5429, n2_adj_5430, n3_adj_5431, 
        n30650, n2_adj_5432, n2_adj_5433, n2_adj_5434, n2_adj_5435, 
        n2_adj_5436, n2_adj_5437, n2_adj_5438, n2_adj_5439, n2_adj_5440, 
        n2_adj_5441, n2_adj_5442, n2_adj_5443, n2_adj_5444, n2_adj_5445, 
        n2_adj_5446, n2_adj_5447, n2_adj_5448, n2_adj_5449, n2_adj_5450, 
        n2_adj_5451, n2_adj_5452, n2_adj_5453, n2_adj_5454, n2_adj_5455, 
        n30649, n78594, n30648, n26244, n26846, n66860, n28323, 
        n30647, n60664, n66666, n66827, n26343, n26362, n66212, 
        n2_adj_5458, n2_adj_5459, n2_adj_5460, n26378, n2_adj_5461, 
        n2_adj_5462, n2_adj_5463, n30646, n76848, n74635, n78987, 
        n78624, n76846, n74611, n78975, n78606, n2_adj_5466, n2_adj_5467, 
        n2_adj_5468, n7_adj_5469, n68344, n26743, n26827, n68553, 
        n66447, n12_adj_5470, n30645, n66391, n66574, n66378, n30644, 
        n66734, n12_adj_5471, n30643, n60778, n14_c, n2_adj_5472, 
        n2_adj_5473, n30784, n30642, n61533, n66748, n22_adj_5474, 
        n21_adj_5475, n60763, n23_adj_5476, n30641, n16_adj_5477, 
        n30640, n66491, n60624, n22_adj_5478, n30639, n30638, n30637, 
        n30636, n30635, n60581, n24, n30634, n30633, n30654, n20_adj_5479, 
        n60607, n66692, n10_adj_5480, n66497, n30783, n30779, n66587, 
        n66531, n60780, n10_adj_5481, n37697, n30777, n30776, n30775, 
        n30773, n30772, n30771, n30768, n29738, n29741, n29744, 
        n29747, n29750, n66571, n29754, n28674;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(99[12:25])
    
    wire n65364, n29757, n29761, n29792;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    
    wire n29795, n29798, n29801, n30268, n30271, n30278, n65368, 
        n30284, n30288, n29804, n29807, n30291, n29810, n29813, 
        n30321, n29816, n30324, n30337, n30340, n30344, n30347, 
        n30350, n30353, n30357, n30360;
    wire [7:0]\data_in_frame[13]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30363, n30366, n30370, n30373, n30376, n30380, n30383;
    wire [7:0]\data_in_frame[14]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30386, n30390, n30393, n30396, n30400, n30403, n30406, 
        n30410, n15, n30416, n30420, n30423, n29819, n29822, n29825, 
        n29828, n29831, n29834, n29837, n61555, n29889, n29892, 
        n60269, n61645, n29895, n29898, n29901, n29905, n29909, 
        n66231, n7_adj_5482, n29914, n61607, n66604, n29917, n29920, 
        n66528, n29923, n2_adj_5483, n2_adj_5484, n2_adj_5485, n2_adj_5486, 
        n66453, n1720, n68559, n68131, n26537, n61678, n66488, 
        n29926, n29929, n2_adj_5487, n2_adj_5488, n66794, n66608, 
        n12_adj_5489, n71788, n28441, n24165, n79076, n61308, n66524, 
        n27427, \FRAME_MATCHER.i_31__N_2508 , n2046, n2047, n20637, 
        n65018, \FRAME_MATCHER.i_31__N_2512 , n2058, n27430, \FRAME_MATCHER.i_31__N_2514 , 
        n26870, n61658, n66776, n2_adj_5490, n61605, n2_adj_5491, 
        n2_adj_5492, n2_adj_5493, n66495, n78648, n66568, n71177, 
        n6_adj_5494, n71059, n2_adj_5495, n2_adj_5496, n2_adj_5497, 
        n2_adj_5498, n2_adj_5499, n2_adj_5500, n2_adj_5501, n2_adj_5502, 
        n2_adj_5503, n2_adj_5504, n2_adj_5505, n2_adj_5506, n61240, 
        n10_adj_5507, n44101, n68457, n66683, n71785, n26583, n68646, 
        n61528, n25588, n66407, n60640, n10_adj_5508, n60658, n2_adj_5509, 
        n2_adj_5510, n26722, Kp_23__N_799, n2_adj_5511, n78852, n2_adj_5512, 
        n1835, n26941, n10_adj_5513, n2_adj_5514, n78564, n29753, 
        n2_adj_5515, n2_adj_5516, n2_adj_5517, n2_adj_5518, n2_adj_5519, 
        n2_adj_5520, n2_adj_5521, n2_adj_5522, n2_adj_5523, n2_adj_5524, 
        n2_adj_5525, n2_adj_5526, n2_adj_5527, n2_adj_5528, n61749, 
        n71157, n2_adj_5529, n2_adj_5530, n2_adj_5531, n2_adj_5532, 
        n2_adj_5533, n2_adj_5534, n2_adj_5535, n2_adj_5536, n2_adj_5537, 
        n2_adj_5538, n2_adj_5539, n2_adj_5540, n2_adj_5541, n2_adj_5542, 
        n2_adj_5543, n2_adj_5544, n3_adj_5545, n3_adj_5546, n3_adj_5547, 
        n3_adj_5548, n29199;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n29193, n1_adj_5549;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n65830, n1_adj_5550, n65831, n29725, n1_adj_5551, n65827, 
        n60687, n66435, n10_adj_5552, n66562, n12_adj_5553, n1_adj_5554, 
        n65832, n61543, n26898, n1_adj_5555, n65828, n1_adj_5556, 
        n65833, n1_adj_5557, n65834, n60291, n66616, n1_adj_5558, 
        n65829, n66597, n61601, n78921, n66438, n5_adj_5559, n66356, 
        n26087, n9_adj_5560, n68678, n66851, n66725, n20_adj_5561, 
        n26058, n26459, n66809, n19_adj_5562, n61358, n21_adj_5563, 
        n27087, n26781, n1699, n66521, n26617, n6_adj_5564, n78588, 
        n6_adj_5566, n66669, n66196, n27192, n66806, n10_adj_5567, 
        n771, n25857, n4, n61760, n27182, n6_adj_5568, n68217, 
        n78915, n71761, n78909, n60767, n66103, n60988, n18, n60810, 
        n19_adj_5570, n12_adj_5571, n68158, n58266, n65826, n58265, 
        n28, n26_adj_5572, n66821, n27_adj_5573, n25, n61583, n66619, 
        n58264, n58263, n58262, n58261, n58260, n66206, n66628, 
        n66760, n14_adj_5574, n66728, n13_c, n27256, n66779, n7_adj_5575, 
        n60592, n60445, n18_adj_5576, n66641, n66181, n66800, n10_adj_5577, 
        n66190, n27290, n66757, n66836, n66803, n6_adj_5578, n66866, 
        n10_adj_5579, n66622, n66647, n12_adj_5580, n26811, n6_adj_5581, 
        n66503, n66504, n66251, n6_adj_5582, n1668, n1130, n12_adj_5583, 
        n27211, n26062, n66372, n10_adj_5584, n66304, n29_adj_5585, 
        n10_adj_5586, n66375, n66631, n66742, n10_adj_5587, n66200, 
        n66654, n6_adj_5588, n1516, n26067, n66228, n66782, n10_adj_5589, 
        n66839, n66611, n26051, n66342, n24_adj_5590, n17_adj_5591, 
        n66818, n22_adj_5592, n26_adj_5593, n10_adj_5594, n66441, 
        n14_adj_5595, n69125, n68714, n12_adj_5596, n66169, n61520, 
        n61566, n27056, n10_adj_5597, n14_adj_5598, n6_adj_5599, n1193, 
        n16_adj_5600, n66812, n17_adj_5601, n60693, n66325, n40_adj_5602, 
        n68749, n26910, n30, n28_adj_5603, n29_adj_5604, n26473, 
        n27_adj_5605, n68184, n14_adj_5606, n13_adj_5607, n26590, 
        n68332, n26309, n8_adj_5608, n6_adj_5609, n8_adj_5610, n66650, 
        n66704, n6_adj_5611, n10_adj_5612, n14_adj_5613, n6_adj_5614, 
        n6_adj_5615, n8_adj_5616, n45273, n68152, n1949, n1952, 
        n25866, n4452, n1955, n68081, n67901, n66318, n61665, 
        n66481, n69075, n66254, n26315, n27050, n26716, n66815, 
        n6_adj_5619, n26673, n66686, n26719, n66362, n78864, n78546, 
        n66394, n18_adj_5620, n66701, n26816, n4_adj_5621, n78897, 
        n71165, n66301, n27115, n61180, n66479, n71770, n70987, 
        n18_adj_5622, n27_adj_5623, n61599, n10_adj_5624, n66163, 
        n66459, n66512, n8_adj_5625, n25479, n71109, n70891, n66248, 
        n66485, n66634, n68740, n60648, n71115, Kp_23__N_1564, n66486, 
        n66713, n66369, n66577, n71253, n71259, n66833, n66273, 
        n71217, n71223, n71229, n14_adj_5627, n66538, n60628, n71233, 
        n66429, n66336, n71239, n26522, n66193, n71243, n68427, 
        n66558, n66785, n68895, n66384, n61660, n20_adj_5628, n6_adj_5629, 
        n26794, n27043, n66494, n66500, n66329, n71075, n7_adj_5631, 
        n26843, Kp_23__N_1067, Kp_23__N_1389, n71081, n77669, n71087, 
        n66580, n28088, n8_adj_5632, Kp_23__N_1607, n6_adj_5633, n68908, 
        n25505, n66432, n77665, n61577, n66677, n71065, n30_adj_5634, 
        n66279, n71281, n71285, n61525, n10_adj_5635, n66857, n14_adj_5636, 
        Kp_23__N_1256, n78645, n66535, n61778, n24_adj_5637, n22_adj_5638, 
        n66830, n26_adj_5639, n66722, n66456, n24_adj_5640, n61328, 
        n22_adj_5641, n26_adj_5642, n27071, n66401, n24268, n26098, 
        n70977, n66315, n70985, n70993, n70999, n66565, n66322, 
        n71005, n66854, n6_adj_5643, n18_adj_5644, n19_adj_5645, n60723, 
        n25467, n71171, n66754, n78861, n26321, n66219, n71265, 
        n78633, n27223, n26280, n26777, n61449, n6_adj_5647, n6_adj_5648, 
        n6_adj_5649, n78636, n26294, Kp_23__N_869, n14_adj_5650, n66420, 
        n15_adj_5651, n66209, n26306, n66286, n12_adj_5652, n7_adj_5653, 
        n66397, n66470, n26137, n26297, n66365, n26284, n66175, 
        n78849, n6_adj_5655, n69112, n66404, n26266, n78840, n76803, 
        n78540, n66657, n71027, n71025, n71023, n71037, n71035, 
        n71041, n71049, n71051, n15_adj_5656, n69110, n21_adj_5657, 
        n27_adj_5658, n26_adj_5659, n71362, n71486, n31_adj_5660, 
        n12_adj_5661, n6_adj_5662, n8_adj_5663, n68484, n70941, n66430, 
        n78621, n68439, n68725, n20632, n8_adj_5664, n70947, n66261, 
        n70949, n6_adj_5665, n70951, n23015, n71153, n3303, n68677, 
        n71149, n71123, n67899, n70953, n68042, n70959, n70961, 
        n68851, n71127, n70965, n71310, n68441, n66732, n1953, 
        n25747, n27992, n68490, n78603, n78597, n10_adj_5666, n68362, 
        n14_adj_5667, n68038, n14_adj_5668, n13_adj_5669, n20_adj_5670, 
        n13_adj_5671, n18_adj_5672, n22_adj_5673, n25913, n16_adj_5674, 
        n17_adj_5675, n25954, n10_adj_5676, n14_adj_5677, n25907, 
        n20_adj_5678, n25777, n19_adj_5679, n71490, n78591, n71389, 
        n18_adj_5680, n19_adj_5681, n14_adj_5682, n15_adj_5683, n16_adj_5684, 
        n17_adj_5685, n66134, n4_adj_5686, n4_adj_5687, n6_adj_5688, 
        n78585, n78837, n78831, n78561, n78825, n78819, n78543, 
        n78537, n78525, n78501, n78495;
    
    SB_LUT4 select_787_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30241));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30238));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30235));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_33_lut  (.I0(n74525), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n59509), .O(n28325)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_32_lut  (.I0(n74524), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n59508), .O(n28327)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_32  (.CI(n59508), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n59509));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_31_lut  (.I0(n74523), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n59507), .O(n28329)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_31  (.CI(n59507), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n59508));
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5309), .S(n66000));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5310), .S(n65999));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30232));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_30_lut  (.I0(n74520), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n59506), .O(n28331)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_30  (.CI(n59506), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n59507));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_29_lut  (.I0(n74517), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n59505), .O(n28335)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_29  (.CI(n59505), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n59506));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_28_lut  (.I0(n74509), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n59504), .O(n28337)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_28  (.CI(n59504), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n59505));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_27_lut  (.I0(n74487), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n59503), .O(n28339)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62913 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n78801));
    defparam byte_transmit_counter_0__bdd_4_lut_62913.LUT_INIT = 16'he4aa;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_27  (.CI(n59503), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n59504));
    SB_LUT4 n78801_bdd_4_lut (.I0(n78801), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n78804));
    defparam n78801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14187_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n28398));   // verilog/coms.v(109[34:55])
    defparam i14187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55974_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71809));
    defparam i55974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55975_4_lut (.I0(n71809), .I1(n28398), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n71810));
    defparam i55975_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i55973_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71808));
    defparam i55973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61822_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[0] [4]), .I2(n7), 
            .I3(GND_net), .O(n65402));   // verilog/coms.v(94[13:20])
    defparam i61822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61821_3_lut (.I0(rx_data[2]), .I1(\data_in_frame[0] [2]), .I2(n7), 
            .I3(GND_net), .O(n65400));   // verilog/coms.v(94[13:20])
    defparam i61821_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30229));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30226));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30223));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30220));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30217));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
           .D(n29951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30213));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30210));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30204));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30201));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30198));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30195));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59743_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74517));   // verilog/coms.v(158[12:15])
    defparam i59743_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
           .D(n29960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30191));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30188));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30185));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30182));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30179));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30176));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_26_lut  (.I0(n74486), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n59502), .O(n28341)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_26  (.CI(n59502), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n59503));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62908 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n78795));
    defparam byte_transmit_counter_0__bdd_4_lut_62908.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_25_lut  (.I0(n74469), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n59501), .O(n28343)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i16234_3_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(n28715), .I3(GND_net), .O(n30446));   // verilog/coms.v(130[12] 305[6])
    defparam i16234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16231_3_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(n28715), .I3(GND_net), .O(n30443));   // verilog/coms.v(130[12] 305[6])
    defparam i16231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n78795_bdd_4_lut (.I0(n78795), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n78798));
    defparam n78795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_25  (.CI(n59501), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n59502));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_24_lut  (.I0(n74468), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n59500), .O(n28345)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_24  (.CI(n59500), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n59501));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_23_lut  (.I0(n74467), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n59499), .O(n28347)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_23  (.CI(n59499), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n59500));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_22_lut  (.I0(n74465), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n59498), .O(n28349)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_22  (.CI(n59498), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n59499));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_21_lut  (.I0(n74463), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n59497), .O(n28351)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_21  (.CI(n59497), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n59498));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_20_lut  (.I0(n74448), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n59496), .O(n28353)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_20  (.CI(n59496), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n59497));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_19_lut  (.I0(n74447), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n59495), .O(n28355)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_19  (.CI(n59495), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n59496));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_18_lut  (.I0(n74446), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n59494), .O(n28357)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_18  (.CI(n59494), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n59495));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_17_lut  (.I0(n74440), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n59493), .O(n28359)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30173));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5312), .S(n65854));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62903 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n78789));
    defparam byte_transmit_counter_0__bdd_4_lut_62903.LUT_INIT = 16'he4aa;
    SB_LUT4 n78789_bdd_4_lut (.I0(n78789), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71834));
    defparam n78789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_17  (.CI(n59493), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n59494));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_16_lut  (.I0(n74439), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n59492), .O(n28361)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2066), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_16  (.CI(n59492), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n59493));
    SB_LUT4 i59074_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74520));   // verilog/coms.v(158[12:15])
    defparam i59074_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_15_lut  (.I0(n74435), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n59491), .O(n28363)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i15674_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29886));
    defparam i15674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n28129), 
            .D(n4930[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5313), .S(n65998));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30170));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_15  (.CI(n59491), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n59492));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_14_lut  (.I0(n74434), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n59490), .O(n28365)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_14  (.CI(n59490), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n59491));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_13_lut  (.I0(n74433), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n59489), .O(n28367)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[1][7] ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5314));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_3_lut_adj_1070 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[1][6] ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5315));
    defparam i1_3_lut_adj_1070.LUT_INIT = 16'ha8a8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_13  (.CI(n59489), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n59490));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_12_lut  (.I0(n74430), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n59488), .O(n28369)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_12  (.CI(n59488), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n59489));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_11_lut  (.I0(n74427), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n59487), .O(n28371)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_11  (.CI(n59487), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n59488));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_10_lut  (.I0(n74422), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n59486), .O(n28373)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30167));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_10  (.CI(n59486), .I0(n28649), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n59487));
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5316), .S(n65997));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5317), .S(n66003));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5318), .S(n65996));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5319), .S(n66040));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_9_lut  (.I0(n74421), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n59485), .O(n28375)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5320), .S(n65995));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5321), .S(n65994));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5322), .S(n65993));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5323), .S(n65992));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5324), .S(n65991));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5325), .S(n65990));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5326), .S(n65989));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5327), .S(n65855));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5328), .S(n65988));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5329), .S(n65987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5330), .S(n65986));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5331), .S(n65985));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5332), .S(n65984));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_9  (.CI(n59485), .I0(n28649), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n59486));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_8_lut  (.I0(n74417), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n59484), .O(n28377)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_8  (.CI(n59484), .I0(n28649), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n59485));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_7_lut  (.I0(n74415), .I1(n28649), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n59483), .O(n28379)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_7  (.CI(n59483), .I0(n28649), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n59484));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_6_lut  (.I0(n74414), .I1(n28649), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n59482), .O(n28381)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_6  (.CI(n59482), .I0(n28649), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n59483));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_5_lut  (.I0(n74411), .I1(n28649), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n59481), .O(n28383)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_5  (.CI(n59481), .I0(n28649), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n59482));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_4_lut  (.I0(n74410), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n59480), .O(n28385)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_4  (.CI(n59480), .I0(n28649), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n59481));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_3_lut  (.I0(n74409), .I1(n28649), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n59479), .O(n28387)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_3  (.CI(n59479), .I0(n28649), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n59480));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n59479));
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5333), .S(n65983));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5334), .S(n65982));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5335), .S(n65981));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5336), .S(n65980));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5337), .S(n65979));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5338), .S(n65978));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5339), .S(n65977));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5340), .S(n65976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5341), .S(n65975));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5342), .S(n65871));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5343), .S(n65973));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5344), .S(n65972));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5345), .S(n65971));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5346), .S(n65970));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5347), .S(n65969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5348), .S(n65968));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15671_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[1][0] ), .O(n29883));
    defparam i15671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5350), .S(n65967));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30164));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59183_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n74621));
    defparam i59183_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5351), .S(n65966));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62898 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n78771));
    defparam byte_transmit_counter_0__bdd_4_lut_62898.LUT_INIT = 16'he4aa;
    SB_LUT4 i55965_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71800));
    defparam i55965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55966_4_lut (.I0(n71800), .I1(n74621), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n71801));
    defparam i55966_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 n78771_bdd_4_lut (.I0(n78771), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n78774));
    defparam n78771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i55964_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71799));
    defparam i55964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62884 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n78765));
    defparam byte_transmit_counter_0__bdd_4_lut_62884.LUT_INIT = 16'he4aa;
    SB_LUT4 n78765_bdd_4_lut (.I0(n78765), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n78768));
    defparam n78765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59276_2_lut (.I0(n78828), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74612));
    defparam i59276_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i60845_3_lut (.I0(n78774), .I1(n78504), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76680));
    defparam i60845_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5352), .S(n65965));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[2]_c [2]), .I1(\data_in_frame[0][0] ), 
            .I2(\data_in_frame[0][1] ), .I3(GND_net), .O(n26750));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut (.I0(ID[7]), .I1(ID[1]), .I2(\data_in_frame[0][7] ), 
            .I3(\data_in_frame[0][1] ), .O(n12));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30161));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30158));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30155));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30152));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30149));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5353), .S(n65964));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30146));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59480_2_lut (.I0(n78822), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74610));
    defparam i59480_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i60965_3_lut (.I0(n78738), .I1(n78528), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76800));
    defparam i60965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [7]), 
            .I2(encoder0_position[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [0]), 
            .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n7_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'ha088;
    SB_LUT4 i2_4_lut (.I0(ID[3]), .I1(\data_in_frame[0][6] ), .I2(\data_in_frame[0][3] ), 
            .I3(ID[6]), .O(n10));   // verilog/coms.v(99[12:25])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 select_787_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[0][5] ), .I1(ID[2]), .I2(ID[5]), 
            .I3(\data_in_frame[0] [2]), .O(n11));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i61816_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[20] [7]), 
            .I2(n66998), .I3(GND_net), .O(n65224));   // verilog/coms.v(94[13:20])
    defparam i61816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15574_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n66998), .I3(GND_net), .O(n29786));   // verilog/coms.v(130[12] 305[6])
    defparam i15574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(ID[4]), .I1(\data_in_frame[0][0] ), .I2(\data_in_frame[0] [4]), 
            .I3(ID[0]), .O(n9));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'h7bde;
    SB_LUT4 i61815_3_lut (.I0(rx_data[5]), .I1(\data_in_frame[20] [5]), 
            .I2(n66998), .I3(GND_net), .O(n65218));   // verilog/coms.v(94[13:20])
    defparam i61815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n11), .I2(n10), .I3(n12), .O(n69189));   // verilog/coms.v(99[12:25])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 select_787_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[0][0] ), .I1(Kp_23__N_748), .I2(GND_net), 
            .I3(GND_net), .O(n66309));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[0][3] ), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66267));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n66417));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_0__7__I_0_4044_2_lut (.I0(\data_in_frame[0][7] ), 
            .I1(\data_in_frame[0][6] ), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_753));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_0__7__I_0_4044_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\data_in_frame[2][4] ), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66359));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1076 (.I0(Kp_23__N_753), .I1(n66417), .I2(n66267), 
            .I3(\data_in_frame[0][5] ), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1077 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [2]), 
            .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1077.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_adj_1078 (.I0(\data_in_frame[2][6] ), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0][5] ), .I3(GND_net), .O(n27046));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1078.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5365), .S(n65963));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_2035_i10_2_lut (.I0(\data_in_frame[0][7] ), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5367));   // verilog/coms.v(169[9:87])
    defparam equal_2035_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut (.I0(n27046), .I1(\data_in_frame[0][7] ), .I2(\data_in_frame[1][0] ), 
            .I3(\data_in_frame[0][6] ), .O(n23_c));
    defparam i6_4_lut.LUT_INIT = 16'h4114;
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30143));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i10_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1][6] ), .O(n27_c));
    defparam i10_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 select_787_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n29978));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut (.I0(\data_in_frame[2][0] ), .I1(n10_adj_5367), .I2(n66309), 
            .I3(\data_in_frame[1] [5]), .O(n26));
    defparam i9_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(current_limit[14]), .I1(current_limit[12]), 
            .I2(GND_net), .I3(GND_net), .O(n71103));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(current_limit[15]), .I1(n71103), .I2(n65), 
            .I3(current_limit[13]), .O(n51));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'h5554;
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30139));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i12_4_lut (.I0(n23_c), .I1(\data_in_frame[1] [7]), .I2(n26188), 
            .I3(n66309), .O(n29_c));
    defparam i12_4_lut.LUT_INIT = 16'h0208;
    SB_LUT4 i65_3_lut (.I0(n22), .I1(\current[11] ), .I2(current_limit[11]), 
            .I3(GND_net), .O(n65));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i65_3_lut.LUT_INIT = 16'hb2b2;
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30136));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59010_4_lut (.I0(current_limit[14]), .I1(n65), .I2(current_limit[13]), 
            .I3(current_limit[12]), .O(n74457));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i59010_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i14_4_lut (.I0(n27_c), .I1(n69189), .I2(n22_adj_5369), .I3(n26750), 
            .O(n31));
    defparam i14_4_lut.LUT_INIT = 16'h0020;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30133));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i23533_4_lut (.I0(n51), .I1(n74457), .I2(\current[15] ), .I3(current_limit[15]), 
            .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i23533_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 select_787_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16_4_lut (.I0(n31), .I1(n29_c), .I2(n71370), .I3(n26), 
            .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62879 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n78759));
    defparam byte_transmit_counter_0__bdd_4_lut_62879.LUT_INIT = 16'he4aa;
    SB_LUT4 n78759_bdd_4_lut (.I0(n78759), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71867));
    defparam n78759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62874 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n78753));
    defparam byte_transmit_counter_0__bdd_4_lut_62874.LUT_INIT = 16'he4aa;
    SB_LUT4 n78753_bdd_4_lut (.I0(n78753), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n78756));
    defparam n78753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63008 (.I0(byte_transmit_counter[3]), 
            .I1(n76680), .I2(n74612), .I3(byte_transmit_counter[4]), .O(n78747));
    defparam byte_transmit_counter_3__bdd_4_lut_63008.LUT_INIT = 16'he4aa;
    SB_LUT4 n78747_bdd_4_lut (.I0(n78747), .I1(n78600), .I2(n65728), .I3(byte_transmit_counter[4]), 
            .O(tx_data[2]));
    defparam n78747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62860 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n78735));
    defparam byte_transmit_counter_0__bdd_4_lut_62860.LUT_INIT = 16'he4aa;
    SB_LUT4 n78735_bdd_4_lut (.I0(n78735), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n78738));
    defparam n78735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62850 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n78723));
    defparam byte_transmit_counter_0__bdd_4_lut_62850.LUT_INIT = 16'he4aa;
    SB_LUT4 n78723_bdd_4_lut (.I0(n78723), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n78726));
    defparam n78723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30130));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30127));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30124));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59041_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74487));   // verilog/coms.v(158[12:15])
    defparam i59041_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30121));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30118));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_223_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n66444), .I3(\data_out_frame[25] [5]), 
            .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_222_i3_4_lut (.I0(n68828), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_c), .I3(n60670), .O(n3_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2872));   // verilog/coms.v(94[13:20])
    defparam i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 select_787_Select_221_i3_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n66546), .I3(\data_out_frame[25] [4]), 
            .O(n3_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_221_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 mux_1087_i24_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i24_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_787_Select_220_i3_4_lut (.I0(n66381), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n66416), .I3(n61341), .O(n3_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51197_2_lut_3_lut (.I0(n3474), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n66982));
    defparam i51197_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
           .D(n30002));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
           .D(n30007));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n30012));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i23_3_lut_4_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1][6] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i23_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_787_Select_219_i3_4_lut (.I0(n69031), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[25] [2]), .I3(\data_out_frame[25] [1]), 
            .O(n3_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_219_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30095));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i22_3_lut_4_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i22_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i21_3_lut_4_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i21_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i59076_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74523));   // verilog/coms.v(158[12:15])
    defparam i59076_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1087_i20_3_lut_4_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i20_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i19_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i19_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i18_3_lut_4_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i18_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_787_Select_218_i3_4_lut (.I0(n66339), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n66710), .I3(\data_out_frame[25] [1]), .O(n3_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i58903_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74509));   // verilog/coms.v(158[12:15])
    defparam i58903_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1087_i16_3_lut_4_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i16_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i15_3_lut_4_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2][6] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i15_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [0]), 
            .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1087_i14_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2]_c [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i14_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i13_3_lut_4_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2][4] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i13_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_787_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i12_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2][3] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i12_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i11_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2]_c [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i11_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_787_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1082 (.I0(n66348), .I1(n66716), .I2(n60565), 
            .I3(GND_net), .O(n60670));
    defparam i2_3_lut_adj_1082.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut (.I0(n60666), .I1(n66772), .I2(\data_out_frame[23] [1]), 
            .I3(n66474), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1083 (.I0(n66413), .I1(\data_out_frame[21] [1]), 
            .I2(n26201), .I3(n66518), .O(n19));
    defparam i7_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
           .D(n30015));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n30093), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n30092), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1084 (.I0(n60585), .I1(\data_out_frame[23] [2]), 
            .I2(n26659), .I3(n60698), .O(n21));
    defparam i9_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19), .I2(n20), .I3(GND_net), .O(n61341));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1087_i10_3_lut_4_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2][1] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i10_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\data_out_frame[21] [0]), .I1(n25417), 
            .I2(GND_net), .I3(GND_net), .O(n66348));
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1086 (.I0(\data_out_frame[20] [7]), .I1(n66348), 
            .I2(n61545), .I3(n66413), .O(n16));
    defparam i6_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i9_3_lut_4_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2][0] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i9_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i7_4_lut_adj_1087 (.I0(n66518), .I1(n61568), .I2(\data_out_frame[16] [4]), 
            .I3(n61315), .O(n17_c));
    defparam i7_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1088 (.I0(n17_c), .I1(n60677), .I2(n16), .I3(n26605), 
            .O(n66416));
    defparam i9_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1089 (.I0(n66797), .I1(n66745), .I2(n66572), 
            .I3(n66845), .O(n10_adj_5377));
    defparam i4_4_lut_adj_1089.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1087_i8_3_lut_4_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[7]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i8_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(n61315), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66710));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1087_i7_3_lut_4_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i7_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[20] [5]), .I1(n66552), .I2(n66416), 
            .I3(n69046), .O(n12_adj_5378));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n30091), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1091 (.I0(\data_out_frame[22] [6]), .I1(n12_adj_5378), 
            .I2(n66710), .I3(\data_out_frame[24] [7]), .O(n69031));
    defparam i6_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i6_3_lut_4_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i6_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i5_3_lut_4_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i5_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[23] [5]), .I1(n68518), 
            .I2(n61070), .I3(n26526), .O(n66707));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1087_i4_3_lut_4_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i4_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i3_3_lut_4_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i3_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1087_i2_3_lut_4_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i2_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(n26526), .I1(n66444), .I2(GND_net), 
            .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n82), .I2(reset), 
            .I3(n3474), .O(n66099));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n30090), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_217_i3_4_lut (.I0(n5), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n66546), .I3(n69031), .O(n3_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n30089), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1093 (.I0(\data_out_frame[24] [6]), .I1(n61587), 
            .I2(\data_out_frame[25] [0]), .I3(n66515), .O(n66339));
    defparam i3_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n30088), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n30087), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_216_i3_3_lut (.I0(n66339), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n66707), .I3(GND_net), .O(n3_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n30086), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n30085), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1094 (.I0(\data_out_frame[20] [2]), .I1(n61643), 
            .I2(\data_out_frame[20] [3]), .I3(n61306), .O(n61603));
    defparam i1_2_lut_3_lut_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_4_lut_adj_1095 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n3474), .O(n66108));   // verilog/coms.v(157[7:23])
    defparam i2_3_lut_4_lut_4_lut_adj_1095.LUT_INIT = 16'hfbff;
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n30084), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_1745_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n30083), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n30082), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n30081), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n30080), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1096 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5381), .I3(n66131), .O(n27316));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'haaa8;
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n30079), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n30078), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i55925_4_lut (.I0(\data_out_frame[0][4] ), .I1(\data_out_frame[3][4] ), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n71760));
    defparam i55925_4_lut.LUT_INIT = 16'hc00a;
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n30077), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n30076), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n30075), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66381));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i59078_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74524));   // verilog/coms.v(158[12:15])
    defparam i59078_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n30074), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n30073), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n30072), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n30071), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5383));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55928_4_lut (.I0(n1_adj_5383), .I1(\data_out_frame[3][3] ), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n71763));
    defparam i55928_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i55994_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71829));
    defparam i55994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55995_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71830));
    defparam i55995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1098 (.I0(n66672), .I1(n66381), .I2(\data_out_frame[25] [1]), 
            .I3(n66824), .O(n10_adj_5384));
    defparam i4_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n30070), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n30069), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n30068), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56064_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71899));
    defparam i56064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56063_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71898));
    defparam i56063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1087_i1_3_lut_4_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n4930[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i1_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i55991_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71826));
    defparam i55991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55992_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71827));
    defparam i55992_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n30067), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n30066), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n30065), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(n25877), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_5385));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i56001_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71836));
    defparam i56001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56000_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71835));
    defparam i56000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56012_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71847));
    defparam i56012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56013_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71848));
    defparam i56013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56022_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71857));
    defparam i56022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56021_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71856));
    defparam i56021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56039_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71874));
    defparam i56039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56040_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71875));
    defparam i56040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55941_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71776));
    defparam i55941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55940_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71775));
    defparam i55940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1099 (.I0(\data_in_frame[18] [3]), .I1(n60757), 
            .I2(\data_in_frame[20] [5]), .I3(\data_in_frame[22] [7]), .O(n70933));
    defparam i1_3_lut_4_lut_adj_1099.LUT_INIT = 16'h9669;
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n30064), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n30063), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n30062), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56078_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71913));
    defparam i56078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_215_i3_4_lut (.I0(n66333), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n66707), .I3(\data_out_frame[25] [0]), .O(n3_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_215_i3_4_lut.LUT_INIT = 16'h8448;
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n30061), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56079_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71914));
    defparam i56079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59079_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74525));   // verilog/coms.v(158[12:15])
    defparam i59079_2_lut.LUT_INIT = 16'h2222;
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n30060), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i56082_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71917));
    defparam i56082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56081_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71916));
    defparam i56081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1100 (.I0(reset), .I1(n10_adj_5387), 
            .I2(n3474), .I3(n161), .O(n66156));
    defparam i1_2_lut_3_lut_4_lut_adj_1100.LUT_INIT = 16'hefff;
    SB_LUT4 i56033_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71868));
    defparam i56033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56034_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71869));
    defparam i56034_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n30059), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n30058), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n30057), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n30056), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n30055), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n30054), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2), .S(n65962));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2872), .D(n6_adj_5388), .S(n65961));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5389), .S(n65960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n30053), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5390), .S(n65959));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5391), .S(n65958));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n30052), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5392), .S(n65957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5393), .S(n65956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n30051), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i55968_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71803));
    defparam i55968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55967_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71802));
    defparam i55967_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n30050), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n30049), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n30048), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n30047), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n65839));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1101 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n65841));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1101.LUT_INIT = 16'h5100;
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5364), .S(n65955));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1102 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n65842));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1102.LUT_INIT = 16'h5100;
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n30046), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1103 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n65843));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1103.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1104 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n65844));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1104.LUT_INIT = 16'h5100;
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n30045), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n30044), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n30043), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n30042), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5361), .S(n65954));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5360), .S(n65953));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5359), .S(n65952));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5358), .S(n65951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5357), .S(n65950));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n30041), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1105 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n65837));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1105.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1106 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n65845));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1106.LUT_INIT = 16'h5100;
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n30040), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n30039), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1107 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n65836));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1107.LUT_INIT = 16'h5100;
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2872), .D(n7_adj_5356), .S(n65949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5355), .S(n65948));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1108 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n65840));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1108.LUT_INIT = 16'h5100;
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n30038), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1109 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n65846));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1109.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1110 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n65847));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1110.LUT_INIT = 16'h5100;
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n30037), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n30036), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1111 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n65848));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1111.LUT_INIT = 16'h5100;
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5394), .S(n65947));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1112 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n65849));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1112.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1113 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n65838));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1113.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(n66276), .I3(GND_net), .O(Kp_23__N_767));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5395), .S(n65946));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5396), .S(n65945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n30035), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1114 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n65850));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1114.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1115 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n65851));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1115.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1116 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(n61751), .I3(\data_out_frame[17] [2]), .O(n6_adj_5397));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1117 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(n61751), .I3(n27157), .O(n66594));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n30034), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n30033), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n30032), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1118 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n70901));
    defparam i1_2_lut_3_lut_adj_1118.LUT_INIT = 16'h9696;
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n30031), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n30030), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5398), .S(n65944));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5399), .S(n65853));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n65378));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1119 (.I0(n28670), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n65432));
    defparam i1_4_lut_4_lut_4_lut_adj_1119.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1120 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n66216));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1120.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5400), .S(n65943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5401), .S(n65856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n30029), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n30028), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1121 (.I0(n28670), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n65434));
    defparam i1_4_lut_4_lut_4_lut_adj_1121.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1122 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[4] [3]), .O(n66264));   // verilog/coms.v(76[16:42])
    defparam i1_3_lut_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3] [6]), .I3(GND_net), .O(n6_adj_5402));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5403), .S(n65942));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(n66689), .I3(Kp_23__N_772), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1124 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[0][0] ), 
            .I2(\data_in_frame[2][1] ), .I3(\data_in_frame[3] [7]), .O(n66689));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n30027), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i30396_2_lut (.I0(LED_c), .I1(LED_N_3408), .I2(GND_net), .I3(GND_net), 
            .O(LED_N_3407));   // verilog/coms.v(253[15] 255[9])
    defparam i30396_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14997_4_lut (.I0(n2872), .I1(LED_N_3407), .I2(n27768), .I3(\FRAME_MATCHER.i_31__N_2513 ), 
            .O(n29209));   // verilog/coms.v(130[12] 305[6])
    defparam i14997_4_lut.LUT_INIT = 16'ha8a0;
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n30026), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5404), .S(n65861));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_1743_Select_0_i3_3_lut (.I0(LED_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n3_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_1743_Select_0_i3_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1125 (.I0(LED_c), .I1(n3_adj_5405), .I2(Kp_23__N_1748), 
            .I3(Kp_23__N_612), .O(n5_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1125.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[24] [5]), .I1(n24043), 
            .I2(GND_net), .I3(GND_net), .O(n66333));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[9] [7]), .I1(n24272), .I2(n27046), 
            .I3(n66763), .O(n66719));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5407), .S(n65865));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5408), .S(n65866));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(n24272), .I1(n27046), .I2(n66763), 
            .I3(GND_net), .O(n66352));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n30025), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n30024), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n30023), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5409), .S(n65867));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n30022), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5410), .S(n65868));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5411), .S(n65869));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5412), .S(n65872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n30021), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5413), .S(n65875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5414), .S(n29286));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5415), .S(n65876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5416), .S(n65877));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n30020), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n30019), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n30018), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5417), .S(n65878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5418), .S(n65879));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[24] [4]), .I1(n25456), 
            .I2(GND_net), .I3(GND_net), .O(n66549));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5419), .S(n65880));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5420), .S(n65874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5421), .S(n65881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5422), .S(n65882));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5423), .S(n65883));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1129 (.I0(n26873), .I1(n61123), .I2(\data_in_frame[12] [4]), 
            .I3(n26416), .O(n61589));
    defparam i2_3_lut_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5424), .S(n65884));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16420_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30632));   // verilog/coms.v(130[12] 305[6])
    defparam i16420_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15737_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29949));   // verilog/coms.v(130[12] 305[6])
    defparam i15737_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n30005));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n30001));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1130 (.I0(n26424), .I1(\data_in_frame[12] [5]), 
            .I2(n26873), .I3(GND_net), .O(n26416));
    defparam i1_2_lut_3_lut_adj_1130.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1131 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'ha088;
    SB_LUT4 i16450_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30662));   // verilog/coms.v(130[12] 305[6])
    defparam i16450_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n76856), .I2(n74616), .I3(byte_transmit_counter[4]), .O(n79011));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n79011_bdd_4_lut (.I0(n79011), .I1(n78618), .I2(n7_adj_7), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n79011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1132 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(\data_in_frame[10] [3]), .I3(GND_net), .O(n71295));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1132.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n30000));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29999));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29998));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29997));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29996));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_213_i3_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n66549), .I3(n68582), .O(n3_adj_5426));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_213_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i16449_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30661));   // verilog/coms.v(130[12] 305[6])
    defparam i16449_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29995));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16448_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30660));   // verilog/coms.v(130[12] 305[6])
    defparam i16448_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29994));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1133 (.I0(n68633), .I1(n66863), .I2(\data_in_frame[17] [7]), 
            .I3(\data_in_frame[17] [6]), .O(n66584));
    defparam i2_3_lut_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1134 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [2]), 
            .I2(n66698), .I3(n26685), .O(n26957));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1135 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n66698));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i16447_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30659));   // verilog/coms.v(130[12] 305[6])
    defparam i16447_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29993));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16446_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30658));   // verilog/coms.v(130[12] 305[6])
    defparam i16446_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16445_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30657));   // verilog/coms.v(130[12] 305[6])
    defparam i16445_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16444_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30656));   // verilog/coms.v(130[12] 305[6])
    defparam i16444_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1136 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [4]), 
            .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n6_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1136.LUT_INIT = 16'ha088;
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29992));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29991));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29990));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16443_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30655));   // verilog/coms.v(130[12] 305[6])
    defparam i16443_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut (.I0(n24039), .I1(\data_out_frame[24] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5427));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63083 (.I0(byte_transmit_counter[3]), 
            .I1(n76854), .I2(n74617), .I3(byte_transmit_counter[4]), .O(n79005));
    defparam byte_transmit_counter_3__bdd_4_lut_63083.LUT_INIT = 16'he4aa;
    SB_LUT4 i16441_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30653));   // verilog/coms.v(130[12] 305[6])
    defparam i16441_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_211_i3_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5427), .I3(n61765), 
            .O(n3_adj_5428));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i16440_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30652));   // verilog/coms.v(130[12] 305[6])
    defparam i16440_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16439_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30651));   // verilog/coms.v(130[12] 305[6])
    defparam i16439_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29988));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29987));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode_c[2]), .C(clk16MHz), .D(n53030));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode_c[3]), .C(clk16MHz), .D(n29985));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode_c[4]), .C(clk16MHz), .D(n29983));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(\control_mode[5] ), .C(clk16MHz), .D(n29982));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk16MHz), .D(n29981));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(\control_mode[7] ), .C(clk16MHz), .D(n29977));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(\current_limit[1] ), .C(clk16MHz), .D(n29974));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(\current_limit[2] ), .C(clk16MHz), .D(n29973));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(\current_limit[3] ), .C(clk16MHz), .D(n29972));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(\current_limit[4] ), .C(clk16MHz), .D(n29971));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(\current_limit[5] ), .C(clk16MHz), .D(n29970));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29942), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(\current_limit[0] ), .C(clk16MHz), .D(n29941));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(\control_mode[0] ), .C(clk16MHz), .D(n29940));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29938), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29937), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29936), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29933), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1137 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(n66312), .I3(n66695), .O(n71181));
    defparam i1_3_lut_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1138 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [0]), 
            .I2(\data_out_frame[24] [1]), .I3(n66739), .O(n10_adj_5429));
    defparam i4_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5430), .S(n65885));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_210_i3_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n10_adj_5429), .I3(n68518), 
            .O(n3_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_210_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i16438_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30650));   // verilog/coms.v(130[12] 305[6])
    defparam i16438_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5432), .S(n65886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5433), .S(n65887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5434), .S(n65888));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5435), .S(n65889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5436), .S(n65890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5437), .S(n65891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5438), .S(n65892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5439), .S(n65893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5440), .S(n65894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5441), .S(n65895));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5442), .S(n65896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5443), .S(n65897));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5444), .S(n65898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5445), .S(n65899));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5446), .S(n65900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5447), .S(n65901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5448), .S(n65902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5449), .S(n65903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5450), .S(n65904));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5451), .S(n65905));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5452), .S(n65906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5453), .S(n65907));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5454), .S(n65908));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5455), .S(n65909));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16437_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30649));   // verilog/coms.v(130[12] 305[6])
    defparam i16437_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n79005_bdd_4_lut (.I0(n79005), .I1(n78594), .I2(n7_adj_8), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n79005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16436_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30648));   // verilog/coms.v(130[12] 305[6])
    defparam i16436_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1139 (.I0(n26244), .I1(n26329), .I2(n26685), 
            .I3(n26846), .O(n66860));
    defparam i1_2_lut_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i20958_3_lut_4_lut (.I0(\Kp[10] ), .I1(\data_in_frame[2]_c [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30038));
    defparam i20958_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i14487_4_lut (.I0(n10_adj_5387), .I1(reset), .I2(n66982), 
            .I3(n8_adj_9), .O(n7));
    defparam i14487_4_lut.LUT_INIT = 16'hffef;
    SB_DFFR \FRAME_MATCHER.i_2043__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n28323), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i16435_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30647));   // verilog/coms.v(130[12] 305[6])
    defparam i16435_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1140 (.I0(n60664), .I1(n70901), .I2(n66666), 
            .I3(GND_net), .O(n66827));
    defparam i1_2_lut_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1141 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [5]), 
            .I2(n26343), .I3(n26362), .O(n66212));
    defparam i1_2_lut_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2043__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n28325), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n28327), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n28329), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n28331), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n28335), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n28337), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n28339), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n28341), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n28343), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n28345), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28347), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28349), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28351), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28353), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28355), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28357), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28359), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28361), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28363), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28365), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28367), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28369), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28371), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28373), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28375), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28377), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n28379), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n28381), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n28383), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28385), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28387), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5458), .S(n65910));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5459), .S(n29249));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5460), .S(n65911));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1142 (.I0(\data_in_frame[13] [5]), .I1(n26343), 
            .I2(n26362), .I3(GND_net), .O(n26378));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5461), .S(n65912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5462), .S(n65913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5463), .S(n65914));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16434_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30646));   // verilog/coms.v(130[12] 305[6])
    defparam i16434_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63078 (.I0(byte_transmit_counter[3]), 
            .I1(n76848), .I2(n74635), .I3(byte_transmit_counter[4]), .O(n78987));
    defparam byte_transmit_counter_3__bdd_4_lut_63078.LUT_INIT = 16'he4aa;
    SB_LUT4 n78987_bdd_4_lut (.I0(n78987), .I1(n78624), .I2(n7_adj_10), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n78987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63063 (.I0(byte_transmit_counter[3]), 
            .I1(n76846), .I2(n74611), .I3(byte_transmit_counter[4]), .O(n78975));
    defparam byte_transmit_counter_3__bdd_4_lut_63063.LUT_INIT = 16'he4aa;
    SB_LUT4 n78975_bdd_4_lut (.I0(n78975), .I1(n78606), .I2(n7_adj_11), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n78975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5466), .S(n65873));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5467), .S(n66039));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5468), .S(n66038));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1143 (.I0(n7_adj_5469), .I1(n68344), .I2(n69046), 
            .I3(n26743), .O(n26827));
    defparam i4_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1144 (.I0(n68553), .I1(n66447), .I2(n26827), 
            .I3(n61306), .O(n12_adj_5470));
    defparam i5_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i16433_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30645));   // verilog/coms.v(130[12] 305[6])
    defparam i16433_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1145 (.I0(\data_out_frame[22] [1]), .I1(n12_adj_5470), 
            .I2(n66745), .I3(n61643), .O(n61765));
    defparam i6_4_lut_adj_1145.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1146 (.I0(n26827), .I1(n66391), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n68582));
    defparam i2_3_lut_adj_1146.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1147 (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n66574));
    defparam i1_2_lut_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66378));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i16432_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30644));   // verilog/coms.v(130[12] 305[6])
    defparam i16432_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26605));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i20933_3_lut_4_lut (.I0(\Kp[13] ), .I1(\data_in_frame[2]_c [5]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30035));
    defparam i20933_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_adj_1150 (.I0(n26343), .I1(n26957), .I2(n66734), 
            .I3(GND_net), .O(n12_adj_5471));
    defparam i1_2_lut_3_lut_adj_1150.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n66716));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i16431_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30643));   // verilog/coms.v(130[12] 305[6])
    defparam i16431_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26201));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(\data_out_frame[19] [3]), .I1(n60778), 
            .I2(GND_net), .I3(GND_net), .O(n14_c));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5472), .S(n66037));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5473), .S(n66036));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(\current_limit[8] ), .C(clk16MHz), .D(n30784));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16430_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30642));   // verilog/coms.v(130[12] 305[6])
    defparam i16430_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1154 (.I0(\data_out_frame[17] [3]), .I1(n61533), 
            .I2(n66748), .I3(\data_out_frame[17] [7]), .O(n22_adj_5474));
    defparam i9_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1155 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [6]), 
            .I2(n66450), .I3(\data_out_frame[16] [5]), .O(n21_adj_5475));
    defparam i8_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i10_4_lut_adj_1156 (.I0(n60763), .I1(n26201), .I2(\data_out_frame[17] [4]), 
            .I3(n14_c), .O(n23_adj_5476));
    defparam i10_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i16429_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30641));   // verilog/coms.v(130[12] 305[6])
    defparam i16429_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1157 (.I0(n23_adj_5476), .I1(n66166), .I2(n21_adj_5475), 
            .I3(n22_adj_5474), .O(n16_adj_5477));
    defparam i3_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i16428_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30640));   // verilog/coms.v(130[12] 305[6])
    defparam i16428_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1158 (.I0(n61533), .I1(n66491), .I2(\data_out_frame[19] [4]), 
            .I3(n60624), .O(n22_adj_5478));
    defparam i9_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16427_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30639));   // verilog/coms.v(130[12] 305[6])
    defparam i16427_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16426_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30638));   // verilog/coms.v(130[12] 305[6])
    defparam i16426_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16425_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30637));   // verilog/coms.v(130[12] 305[6])
    defparam i16425_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16424_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30636));   // verilog/coms.v(130[12] 305[6])
    defparam i16424_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16423_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30635));   // verilog/coms.v(130[12] 305[6])
    defparam i16423_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_4_lut (.I0(n60581), .I1(n22_adj_5478), .I2(n16_adj_5477), 
            .I3(\data_out_frame[18] [7]), .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16422_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30634));   // verilog/coms.v(130[12] 305[6])
    defparam i16422_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16421_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30633));   // verilog/coms.v(130[12] 305[6])
    defparam i16421_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16442_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30654));   // verilog/coms.v(130[12] 305[6])
    defparam i16442_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12_4_lut_adj_1159 (.I0(\data_out_frame[14] [3]), .I1(n24), 
            .I2(n20_adj_5479), .I3(\data_out_frame[18] [2]), .O(n66772));
    defparam i12_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(n60607), .I1(n66312), .I2(\data_in_frame[12] [1]), 
            .I3(GND_net), .O(n66692));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(n27157), .I1(n66772), .I2(GND_net), 
            .I3(GND_net), .O(n66845));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1161 (.I0(n69038), .I1(n10_adj_5480), .I2(\data_in_frame[15] [5]), 
            .I3(\data_in_frame[18] [1]), .O(n66497));
    defparam i1_2_lut_4_lut_adj_1161.LUT_INIT = 16'h9669;
    SB_DFF current_limit_i0_i9 (.Q(\current_limit[9] ), .C(clk16MHz), .D(n30783));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(\current_limit[10] ), .C(clk16MHz), 
           .D(n30779));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1162 (.I0(n66587), .I1(n66531), .I2(n60780), 
            .I3(n66845), .O(n10_adj_5481));
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n37697));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n30777));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n30776));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n30775));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n65176));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n30773));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n30772), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30771), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30770), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30768), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n65172));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30766), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30764), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n30761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n65168));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n65164));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29729));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29732));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n65160));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
           .D(n29738));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30735), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30734), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29741));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n30732));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30731), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30730), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n29744));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30728), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30725));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
           .D(n29747));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30723), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
           .D(n29750));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30721), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30720), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(n66571), .I1(n10_adj_5481), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n61545));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30697), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30679), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
           .D(n29754));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30677), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n30676));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1163 (.I0(n28674), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[10]_c [2]), .O(n65364));
    defparam i1_4_lut_4_lut_4_lut_adj_1163.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n30664));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30663), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30662));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30661));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30660));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30659));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30658));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30657));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30656));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30654));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30653));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30652));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30651));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30650));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30649));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30648));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30647));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30646));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30645));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30644));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30643));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30642));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30641));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30640));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30639));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5370), .S(n66035));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30637));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30634));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30633));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30631), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n30630));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30629), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30628), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n30247));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n29757));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n30250));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30624), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n30253));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30622), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
           .D(n29761));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n30256));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n30259));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n30262));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n30617));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5366), .S(n66034));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20][0] ), .C(clk16MHz), 
           .D(n29764));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20][1] ), .C(clk16MHz), 
           .D(n29767));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20][2] ), .C(clk16MHz), 
           .D(n29770));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0][1] ), .C(clk16MHz), 
           .D(n65360));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20][3] ), .C(clk16MHz), 
           .D(n29777));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20][4] ), .C(clk16MHz), 
           .D(n29780));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n65218));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29786));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n65224));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29792));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29795));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30265));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n30601));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29798));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29801));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10][0] ), .C(clk16MHz), 
           .D(n30268));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10]_c [1]), .C(clk16MHz), 
           .D(n30271));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10]_c [2]), .C(clk16MHz), 
           .D(n65364));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
           .D(n30278));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10]_c [4]), .C(clk16MHz), 
           .D(n65368));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10][5] ), .C(clk16MHz), 
           .D(n30284));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10][6] ), .C(clk16MHz), 
           .D(n30288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30591));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29804));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n30587));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n30586));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29807));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10][7] ), .C(clk16MHz), 
           .D(n30291));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n30583));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29810));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29813));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n30294));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n30298));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n65336));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n30304));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n30308));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n65318));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30314));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30318));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30321));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29816));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30324));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n65378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n65432));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n65434));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n30337));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n30340));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30344));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30347));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30350));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30353));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30357));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13]_c [4]), .C(clk16MHz), 
           .D(n30360));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30363));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13][6] ), .C(clk16MHz), 
           .D(n30366));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13][7] ), .C(clk16MHz), 
           .D(n30370));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n30373));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5315), .S(n65863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5314), .S(n65860));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n30376));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
           .D(n30380));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i116 (.Q(\data_in_frame[14]_c [3]), .C(clk16MHz), 
           .D(n30383));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14][4] ), .C(clk16MHz), 
           .D(n30386));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14][5] ), .C(clk16MHz), 
           .D(n30390));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14][6] ), .C(clk16MHz), 
           .D(n30393));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14][7] ), .C(clk16MHz), 
           .D(n30396));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
           .D(n30400));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
           .D(n30403));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
           .D(n30406));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
           .D(n30410));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
           .D(n15));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n30416));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
           .D(n30420));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
           .D(n30423));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
           .D(n65154));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
           .D(n30430));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
           .D(n65150));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n65146));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n65094));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n30443));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n30446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
           .D(n65142));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n65244));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n30456));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n65276));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n65272));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n65268));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n30515));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5311), .S(n66033));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29819));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29822));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29825));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29828));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29831));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29834));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29837));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29840));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29843));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n65400));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0][3] ), .C(clk16MHz), 
           .D(n29849));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n65402));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n65134));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29858));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29861));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n65132));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n65130));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29870));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0][5] ), .C(clk16MHz), 
           .D(n29874));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0][6] ), .C(clk16MHz), 
           .D(n29877));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0][7] ), .C(clk16MHz), 
           .D(n65398));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1164 (.I0(\data_in_frame[9] [3]), .I1(n60664), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n61555));
    defparam i1_2_lut_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i9 (.Q(\data_in_frame[1][0] ), .C(clk16MHz), 
           .D(n29883));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
           .D(n29886));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i58846_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74409));   // verilog/coms.v(158[12:15])
    defparam i58846_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
           .D(n29889));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
           .D(n29892));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_out_frame[18] [3]), .I1(n60269), 
            .I2(GND_net), .I3(GND_net), .O(n60677));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_out_frame[16] [3]), .I1(n61645), 
            .I2(GND_net), .I3(GND_net), .O(n61568));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
           .D(n29895));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
           .D(n29898));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i59199_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74410));   // verilog/coms.v(158[12:15])
    defparam i59199_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i15 (.Q(\data_in_frame[1][6] ), .C(clk16MHz), 
           .D(n29901));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i58847_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74411));   // verilog/coms.v(158[12:15])
    defparam i58847_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i58946_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74414));   // verilog/coms.v(158[12:15])
    defparam i58946_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
           .D(n29905));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i17 (.Q(\data_in_frame[2][0] ), .C(clk16MHz), 
           .D(n29909));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1167 (.I0(\data_out_frame[18] [2]), .I1(n66231), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5482));
    defparam i2_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i18 (.Q(\data_in_frame[2][1] ), .C(clk16MHz), 
           .D(n29914));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1168 (.I0(n7_adj_5482), .I1(\data_out_frame[18] [1]), 
            .I2(n61607), .I3(n66604), .O(n61306));
    defparam i4_4_lut_adj_1168.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i19 (.Q(\data_in_frame[2]_c [2]), .C(clk16MHz), 
           .D(n29917));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i20 (.Q(\data_in_frame[2][3] ), .C(clk16MHz), 
           .D(n29920));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66528));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1170 (.I0(n28674), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[10]_c [4]), .O(n65368));
    defparam i1_4_lut_4_lut_4_lut_adj_1170.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i21 (.Q(\data_in_frame[2][4] ), .C(clk16MHz), 
           .D(n29923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5308), .S(n66032));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5483), .S(n66031));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5484), .S(n65870));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5485), .S(n65864));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5486), .S(n66030));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1171 (.I0(\data_out_frame[17] [6]), .I1(n66604), 
            .I2(n66453), .I3(n1720), .O(n68559));
    defparam i3_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1172 (.I0(n68131), .I1(n26537), .I2(n61678), 
            .I3(GND_net), .O(n66488));
    defparam i1_2_lut_3_lut_adj_1172.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF data_in_frame_0___i22 (.Q(\data_in_frame[2]_c [5]), .C(clk16MHz), 
           .D(n29926));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i23 (.Q(\data_in_frame[2][6] ), .C(clk16MHz), 
           .D(n29929));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i58853_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74415));   // verilog/coms.v(158[12:15])
    defparam i58853_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5487), .S(n66029));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5488), .S(n66028));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i58947_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74417));   // verilog/coms.v(158[12:15])
    defparam i58947_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_adj_1173 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\data_out_frame[0][2] ), .I3(GND_net), .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_adj_1173.LUT_INIT = 16'ha8a8;
    SB_LUT4 i5_4_lut_adj_1174 (.I0(n68559), .I1(\data_out_frame[15] [7]), 
            .I2(n66794), .I3(n66608), .O(n12_adj_5489));
    defparam i5_4_lut_adj_1174.LUT_INIT = 16'h9669;
    SB_LUT4 i55953_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71788));
    defparam i55953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1175 (.I0(n61533), .I1(n12_adj_5489), .I2(n66166), 
            .I3(n66528), .O(n61643));
    defparam i6_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i55954_4_lut (.I0(n71788), .I1(n28441), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][5] ), .O(n71789));
    defparam i55954_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i55952_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71787));
    defparam i55952_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n28129), 
            .D(n4930[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1176 (.I0(n68633), .I1(\data_in_frame[15] [5]), 
            .I2(n24165), .I3(GND_net), .O(n61678));
    defparam i1_2_lut_3_lut_adj_1176.LUT_INIT = 16'h6969;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n28129), 
            .D(n4930[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n28129), 
            .D(n4930[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n28129), 
            .D(n4930[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n28129), 
            .D(n4930[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n28129), 
            .D(n4930[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n28129), 
            .D(n4930[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n28129), 
            .D(n4938), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n28129), 
            .D(n4930[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n28129), 
            .D(n4930[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n28129), 
            .D(n4930[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n28129), 
            .D(n4930[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n28129), 
            .D(n4930[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n28129), 
            .D(n4930[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n28129), 
            .D(n4930[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n28129), 
            .D(n4930[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n28129), 
            .D(n4930[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n28129), 
            .D(n4930[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n28129), 
            .D(n4930[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n28129), 
            .D(n4930[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n28129), 
            .D(n4930[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n28129), 
            .D(n4930[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n28129), 
            .D(n4930[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n79076), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i1_2_lut_4_lut_adj_1177 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[13][7] ), 
            .I2(\data_in_frame[13][6] ), .I3(n61308), .O(n66524));
    defparam i1_2_lut_4_lut_adj_1177.LUT_INIT = 16'h9669;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n27427), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2046), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2047), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20637), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n65018), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2058), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27430), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i1_3_lut_4_lut_adj_1178 (.I0(\data_in_frame[14][7] ), .I1(n26362), 
            .I2(n26870), .I3(n61658), .O(n66776));
    defparam i1_3_lut_4_lut_adj_1178.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5490), .S(n66027));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[20] [3]), .I1(n61306), 
            .I2(GND_net), .I3(GND_net), .O(n61605));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59117_2_lut (.I0(n78798), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74611));
    defparam i59117_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5491), .S(n66026));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5492), .S(n66025));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5493), .S(n66024));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1180 (.I0(\data_in_frame[16] [6]), .I1(n60656), 
            .I2(n26758), .I3(GND_net), .O(n66495));
    defparam i1_2_lut_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i61011_3_lut (.I0(n78756), .I1(n78648), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76846));
    defparam i61011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1181 (.I0(\data_in_frame[9] [3]), .I1(n66568), 
            .I2(n71177), .I3(\data_in_frame[12] [1]), .O(n6_adj_5494));
    defparam i1_2_lut_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1182 (.I0(\data_in_frame[14][6] ), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[17] [2]), .O(n71059));
    defparam i1_3_lut_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5495), .S(n66023));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5496), .S(n66022));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5497), .S(n66021));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5498), .S(n66020));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5499), .S(n66019));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5500), .S(n66018));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5501), .S(n65974));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5502), .S(n66017));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5503), .S(n66016));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5504), .S(n66015));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5505), .S(n66014));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5506), .S(n66013));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1183 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [0]), 
            .I2(encoder1_position[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1183.LUT_INIT = 16'ha088;
    SB_LUT4 i4_4_lut_adj_1184 (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[20] [0]), 
            .I2(\data_out_frame[17] [6]), .I3(n61240), .O(n10_adj_5507));
    defparam i4_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i30012_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n44101));   // verilog/coms.v(105[12:33])
    defparam i30012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1185 (.I0(\data_in_frame[20] [7]), .I1(n66495), 
            .I2(n68457), .I3(\data_in_frame[18] [6]), .O(n66683));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i55950_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71785));
    defparam i55950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1186 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0][5] ), 
            .I2(\data_in_frame[1][0] ), .I3(Kp_23__N_767), .O(n26583));
    defparam i1_2_lut_3_lut_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1187 (.I0(n68646), .I1(\data_in_frame[14] [2]), 
            .I2(n61528), .I3(GND_net), .O(n25588));
    defparam i1_2_lut_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i55951_4_lut (.I0(n71785), .I1(n44101), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n71786));
    defparam i55951_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i55949_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71784));
    defparam i55949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1188 (.I0(\data_in_frame[13] [0]), .I1(n26424), 
            .I2(\data_in_frame[12] [5]), .I3(n26873), .O(n26870));
    defparam i1_2_lut_3_lut_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1189 (.I0(n26758), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n66407));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1189.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1190 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n60640), .I3(GND_net), .O(n60698));
    defparam i2_3_lut_adj_1190.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1191 (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(n66108), .I3(n10_adj_5508), .O(n28670));
    defparam i1_2_lut_3_lut_4_lut_adj_1191.LUT_INIT = 16'hfffd;
    SB_LUT4 select_787_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1192 (.I0(n60658), .I1(n60269), .I2(\data_out_frame[18] [3]), 
            .I3(\data_out_frame[18] [4]), .O(n69046));
    defparam i2_3_lut_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i58949_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74421));   // verilog/coms.v(158[12:15])
    defparam i58949_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5509), .S(n66012));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5510), .S(n66011));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1193 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[4] [5]), .I3(n66666), .O(Kp_23__N_993));
    defparam i1_2_lut_3_lut_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1194 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1194.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1195 (.I0(\data_in_frame[0][3] ), .I1(\data_in_frame[2][4] ), 
            .I2(\data_in_frame[0] [2]), .I3(n26722), .O(Kp_23__N_799));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5511), .S(n66010));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1196 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1196.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(\data_out_frame[16] [1]), .I1(n60698), 
            .I2(GND_net), .I3(GND_net), .O(n61607));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59268_2_lut (.I0(n78852), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n74635));
    defparam i59268_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5512), .S(n65915));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1198 (.I0(n1835), .I1(n26941), .I2(n60677), .I3(n66528), 
            .O(n10_adj_5513));
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5514), .S(n65916));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i61013_3_lut (.I0(n78726), .I1(n78564), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76848));
    defparam i61013_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF current_limit_i0_i6 (.Q(\current_limit[6] ), .C(clk16MHz), .D(n29753));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5515), .S(n65917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5516), .S(n65918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5517), .S(n65919));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5518), .S(n65920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5519), .S(n65921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5520), .S(n65922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5521), .S(n65923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5522), .S(n65924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5523), .S(n65925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5524), .S(n65926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5525), .S(n65927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5526), .S(n65928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5527), .S(n65929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5528), .S(n66009));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_3_lut (.I0(LED_N_3408), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(reset), .I3(GND_net), .O(n23023));   // verilog/coms.v(130[12] 305[6])
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1199 (.I0(\data_in_frame[16] [3]), .I1(n68646), 
            .I2(n61749), .I3(\data_in_frame[18] [4]), .O(n71157));
    defparam i1_2_lut_3_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5529), .S(n65862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5530), .S(n66008));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5531), .S(n65859));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5532), .S(n65930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5533), .S(n65931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5534), .S(n65932));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5535), .S(n65933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5536), .S(n65934));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5537), .S(n65935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5538), .S(n65936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5539), .S(n65937));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5540), .S(n65938));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5541), .S(n65939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5542), .S(n65857));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5543), .S(n65940));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5544), .S(n65941));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5545), .S(n65839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5546), .S(n65841));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5431), .S(n65842));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5428), .S(n65843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5547), .S(n65844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5426), .S(n65837));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5548), .S(n65845));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2872), .D(n5_adj_5406), 
            .S(n29209));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5386), .S(n65836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5382), .S(n66007));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2872), .D(n27316), 
            .S(n29199));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2872), .D(n1), .S(n29193));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5380), .S(n65840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5379), .S(n65846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5376), .S(n65847));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5375), .S(n65848));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5374), .S(n65849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5373), .S(n65838));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2872), .D(n3_adj_5372), .S(n65850));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2872), .D(n3), .S(n65851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2872), .D(n1_adj_5549), .S(n65830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2872), .D(n1_adj_5550), .S(n65831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5371), .S(n66006));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(\current_limit[7] ), .C(clk16MHz), .D(n29725));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5368), .S(n66005));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2872), .D(n1_adj_5551), .S(n65827));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1200 (.I0(\data_out_frame[22] [1]), .I1(n60687), 
            .I2(\data_out_frame[21] [7]), .I3(n66435), .O(n10_adj_5552));
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1201 (.I0(n66562), .I1(n10_adj_5552), .I2(n61603), 
            .I3(GND_net), .O(n66391));
    defparam i5_3_lut_adj_1201.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1202 (.I0(\data_out_frame[19] [0]), .I1(n61568), 
            .I2(n60565), .I3(\data_out_frame[20] [7]), .O(n12_adj_5553));
    defparam i5_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2872), .D(n1_adj_5554), .S(n65832));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1203 (.I0(\data_out_frame[21] [1]), .I1(n12_adj_5553), 
            .I2(n66587), .I3(n61543), .O(n26898));
    defparam i6_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2872), .D(n1_adj_5555), .S(n65828));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2872), .D(n1_adj_5556), .S(n65833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2872), .D(n1_adj_5557), .S(n65834));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5363), .S(n66004));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[16] [3]), .I1(n68646), 
            .I2(n61749), .I3(n68457), .O(n60291));
    defparam i1_2_lut_3_lut_4_lut_adj_1204.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5362), .S(n66002));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1205 (.I0(n68518), .I1(n61070), .I2(GND_net), 
            .I3(GND_net), .O(n66616));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h9999;
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2872), .D(n1_adj_5558), .S(n65829));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5354), .S(n65858));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1206 (.I0(n26343), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[13]_c [4]), .I3(n66597), .O(n61601));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_63053 (.I0(byte_transmit_counter[3]), 
            .I1(n76800), .I2(n74610), .I3(byte_transmit_counter[4]), .O(n78921));
    defparam byte_transmit_counter_3__bdd_4_lut_63053.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2872), .D(n2_adj_5349), .S(n66001));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1207 (.I0(\data_out_frame[17] [5]), .I1(n1720), 
            .I2(n66438), .I3(\data_out_frame[15] [4]), .O(n60624));
    defparam i1_4_lut_adj_1207.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1208 (.I0(n60624), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[22] [0]), .I3(n61240), .O(n5_adj_5559));
    defparam i1_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_out_frame[17] [4]), .I1(n66356), 
            .I2(n26087), .I3(n61751), .O(n61240));
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1210 (.I0(n26685), .I1(n26846), .I2(\data_in_frame[9] [2]), 
            .I3(\data_in_frame[14] [1]), .O(n9_adj_5560));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1211 (.I0(\data_out_frame[19] [5]), .I1(n68678), 
            .I2(n61240), .I3(GND_net), .O(n26743));
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1212 (.I0(n5_adj_5559), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[21] [7]), .I3(n60808), .O(n66739));
    defparam i4_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_4_lut_adj_1213 (.I0(\data_out_frame[11] [7]), .I1(n66851), 
            .I2(\data_out_frame[12] [1]), .I3(n66725), .O(n20_adj_5561));
    defparam i8_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_4_lut_adj_1214 (.I0(n26058), .I1(n26459), .I2(\data_out_frame[13] [7]), 
            .I3(n66809), .O(n19_adj_5562));
    defparam i7_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1215 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [4]), .I3(n61358), .O(n21_adj_5563));
    defparam i9_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1216 (.I0(\data_out_frame[14] [1]), .I1(n21_adj_5563), 
            .I2(n19_adj_5562), .I3(n20_adj_5561), .O(n61645));
    defparam i1_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1217 (.I0(n61645), .I1(n27087), .I2(n26781), 
            .I3(n1699), .O(n66521));
    defparam i3_4_lut_adj_1217.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(n61645), .I1(n60585), .I2(GND_net), 
            .I3(GND_net), .O(n60780));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26617));
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_out_frame[18] [4]), .I1(n60658), 
            .I2(GND_net), .I3(GND_net), .O(n60666));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1221 (.I0(n61543), .I1(n60666), .I2(n26617), 
            .I3(n6_adj_5564), .O(n25417));
    defparam i4_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 n78921_bdd_4_lut (.I0(n78921), .I1(n78588), .I2(n7_adj_12), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n78921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5566));
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1223 (.I0(n25417), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [5]), .I3(n6_adj_5566), .O(n66797));
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[15] [4]), .I1(n61318), 
            .I2(GND_net), .I3(GND_net), .O(n66453));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1225 (.I0(n66669), .I1(n66196), .I2(n27192), 
            .I3(n66806), .O(n10_adj_5567));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1226 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25857), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n4));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1226.LUT_INIT = 16'hfff4;
    SB_LUT4 i2_3_lut_adj_1227 (.I0(n68798), .I1(\data_out_frame[15] [3]), 
            .I2(n26087), .I3(GND_net), .O(n66438));
    defparam i2_3_lut_adj_1227.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(n61760), .I1(n66438), .I2(\data_out_frame[17] [5]), 
            .I3(GND_net), .O(n60581));
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1229 (.I0(\data_out_frame[17] [7]), .I1(n27182), 
            .I2(GND_net), .I3(GND_net), .O(n66794));
    defparam i2_2_lut_adj_1229.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(n65754), .I1(control_mode_c[4]), .I2(control_mode_c[3]), 
            .I3(control_mode_c[2]), .O(n25794));
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_out_frame[18] [0]), .I1(n66604), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5568));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1232 (.I0(\data_out_frame[19] [7]), .I1(n60581), 
            .I2(n61318), .I3(n6_adj_5568), .O(n68553));
    defparam i4_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n68553), .I3(GND_net), .O(n68217));
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(byte_transmit_counter[1]), 
            .O(n78915));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n78915_bdd_4_lut (.I0(n78915), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71761));
    defparam n78915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_63003 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(byte_transmit_counter[1]), 
            .O(n78909));
    defparam byte_transmit_counter_0__bdd_4_lut_63003.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_3_lut (.I0(n5_adj_5559), .I1(n60767), .I2(\data_out_frame[21] [6]), 
            .I3(GND_net), .O(n66447));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1234 (.I0(n10_adj_5508), .I1(n3474), 
            .I2(n161), .I3(reset), .O(n66103));
    defparam i1_2_lut_3_lut_4_lut_adj_1234.LUT_INIT = 16'hffbf;
    SB_LUT4 i3_4_lut_adj_1235 (.I0(n66739), .I1(\data_out_frame[23] [7]), 
            .I2(n60767), .I3(n26743), .O(n24039));
    defparam i3_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1236 (.I0(\data_out_frame[21] [2]), .I1(n60988), 
            .I2(n66571), .I3(GND_net), .O(n60565));
    defparam i1_2_lut_3_lut_adj_1236.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1237 (.I0(n10_adj_5508), .I1(n3474), 
            .I2(n161), .I3(n8_adj_13), .O(n28674));
    defparam i1_2_lut_3_lut_4_lut_adj_1237.LUT_INIT = 16'hffbf;
    SB_LUT4 i7_4_lut_adj_1238 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [0]), 
            .I2(n66447), .I3(n68217), .O(n18));
    defparam i7_4_lut_adj_1238.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1239 (.I0(n66616), .I1(n26898), .I2(n66391), 
            .I3(n60810), .O(n19_adj_5570));
    defparam i8_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1240 (.I0(n19_adj_5570), .I1(n69046), .I2(n18), 
            .I3(n12_adj_5571), .O(n68158));
    defparam i10_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 add_1194_9_lut (.I0(n65826), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n58266), .O(n65830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1194_8_lut (.I0(n65826), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n58265), .O(n65829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12_4_lut_adj_1241 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(n26605), .I3(\data_out_frame[24] [6]), .O(n28));
    defparam i12_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1242 (.I0(n66716), .I1(n60810), .I2(\data_out_frame[24] [5]), 
            .I3(\data_out_frame[23] [5]), .O(n26_adj_5572));
    defparam i10_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1243 (.I0(n66821), .I1(n68158), .I2(n66378), 
            .I3(\data_out_frame[23] [7]), .O(n27_adj_5573));
    defparam i11_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1244 (.I0(n60687), .I1(n61605), .I2(\data_out_frame[24] [1]), 
            .I3(\data_out_frame[24] [7]), .O(n25));
    defparam i9_4_lut_adj_1244.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27_adj_5573), .I2(n26_adj_5572), 
            .I3(n28), .O(n61583));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_1194_8 (.CI(n58265), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n58266));
    SB_LUT4 i1_2_lut_3_lut_adj_1245 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n66619));
    defparam i1_2_lut_3_lut_adj_1245.LUT_INIT = 16'h9696;
    SB_LUT4 add_1194_7_lut (.I0(n65826), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n58264), .O(n65834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_7 (.CI(n58264), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n58265));
    SB_LUT4 add_1194_6_lut (.I0(n65826), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n58263), .O(n65833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_6 (.CI(n58263), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n58264));
    SB_LUT4 add_1194_5_lut (.I0(n65826), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n58262), .O(n65832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_5 (.CI(n58262), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n58263));
    SB_LUT4 add_1194_4_lut (.I0(n65826), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n58261), .O(n65827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_4 (.CI(n58261), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n58262));
    SB_LUT4 add_1194_3_lut (.I0(n65826), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n58260), .O(n65831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_3 (.CI(n58260), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n58261));
    SB_LUT4 add_1194_2_lut (.I0(n65826), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n65828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n58260));
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n66206));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1247 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[5] [3]), .O(n66628));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [1]), .I3(GND_net), .O(n66760));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1249 (.I0(n66824), .I1(n24043), .I2(n66515), 
            .I3(n25456), .O(n14_adj_5574));
    defparam i6_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1250 (.I0(\data_out_frame[25] [7]), .I1(n66728), 
            .I2(n61583), .I3(n24039), .O(n13_c));
    defparam i5_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_209_i3_3_lut (.I0(n13_c), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n14_adj_5574), .I3(GND_net), .O(n3_adj_5546));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_209_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(n27256), .I1(n66531), .I2(GND_net), 
            .I3(GND_net), .O(n66779));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66450));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1253 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5575));
    defparam i2_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1254 (.I0(n7_adj_5575), .I1(\data_out_frame[15] [2]), 
            .I2(n60592), .I3(n68798), .O(n68678));
    defparam i4_4_lut_adj_1254.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1255 (.I0(\data_out_frame[11] [5]), .I1(n60445), 
            .I2(n27087), .I3(GND_net), .O(n18_adj_5576));
    defparam i1_2_lut_4_lut_adj_1255.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1256 (.I0(\data_out_frame[19] [4]), .I1(n68678), 
            .I2(n66594), .I3(\data_out_frame[17] [2]), .O(n60767));
    defparam i3_4_lut_adj_1256.LUT_INIT = 16'h9669;
    SB_LUT4 n78909_bdd_4_lut (.I0(n78909), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(byte_transmit_counter[1]), 
            .O(n71764));
    defparam n78909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26659));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1258 (.I0(n66641), .I1(n66181), .I2(\data_out_frame[12] [6]), 
            .I3(n66800), .O(n10_adj_5577));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1259 (.I0(n66190), .I1(n10_adj_5577), .I2(\data_out_frame[10] [5]), 
            .I3(GND_net), .O(n60592));   // verilog/coms.v(76[16:42])
    defparam i5_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1260 (.I0(\data_out_frame[15] [0]), .I1(n27290), 
            .I2(n60592), .I3(\data_out_frame[16] [7]), .O(n60646));
    defparam i3_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_out_frame[17] [0]), .I1(n27256), 
            .I2(GND_net), .I3(GND_net), .O(n66748));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1262 (.I0(n66757), .I1(n66836), .I2(n66463), 
            .I3(n66803), .O(n6_adj_5578));
    defparam i1_2_lut_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[6] [0]), .I1(n66866), .I2(n10_adj_5579), 
            .I3(n66181), .O(n66622));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14112_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3474), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n28323));   // verilog/coms.v(158[12:15])
    defparam i14112_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i5_4_lut_adj_1263 (.I0(n34), .I1(n66647), .I2(\data_out_frame[8] [7]), 
            .I3(\data_out_frame[11] [1]), .O(n12_adj_5580));
    defparam i5_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1264 (.I0(n26811), .I1(n12_adj_5580), .I2(\data_out_frame[15] [5]), 
            .I3(n66240), .O(n66231));
    defparam i6_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(n61318), .I1(n66231), .I2(GND_net), 
            .I3(GND_net), .O(n61533));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1266 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(n66628), .I3(n6_adj_5581), .O(n60778));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(n60778), .I1(n66503), .I2(GND_net), 
            .I3(GND_net), .O(n66504));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66251));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66356));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n66800));
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i30034_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n44122));   // verilog/coms.v(105[12:33])
    defparam i30034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5582));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1272 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [2]), 
            .I2(n26732), .I3(n6_adj_5582), .O(n66647));
    defparam i4_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1273 (.I0(\data_out_frame[8] [3]), .I1(n1668), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[10] [4]), .O(n66725));
    defparam i3_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16_2_lut (.I0(deadband[19]), .I1(n460), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1274 (.I0(n26732), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [4]), .I3(n26478), .O(n12_adj_5583));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1275 (.I0(\data_out_frame[9] [3]), .I1(n12_adj_5583), 
            .I2(n27211), .I3(n1130), .O(n26781));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1276 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n26062));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1276.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1277 (.I0(\data_out_frame[6] [6]), .I1(n66388), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n27211));
    defparam i1_2_lut_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1278 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n26058));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1279 (.I0(n66372), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[10] [6]), .I3(n66725), .O(n10_adj_5584));
    defparam i4_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1280 (.I0(\data_out_frame[13] [0]), .I1(n66304), 
            .I2(n10_adj_5584), .I3(n29_adj_5585), .O(n61751));
    defparam i1_4_lut_adj_1280.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(n66647), .I1(n26062), .I2(n27211), 
            .I3(n66806), .O(n10_adj_5586));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1282 (.I0(n61318), .I1(\data_out_frame[11] [5]), 
            .I2(n60445), .I3(n26781), .O(n26941));
    defparam i1_2_lut_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1283 (.I0(n26459), .I1(n66375), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n27087));
    defparam i2_3_lut_adj_1283.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1284 (.I0(n66631), .I1(n27004), .I2(\data_out_frame[11] [4]), 
            .I3(n66742), .O(n10_adj_5587));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1285 (.I0(\data_out_frame[13] [5]), .I1(n66200), 
            .I2(n10_adj_5587), .I3(\data_out_frame[11] [3]), .O(n27182));
    defparam i1_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1286 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(n26058), .O(n66806));
    defparam i2_3_lut_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27192));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_out_frame[5] [4]), .I1(n66654), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5588));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1289 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[10] [0]), 
            .I2(n26459), .I3(GND_net), .O(n6_adj_5581));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1290 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[4] [0]), 
            .I2(n66206), .I3(n6_adj_5588), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1290.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1291 (.I0(n66757), .I1(n66836), .I2(n66463), 
            .I3(GND_net), .O(n26067));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1291.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1292 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66228));
    defparam i1_2_lut_adj_1292.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1293 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(n66782), .I3(\data_out_frame[19] [1]), .O(n66474));
    defparam i2_3_lut_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1294 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[6] [1]), .O(n66654));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1295 (.I0(n66228), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[9] [3]), .I3(n66619), .O(n10_adj_5589));
    defparam i4_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1296 (.I0(\data_out_frame[9] [4]), .I1(n10_adj_5589), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n60445));
    defparam i5_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1297 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [3]), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1297.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1298 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66631));
    defparam i1_2_lut_adj_1298.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1299 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n27004));
    defparam i2_3_lut_adj_1299.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5436));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1300 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(\data_out_frame[17] [0]), 
            .O(n66531));
    defparam i2_3_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66669));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5435));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5434));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19851_3_lut (.I0(n38), .I1(n460), .I2(n486), .I3(GND_net), 
            .O(n40));
    defparam i19851_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i3_4_lut_adj_1302 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[7] [0]), .O(n66200));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5433));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1303 (.I0(\data_out_frame[8] [2]), .I1(n66866), 
            .I2(n66839), .I3(\data_out_frame[8] [4]), .O(n66190));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n66611));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_150_i2_4_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_150_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1305 (.I0(n26827), .I1(n66391), .I2(\data_out_frame[20] [5]), 
            .I3(n61765), .O(n66728));
    defparam i1_2_lut_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66304));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5585));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5430));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1308 (.I0(\data_out_frame[5] [0]), .I1(n26051), 
            .I2(n66342), .I3(n29_adj_5585), .O(n66388));   // verilog/coms.v(74[16:62])
    defparam i3_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1309 (.I0(\data_out_frame[6] [4]), .I1(n66372), 
            .I2(n26062), .I3(GND_net), .O(n26811));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1309.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1310 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[6] [1]), 
            .I2(n27211), .I3(n26058), .O(n24_adj_5590));
    defparam i10_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1311 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n17_adj_5591));
    defparam i3_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1312 (.I0(n66818), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [7]), .I3(n66304), .O(n22_adj_5592));
    defparam i8_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1313 (.I0(n17_adj_5591), .I1(n24_adj_5590), .I2(n66611), 
            .I3(\data_out_frame[5] [5]), .O(n26_adj_5593));
    defparam i12_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1314 (.I0(\data_out_frame[9] [6]), .I1(n66190), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5594));
    defparam i2_2_lut_adj_1314.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1315 (.I0(n66441), .I1(n66200), .I2(n66669), 
            .I3(\data_out_frame[5] [4]), .O(n14_adj_5595));
    defparam i6_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[4] [4]), .I1(n26_adj_5593), .I2(n22_adj_5592), 
            .I3(n27004), .O(n69125));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1316 (.I0(n69125), .I1(n14_adj_5595), .I2(n10_adj_5594), 
            .I3(\data_out_frame[9] [4]), .O(n68714));
    defparam i7_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1317 (.I0(\data_out_frame[9] [0]), .I1(n66631), 
            .I2(n26811), .I3(\data_out_frame[9] [5]), .O(n12_adj_5596));
    defparam i5_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1318 (.I0(\data_out_frame[9] [2]), .I1(n12_adj_5596), 
            .I2(n68714), .I3(n66169), .O(n61520));
    defparam i6_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(n61520), .I1(n26811), .I2(GND_net), 
            .I3(GND_net), .O(n61566));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66196));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(n27182), .I3(GND_net), .O(n66604));
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27056));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1323 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5597));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1324 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(n27056), .I3(\data_out_frame[11] [6]), .O(n14_adj_5598));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1325 (.I0(n66196), .I1(n14_adj_5598), .I2(n10_adj_5597), 
            .I3(n61566), .O(n66803));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1325.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(n26087), .I1(\data_out_frame[15] [4]), 
            .I2(n61318), .I3(\data_out_frame[15] [5]), .O(n61760));
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n66836));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\data_out_frame[10] [3]), .I1(n26058), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5599));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1329 (.I0(n29_adj_5585), .I1(n1193), .I2(n26062), 
            .I3(n6_adj_5599), .O(n66641));   // verilog/coms.v(76[16:42])
    defparam i4_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(88[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1193));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1331 (.I0(\data_out_frame[8] [3]), .I1(n26062), 
            .I2(\data_out_frame[6] [1]), .I3(n1193), .O(n66644));
    defparam i3_4_lut_adj_1331.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1332 (.I0(n66641), .I1(\data_out_frame[12] [2]), 
            .I2(n66836), .I3(n66803), .O(n16_adj_5600));
    defparam i6_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1333 (.I0(n60445), .I1(n66812), .I2(n66851), 
            .I3(n66654), .O(n17_adj_5601));
    defparam i7_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1334 (.I0(n17_adj_5601), .I1(n1668), .I2(n16_adj_5600), 
            .I3(\data_out_frame[10] [1]), .O(n60693));
    defparam i9_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66181));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66463));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1337 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [0]), 
            .I2(n10_adj_5567), .I3(\data_out_frame[6] [6]), .O(n26087));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n66839));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1339 (.I0(\data_out_frame[14] [6]), .I1(n66839), 
            .I2(n66463), .I3(\data_out_frame[6] [1]), .O(n10_adj_5579));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1340 (.I0(n60693), .I1(\data_out_frame[11] [5]), 
            .I2(n66644), .I3(n6_adj_5578), .O(n61358));
    defparam i4_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1341 (.I0(\data_out_frame[14] [5]), .I1(n1516), 
            .I2(n66325), .I3(\data_out_frame[12] [4]), .O(n27290));
    defparam i1_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1342 (.I0(n40_adj_5602), .I1(\data_out_frame[10] [2]), 
            .I2(n61520), .I3(n26459), .O(n68749));
    defparam i3_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1343 (.I0(\data_out_frame[10] [5]), .I1(n26067), 
            .I2(n61566), .I3(n26910), .O(n67902));
    defparam i3_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1344 (.I0(n1699), .I1(\data_out_frame[14] [4]), 
            .I2(n60585), .I3(n18_adj_5576), .O(n30));
    defparam i13_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1345 (.I0(n68798), .I1(n27290), .I2(n61358), 
            .I3(n66622), .O(n28_adj_5603));
    defparam i11_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1346 (.I0(\data_out_frame[12] [7]), .I1(n1720), 
            .I2(n61751), .I3(n26941), .O(n29_adj_5604));
    defparam i12_4_lut_adj_1346.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1347 (.I0(n61645), .I1(n60585), .I2(n66521), 
            .I3(n26473), .O(n60658));
    defparam i2_3_lut_4_lut_adj_1347.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1348 (.I0(n66503), .I1(n66800), .I2(\data_out_frame[14] [1]), 
            .I3(n60693), .O(n27_adj_5605));
    defparam i10_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1349 (.I0(n27_adj_5605), .I1(n29_adj_5604), .I2(n28_adj_5603), 
            .I3(n30), .O(n68184));
    defparam i16_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1350 (.I0(n66356), .I1(n27182), .I2(n66251), 
            .I3(\data_out_frame[15] [5]), .O(n14_adj_5606));
    defparam i6_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1351 (.I0(n1835), .I1(n27290), .I2(\data_out_frame[15] [4]), 
            .I3(n68184), .O(n13_adj_5607));
    defparam i5_4_lut_adj_1351.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1352 (.I0(n13_adj_5607), .I1(\data_out_frame[16] [0]), 
            .I2(n14_adj_5606), .I3(n61533), .O(n26590));
    defparam i2_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1353 (.I0(\data_out_frame[16] [4]), .I1(n27290), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n68332));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1354 (.I0(n26590), .I1(n68332), .I2(n66504), 
            .I3(n26309), .O(n60763));
    defparam i3_4_lut_adj_1354.LUT_INIT = 16'h9669;
    SB_LUT4 i15803_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n30015));
    defparam i15803_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15883_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n30095));
    defparam i15883_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15800_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n30012));
    defparam i15800_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15795_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n30007));
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26473));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i15790_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n30002));
    defparam i15790_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15906_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n30118));
    defparam i15906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66812));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66818));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1358 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n66169));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1358.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1359 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66866));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66757));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i15766_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29978));
    defparam i15766_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1361 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5609));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'h6666;
    SB_LUT4 i15748_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29960));
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1362 (.I0(n66757), .I1(n66628), .I2(n66760), 
            .I3(n6_adj_5609), .O(n66325));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i15958_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n30170));
    defparam i15958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15961_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n30173));
    defparam i15961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1363 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40_adj_5602));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1363.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1364 (.I0(\data_out_frame[12] [2]), .I1(n66650), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[5] [6]), .O(n66809));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\data_out_frame[14] [4]), .I1(n66325), 
            .I2(GND_net), .I3(GND_net), .O(n66704));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26051));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h6666;
    SB_LUT4 i15964_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n30176));
    defparam i15964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15967_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n30179));
    defparam i15967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15970_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n30182));
    defparam i15970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15973_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n30185));
    defparam i15973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15976_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n30188));
    defparam i15976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15979_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n30191));
    defparam i15979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66742));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1368 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n66441));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1369 (.I0(n66441), .I1(n66742), .I2(\data_out_frame[9] [5]), 
            .I3(GND_net), .O(n26459));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i16008_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n30220));
    defparam i16008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(n66571), .I1(n10_adj_5481), .I2(\data_out_frame[16] [3]), 
            .I3(n26617), .O(n66435));
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i16011_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n30223));
    defparam i16011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16014_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n30226));
    defparam i16014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16017_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n30229));
    defparam i16017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1371 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n66650));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1372 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n66342));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i29_2_lut (.I0(\data_out_frame[10] [0]), .I1(n26459), .I2(GND_net), 
            .I3(GND_net), .O(n26910));
    defparam i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5611));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i16020_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n30232));
    defparam i16020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16023_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n30235));
    defparam i16023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1374 (.I0(n66619), .I1(\data_out_frame[4] [7]), 
            .I2(n26478), .I3(n6_adj_5611), .O(n66375));
    defparam i4_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i16026_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n30238));
    defparam i16026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16029_3_lut_4_lut (.I0(n8_adj_9), .I1(n66103), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n30241));
    defparam i16029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1375 (.I0(\data_out_frame[7] [6]), .I1(n66375), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5612));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1375.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1376 (.I0(n26910), .I1(n66342), .I2(n66650), 
            .I3(\data_out_frame[9] [7]), .O(n14_adj_5613));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1377 (.I0(\data_out_frame[14] [2]), .I1(n14_adj_5613), 
            .I2(n10_adj_5612), .I3(n66812), .O(n60585));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1378 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [5]), 
            .I2(n26473), .I3(\data_out_frame[16] [7]), .O(n26309));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1379 (.I0(n60763), .I1(n26590), .I2(\data_out_frame[18] [7]), 
            .I3(GND_net), .O(n66782));
    defparam i2_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(n27256), .I1(n60585), .I2(GND_net), 
            .I3(GND_net), .O(n61543));
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 equal_305_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_9));   // verilog/coms.v(157[7:23])
    defparam equal_305_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1381 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[16] [6]), 
            .I2(n6_adj_5614), .I3(n66748), .O(n66571));
    defparam i1_4_lut_adj_1381.LUT_INIT = 16'h9669;
    SB_LUT4 equal_304_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam equal_304_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i3_4_lut_adj_1382 (.I0(n61543), .I1(n66782), .I2(\data_out_frame[18] [6]), 
            .I3(n26309), .O(n60988));
    defparam i3_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(n60988), .I1(n66571), .I2(GND_net), 
            .I3(GND_net), .O(n66572));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h6666;
    SB_LUT4 i14513_3_lut_4_lut (.I0(n10_adj_5508), .I1(n66982), .I2(reset), 
            .I3(n8_adj_5608), .O(n66992));
    defparam i14513_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n65826));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut_adj_1384 (.I0(\data_out_frame[21] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(n26659), .I3(n6_adj_5615), .O(n61070));
    defparam i4_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1385 (.I0(\data_out_frame[16] [2]), .I1(n66521), 
            .I2(\data_out_frame[16] [1]), .I3(n60698), .O(n60269));
    defparam i2_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1386 (.I0(n60778), .I1(n66503), .I2(n60988), 
            .I3(n66491), .O(n66587));
    defparam i1_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66672));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1388 (.I0(n60565), .I1(n61070), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n68828));
    defparam i2_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i51252_3_lut_4_lut (.I0(n10_adj_5508), .I1(n66982), .I2(n8), 
            .I3(reset), .O(n67037));
    defparam i51252_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_adj_1389 (.I0(\data_out_frame[23] [6]), .I1(n60767), 
            .I2(GND_net), .I3(GND_net), .O(n66821));
    defparam i1_2_lut_adj_1389.LUT_INIT = 16'h6666;
    SB_LUT4 i59190_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74422));   // verilog/coms.v(158[12:15])
    defparam i59190_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut_adj_1390 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n66131), .I3(LED_c), .O(n27768));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1390.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1391 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3474));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1391.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_306_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5508));   // verilog/coms.v(158[12:15])
    defparam equal_306_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_314_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5387));   // verilog/coms.v(158[12:15])
    defparam equal_314_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i58953_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74427));   // verilog/coms.v(158[12:15])
    defparam i58953_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1392 (.I0(\data_out_frame[21] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(n66779), .I3(n6_adj_5397), .O(n68518));
    defparam i4_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1393 (.I0(\FRAME_MATCHER.i[4] ), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(\FRAME_MATCHER.i[3] ), 
            .O(n82));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1393.LUT_INIT = 16'h0008;
    SB_LUT4 i23449_3_lut_4_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10]_c [1]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30772));
    defparam i23449_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i23437_3_lut_4_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10]_c [2]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30771));
    defparam i23437_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_787_Select_208_i3_4_lut (.I0(n68828), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5616), .I3(n66672), .O(n3_adj_5545));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1394 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5544));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1394.LUT_INIT = 16'ha088;
    SB_LUT4 i2_2_lut_3_lut_adj_1395 (.I0(\data_out_frame[18] [4]), .I1(n60658), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n7_adj_5469));
    defparam i2_2_lut_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1396 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [6]), 
            .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5543));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1396.LUT_INIT = 16'ha088;
    SB_LUT4 i23415_3_lut_4_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10]_c [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30768));
    defparam i23415_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_787_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5542));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5541));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i59009_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74430));   // verilog/coms.v(158[12:15])
    defparam i59009_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1397 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[20] [2]), 
            .I2(n61643), .I3(n61605), .O(n66515));
    defparam i1_2_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i62104_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n45273), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i62104_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_4_lut_adj_1398 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n45273), .I3(\FRAME_MATCHER.i_31__N_2511 ), .O(n25857));
    defparam i1_3_lut_4_lut_adj_1398.LUT_INIT = 16'hef00;
    SB_LUT4 i2_3_lut_4_lut_adj_1399 (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(\FRAME_MATCHER.i_31__N_2511 ), .I3(n45273), .O(n68152));
    defparam i2_3_lut_4_lut_adj_1399.LUT_INIT = 16'h1000;
    SB_LUT4 select_787_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1400 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1949), .I3(n1952), .O(n25866));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1400.LUT_INIT = 16'h4000;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(n1949), .I1(n4452), .I2(n1952), 
            .I3(n1955), .O(n68081));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h2000;
    SB_LUT4 i19_2_lut (.I0(pwm_setpoint[8]), .I1(\pwm_counter[8] ), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/pwm.v(11[19:30])
    defparam i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18_2_lut (.I0(pwm_setpoint[6]), .I1(\pwm_counter[6] ), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/pwm.v(11[19:30])
    defparam i18_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1949), .I1(n4452), .I2(n4), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n67901));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_3_lut_4_lut_adj_1402 (.I0(\data_in_frame[1] [4]), .I1(n66318), 
            .I2(n61665), .I3(n66481), .O(n69075));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1403 (.I0(\data_in_frame[1] [4]), .I1(n66318), 
            .I2(n66680), .I3(n66254), .O(n26315));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1404 (.I0(n27050), .I1(n27046), .I2(n26716), 
            .I3(n66815), .O(n6_adj_5619));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(n27050), .I1(n27046), .I2(n26716), 
            .I3(n66216), .O(n26673));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(n26722), .I1(n66686), .I2(n26719), 
            .I3(GND_net), .O(n66666));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1407 (.I0(n26722), .I1(n66686), .I2(\data_in_frame[6] [5]), 
            .I3(n66362), .O(Kp_23__N_974));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i61019_3_lut (.I0(n78864), .I1(n78546), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n76854));
    defparam i61019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_212_i3_3_lut_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\data_out_frame[24] [2]), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n66728), .O(n3_adj_5547));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_212_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in_frame[1] [5]), .I1(n66394), .I2(\data_in_frame[7] [7]), 
            .I3(\data_in_frame[4] [1]), .O(n18_adj_5620));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1408 (.I0(\data_in_frame[1] [5]), .I1(n66394), 
            .I2(\data_in_frame[7] [7]), .I3(\data_in_frame[5] [7]), .O(n66701));
    defparam i1_2_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1409 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [1]), 
            .I2(encoder0_position[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1409.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(\data_in_frame[9] [6]), .I1(n66719), 
            .I2(\data_in_frame[10][0] ), .I3(\data_in_frame[11] [7]), .O(n66842));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1411 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [7]), 
            .I2(encoder0_position[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1411.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_adj_1412 (.I0(\data_in_frame[9] [6]), .I1(n66719), 
            .I2(\data_in_frame[10][0] ), .I3(\data_in_frame[12] [2]), .O(n66625));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n26816), .I1(n4_adj_5621), .I2(\data_in_frame[10]_c [4]), 
            .I3(GND_net), .O(n26424));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62998 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n78897));
    defparam byte_transmit_counter_0__bdd_4_lut_62998.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1414 (.I0(n26816), .I1(n4_adj_5621), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(n71165));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1415 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[8] [7]), .I3(\data_in_frame[11] [3]), .O(n66815));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1416 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n66301));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1416.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1417 (.I0(n27115), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [4]), .I3(\data_in_frame[9] [3]), .O(n26362));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i58926_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74433));   // verilog/coms.v(158[12:15])
    defparam i58926_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5527));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14230_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n28441));   // verilog/coms.v(109[34:55])
    defparam i14230_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(n61180), .I3(GND_net), .O(n66479));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i55935_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71770));
    defparam i55935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55936_4_lut (.I0(n71770), .I1(n28441), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n71771));
    defparam i55936_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_3_lut_4_lut_adj_1419 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [5]), 
            .I2(n66244), .I3(n66695), .O(n70987));
    defparam i1_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i55934_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n71769));
    defparam i55934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(n3474), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(n8), .I3(n82), .O(n76));
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h0200;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n18_adj_5622));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1421 (.I0(n26343), .I1(n27_adj_5623), .I2(n26957), 
            .I3(n61599), .O(n24165));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i61021_3_lut (.I0(n78810), .I1(n78642), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n76856));
    defparam i61021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5521));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1422 (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[13][6] ), 
            .I2(\data_in_frame[14] [2]), .I3(n10_adj_5624), .O(n66163));   // verilog/coms.v(88[17:28])
    defparam i5_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(n24043), .I2(\FRAME_MATCHER.state[3] ), .I3(n66549), .O(n3_adj_5548));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i58931_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74434));   // verilog/coms.v(158[12:15])
    defparam i58931_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[13][6] ), 
            .I2(n61308), .I3(GND_net), .O(n66459));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n66512), .I3(\data_in_frame[16] [0]), .O(n8_adj_5625));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1424 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n26758), .I3(n25479), .O(n71109));
    defparam i1_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1425 (.I0(control_mode_c[3]), .I1(control_mode_c[2]), 
            .I2(control_mode_c[4]), .I3(GND_net), .O(n22_adj_14));
    defparam i1_3_lut_adj_1425.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1426 (.I0(\control_mode[5] ), .I1(n22_adj_14), 
            .I2(\control_mode[7] ), .I3(\control_mode[6] ), .O(n35278));   // verilog/coms.v(130[12] 305[6])
    defparam i1_4_lut_adj_1426.LUT_INIT = 16'hfffe;
    SB_LUT4 select_787_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1427 (.I0(n60687), .I1(\data_out_frame[22] [5]), 
            .I2(\data_out_frame[20] [3]), .I3(n61306), .O(n61587));
    defparam i1_2_lut_4_lut_adj_1427.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\data_out_frame[22] [5]), .I1(\data_out_frame[20] [3]), 
            .I2(n61306), .I3(GND_net), .O(n66552));
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1429 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(\FRAME_MATCHER.i_31__N_2512 ), .I3(GND_net), .O(n6_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_adj_1429.LUT_INIT = 16'hfefe;
    SB_LUT4 i14987_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n29199));   // verilog/coms.v(130[12] 305[6])
    defparam i14987_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_787_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5424));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14981_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n29193));   // verilog/coms.v(130[12] 305[6])
    defparam i14981_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_787_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5423));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1430 (.I0(n66163), .I1(n66495), .I2(\data_in_frame[20] [6]), 
            .I3(\data_in_frame[21] [0]), .O(n70891));
    defparam i1_4_lut_adj_1430.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1431 (.I0(n21), .I1(n19), .I2(n20), .I3(n60670), 
            .O(n66546));
    defparam i1_2_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5421));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1432 (.I0(n27256), .I1(n66531), .I2(n10_adj_5377), 
            .I3(n66248), .O(n61315));
    defparam i5_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1433 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [0]), 
            .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5420));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1433.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1434 (.I0(n66485), .I1(n66634), .I2(n25588), 
            .I3(n70891), .O(n68740));
    defparam i1_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 n78897_bdd_4_lut (.I0(n78897), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n78900));
    defparam n78897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_out_frame[18] [5]), .I1(n60778), 
            .I2(n66503), .I3(GND_net), .O(n66518));
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1436 (.I0(n60648), .I1(n61749), .I2(n71109), 
            .I3(n60757), .O(n71115));
    defparam i1_4_lut_adj_1436.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1437 (.I0(n60291), .I1(n71115), .I2(Kp_23__N_1564), 
            .I3(n66486), .O(n66713));
    defparam i1_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1438 (.I0(n66212), .I1(n66369), .I2(n66577), 
            .I3(\data_in_frame[15] [7]), .O(n71253));
    defparam i1_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1439 (.I0(n61589), .I1(n66407), .I2(n71253), 
            .I3(n26870), .O(n71259));
    defparam i1_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1440 (.I0(n66488), .I1(n66788), .I2(n68353), 
            .I3(n71259), .O(n60648));
    defparam i1_4_lut_adj_1440.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1441 (.I0(n60291), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n66833));
    defparam i2_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1442 (.I0(\data_in_frame[0][3] ), .I1(n66359), 
            .I2(n26750), .I3(\data_in_frame[4] [4]), .O(n26719));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1443 (.I0(\data_in_frame[0][3] ), .I1(n66359), 
            .I2(\data_in_frame[2][1] ), .I3(Kp_23__N_748), .O(n22_adj_5369));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut_4_lut_adj_1443.LUT_INIT = 16'h0990;
    SB_LUT4 select_787_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1444 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66273));
    defparam i1_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1445 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[19] [0]), 
            .I2(\data_in_frame[21] [1]), .I3(\data_in_frame[17] [7]), .O(n71217));
    defparam i1_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1446 (.I0(n66863), .I1(n66574), .I2(n71217), 
            .I3(n66273), .O(n71223));
    defparam i1_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(n66590), .I1(\data_in_frame[21] [4]), 
            .I2(n71223), .I3(\data_in_frame[21] [3]), .O(n71229));
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1448 (.I0(\data_in_frame[0][3] ), .I1(n66359), 
            .I2(n66254), .I3(\data_in_frame[8] [1]), .O(n14_adj_5627));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1449 (.I0(n66538), .I1(\data_in_frame[19] [7]), 
            .I2(n71229), .I3(n60628), .O(n71233));
    defparam i1_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1450 (.I0(n66833), .I1(n66429), .I2(n71233), 
            .I3(n66336), .O(n71239));
    defparam i1_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1451 (.I0(n26522), .I1(n71239), .I2(n66193), 
            .I3(n66683), .O(n71243));
    defparam i1_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(n68427), .I1(n66558), .I2(GND_net), 
            .I3(GND_net), .O(n66785));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1453 (.I0(n66785), .I1(n60648), .I2(n68895), 
            .I3(n71243), .O(n66384));
    defparam i1_4_lut_adj_1453.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1454 (.I0(\data_in_frame[21] [5]), .I1(n26537), 
            .I2(\data_in_frame[19] [5]), .I3(n61660), .O(n66336));
    defparam i3_4_lut_adj_1454.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1455 (.I0(\data_in_frame[20][0] ), .I1(\data_in_frame[19] [6]), 
            .I2(n61660), .I3(\data_in_frame[20][1] ), .O(n66538));
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n20_adj_5628), .I1(n61349), .I2(n66407), 
            .I3(\data_in_frame[16] [5]), .O(n66485));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5629));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1458 (.I0(\data_in_frame[18] [5]), .I1(n26794), 
            .I2(n27043), .I3(n6_adj_5629), .O(Kp_23__N_1564));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1459 (.I0(n161), .I1(n66108), .I2(n10_adj_5387), 
            .I3(reset), .O(n66150));
    defparam i1_2_lut_3_lut_4_lut_adj_1459.LUT_INIT = 16'hfffd;
    SB_LUT4 select_787_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1460 (.I0(\data_in_frame[16] [5]), .I1(n6), .I2(n66494), 
            .I3(n66500), .O(n66329));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1461 (.I0(\data_in_frame[13][7] ), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[10][6] ), .I3(\data_in_frame[15] [2]), .O(n71075));
    defparam i1_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1462 (.I0(\data_in_frame[16] [3]), .I1(n60656), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5631));
    defparam i2_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 i55550_3_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0][5] ), 
            .I2(\data_in_frame[0][6] ), .I3(n26722), .O(n71370));
    defparam i55550_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i1_4_lut_adj_1463 (.I0(n26843), .I1(Kp_23__N_1067), .I2(Kp_23__N_1389), 
            .I3(n71075), .O(n71081));
    defparam i1_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1464 (.I0(\data_out_frame[21] [5]), .I1(n60808), 
            .I2(\data_out_frame[22] [5]), .I3(GND_net), .O(n60810));
    defparam i1_2_lut_3_lut_adj_1464.LUT_INIT = 16'h9696;
    SB_LUT4 i61834_4_lut (.I0(\data_in_frame[12] [7]), .I1(n7_adj_5631), 
            .I2(\data_in_frame[15] [4]), .I3(n8_adj_5625), .O(n77669));
    defparam i61834_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_out_frame[21] [5]), .I1(n60808), 
            .I2(n66797), .I3(GND_net), .O(n12_adj_5571));
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1466 (.I0(n66329), .I1(n77669), .I2(n60656), 
            .I3(n71081), .O(n71087));
    defparam i1_4_lut_adj_1466.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1467 (.I0(n25588), .I1(n66580), .I2(n66524), 
            .I3(n71087), .O(n66788));
    defparam i1_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1468 (.I0(\data_out_frame[21] [5]), .I1(n60808), 
            .I2(n66821), .I3(n68518), .O(n8_adj_5616));
    defparam i3_3_lut_4_lut_adj_1468.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(Kp_23__N_1564), .I1(n66485), .I2(GND_net), 
            .I3(GND_net), .O(n66486));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27043));
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'h6666;
    SB_LUT4 i15762_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [1]), 
            .I3(\current_limit[1] ), .O(n29974));   // verilog/coms.v(130[12] 305[6])
    defparam i15762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1471 (.I0(n27043), .I1(n66486), .I2(\data_in_frame[19] [0]), 
            .I3(\data_in_frame[18] [2]), .O(n66634));
    defparam i1_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i15729_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [0]), 
            .I3(\current_limit[0] ), .O(n29941));   // verilog/coms.v(130[12] 305[6])
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15601_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29813));
    defparam i15601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21111_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1][0] ), 
            .I3(\control_mode[0] ), .O(n29940));   // verilog/coms.v(130[12] 305[6])
    defparam i21111_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15598_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29810));
    defparam i15598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15595_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29807));
    defparam i15595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16572_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20][0] ), 
            .I3(\current_limit[8] ), .O(n30784));   // verilog/coms.v(130[12] 305[6])
    defparam i16572_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16571_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20][1] ), 
            .I3(\current_limit[9] ), .O(n30783));   // verilog/coms.v(130[12] 305[6])
    defparam i16571_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1472 (.I0(n61349), .I1(n66634), .I2(n66683), 
            .I3(n71157), .O(Kp_23__N_1607));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_in_frame[16] [6]), .I1(n66329), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5633));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i15592_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29804));
    defparam i15592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1474 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[19] [1]), 
            .I2(n20_adj_5628), .I3(n6_adj_5633), .O(n26522));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i15770_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [5]), 
            .I3(\control_mode[5] ), .O(n29982));   // verilog/coms.v(130[12] 305[6])
    defparam i15770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1475 (.I0(\data_in_frame[17] [1]), .I1(n68908), 
            .I2(GND_net), .I3(GND_net), .O(n66580));
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1476 (.I0(n25505), .I1(n66580), .I2(\data_in_frame[19] [3]), 
            .I3(GND_net), .O(n68895));
    defparam i1_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1477 (.I0(\data_in_frame[14][6] ), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66577));
    defparam i1_2_lut_adj_1477.LUT_INIT = 16'h6666;
    SB_LUT4 i61830_4_lut (.I0(n61599), .I1(n66769), .I2(n66776), .I3(n66432), 
            .O(n77665));
    defparam i61830_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i15769_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1][6] ), 
            .I3(\control_mode[6] ), .O(n29981));   // verilog/coms.v(130[12] 305[6])
    defparam i15769_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1478 (.I0(n61577), .I1(n26424), .I2(n66677), 
            .I3(n71059), .O(n71065));
    defparam i1_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i16567_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20][2] ), 
            .I3(\current_limit[10] ), .O(n30779));   // verilog/coms.v(130[12] 305[6])
    defparam i16567_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23550_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20][3] ), 
            .I3(current_limit[11]), .O(n37697));   // verilog/coms.v(130[12] 305[6])
    defparam i23550_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1479 (.I0(n71065), .I1(n61658), .I2(n77665), 
            .I3(n30_adj_5634), .O(n68908));
    defparam i1_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1480 (.I0(n26537), .I1(n68908), .I2(\data_in_frame[19] [4]), 
            .I3(GND_net), .O(n68427));
    defparam i1_3_lut_adj_1480.LUT_INIT = 16'h6969;
    SB_LUT4 i15589_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29801));
    defparam i15589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21164_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [7]), 
            .I3(\control_mode[7] ), .O(n29977));   // verilog/coms.v(130[12] 305[6])
    defparam i21164_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15775_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n29987));   // verilog/coms.v(130[12] 305[6])
    defparam i15775_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16565_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20][4] ), 
            .I3(current_limit[12]), .O(n30777));   // verilog/coms.v(130[12] 305[6])
    defparam i16565_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15586_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29798));
    defparam i15586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(n60656), .I1(n26758), .I2(GND_net), 
            .I3(GND_net), .O(n66494));
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1482 (.I0(\data_in_frame[14] [2]), .I1(n61528), 
            .I2(GND_net), .I3(GND_net), .O(n61749));
    defparam i1_2_lut_adj_1482.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1483 (.I0(\data_in_frame[14]_c [3]), .I1(n27241), 
            .I2(n66301), .I3(n6_adj_5494), .O(n20_adj_5628));
    defparam i4_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1484 (.I0(\data_in_frame[16] [4]), .I1(n20_adj_5628), 
            .I2(n61749), .I3(n6), .O(n68457));
    defparam i3_4_lut_adj_1484.LUT_INIT = 16'h9669;
    SB_LUT4 i38961_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode_c[3]), .O(n29985));   // verilog/coms.v(130[12] 305[6])
    defparam i38961_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1485 (.I0(n66495), .I1(n68457), .I2(\data_in_frame[18] [6]), 
            .I3(GND_net), .O(n66279));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1485.LUT_INIT = 16'h9696;
    SB_LUT4 i23549_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20] [7]), 
            .I3(current_limit[15]), .O(n30773));   // verilog/coms.v(130[12] 305[6])
    defparam i23549_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15761_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [2]), 
            .I3(\current_limit[2] ), .O(n29973));   // verilog/coms.v(130[12] 305[6])
    defparam i15761_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i38974_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode_c[2]), .O(n53030));   // verilog/coms.v(130[12] 305[6])
    defparam i38974_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1486 (.I0(n66279), .I1(\data_in_frame[19] [0]), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n66193));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1486.LUT_INIT = 16'h9696;
    SB_LUT4 i23544_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20] [6]), 
            .I3(current_limit[14]), .O(n30775));   // verilog/coms.v(130[12] 305[6])
    defparam i23544_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15583_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29795));
    defparam i15583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15771_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode_c[4]), .O(n29983));   // verilog/coms.v(130[12] 305[6])
    defparam i15771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15758_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [5]), 
            .I3(\current_limit[5] ), .O(n29970));   // verilog/coms.v(130[12] 305[6])
    defparam i15758_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i23548_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[20] [5]), 
            .I3(current_limit[13]), .O(n30776));   // verilog/coms.v(130[12] 305[6])
    defparam i23548_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15541_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [6]), 
            .I3(\current_limit[6] ), .O(n29753));   // verilog/coms.v(130[12] 305[6])
    defparam i15541_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15580_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66099), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29792));
    defparam i15580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1487 (.I0(n26816), .I1(n69038), .I2(n26244), 
            .I3(n71189), .O(n66769));
    defparam i1_4_lut_adj_1487.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n71281));
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1489 (.I0(\data_in_frame[12] [6]), .I1(n71281), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[15] [2]), .O(n71285));
    defparam i1_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1490 (.I0(n26424), .I1(n66791), .I2(n26244), 
            .I3(n71285), .O(n61525));
    defparam i1_4_lut_adj_1490.LUT_INIT = 16'h6996;
    SB_LUT4 i15760_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [3]), 
            .I3(\current_limit[3] ), .O(n29972));   // verilog/coms.v(130[12] 305[6])
    defparam i15760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_adj_1491 (.I0(\data_in_frame[15] [3]), .I1(n61525), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n61660));
    defparam i1_3_lut_adj_1491.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1492 (.I0(n66524), .I1(n26378), .I2(\data_in_frame[17] [3]), 
            .I3(n66776), .O(n10_adj_5635));
    defparam i4_4_lut_adj_1492.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1493 (.I0(n61525), .I1(n10_adj_5635), .I2(n24165), 
            .I3(GND_net), .O(n26537));
    defparam i5_3_lut_adj_1493.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1494 (.I0(n61660), .I1(n68633), .I2(n68353), 
            .I3(\data_in_frame[17] [5]), .O(n68131));
    defparam i1_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i16079_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[10][7] ), .O(n30291));
    defparam i16079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15759_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [4]), 
            .I3(\current_limit[4] ), .O(n29971));   // verilog/coms.v(130[12] 305[6])
    defparam i15759_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16076_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[10][6] ), .O(n30288));
    defparam i16076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(\data_in_frame[15] [5]), .I1(n24165), 
            .I2(GND_net), .I3(GND_net), .O(n66590));
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i16072_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[10][5] ), .O(n30284));
    defparam i16072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(n68131), .I1(n26537), .I2(GND_net), 
            .I3(GND_net), .O(n27201));
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15513_3_lut_4_lut (.I0(n2872), .I1(n28088), .I2(\data_in_frame[21] [7]), 
            .I3(\current_limit[7] ), .O(n29725));   // verilog/coms.v(130[12] 305[6])
    defparam i15513_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1497 (.I0(n66857), .I1(\data_in_frame[11] [5]), 
            .I2(n66698), .I3(\data_in_frame[13][7] ), .O(n14_adj_5636));
    defparam i6_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1498 (.I0(n9_adj_5560), .I1(n14_adj_5636), .I2(n66827), 
            .I3(n61665), .O(n68646));
    defparam i7_4_lut_adj_1498.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1499 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66512));
    defparam i1_2_lut_adj_1499.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1500 (.I0(Kp_23__N_1256), .I1(n66512), .I2(n68646), 
            .I3(n61601), .O(n60757));
    defparam i3_4_lut_adj_1500.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62845 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[1]), .O(n78645));
    defparam byte_transmit_counter_0__bdd_4_lut_62845.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1501 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66751));
    defparam i1_2_lut_adj_1501.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1502 (.I0(n27_adj_5623), .I1(n66459), .I2(n66751), 
            .I3(\data_in_frame[13] [5]), .O(n61658));
    defparam i1_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i16066_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n30278));
    defparam i16066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(n26870), .I1(n61658), .I2(GND_net), 
            .I3(GND_net), .O(n66535));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i16059_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[10]_c [1]), .O(n30271));
    defparam i16059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1504 (.I0(\data_in_frame[11] [5]), .I1(n66535), 
            .I2(n26673), .I3(n61555), .O(Kp_23__N_1256));
    defparam i3_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1505 (.I0(Kp_23__N_1256), .I1(\data_in_frame[16] [0]), 
            .I2(\data_in_frame[17] [7]), .I3(n66597), .O(n10_adj_5480));
    defparam i4_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1506 (.I0(n66206), .I1(n66809), .I2(n40_adj_5602), 
            .I3(n66704), .O(n27256));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1507 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[16] [0]), 
            .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1507.LUT_INIT = 16'ha088;
    SB_LUT4 i5_3_lut_adj_1508 (.I0(n69038), .I1(n10_adj_5480), .I2(\data_in_frame[15] [5]), 
            .I3(GND_net), .O(n25479));
    defparam i5_3_lut_adj_1508.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1509 (.I0(n66206), .I1(n66809), .I2(n40_adj_5602), 
            .I3(\data_out_frame[14] [3]), .O(n66503));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1509.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_in_frame[18] [3]), .I1(n60757), 
            .I2(GND_net), .I3(GND_net), .O(n61778));
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i16056_3_lut_4_lut (.I0(n28674), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[10][0] ), .O(n30268));
    defparam i16056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1511 (.I0(n61778), .I1(\data_in_frame[20][3] ), 
            .I2(n66497), .I3(\data_in_frame[20][4] ), .O(n66429));
    defparam i3_4_lut_adj_1511.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1512 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66555));
    defparam i1_2_lut_adj_1512.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(n60664), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n66568));
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1514 (.I0(n66719), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[8] [4]), .O(n24_adj_5637));
    defparam i10_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1515 (.I0(n66689), .I1(\data_in_frame[1] [7]), 
            .I2(n66479), .I3(\data_in_frame[8] [3]), .O(n22_adj_5638));
    defparam i8_4_lut_adj_1515.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1516 (.I0(n66830), .I1(n24_adj_5637), .I2(n18_adj_5620), 
            .I3(\data_in_frame[6] [3]), .O(n26_adj_5639));
    defparam i12_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1517 (.I0(\data_in_frame[8] [0]), .I1(n26_adj_5639), 
            .I2(n22_adj_5638), .I3(\data_in_frame[8] [7]), .O(n66857));
    defparam i13_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1518 (.I0(\data_in_frame[2][3] ), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0][1] ), .I3(GND_net), .O(n26722));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1518.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1519 (.I0(n66842), .I1(n66686), .I2(n66722), 
            .I3(n66456), .O(n24_adj_5640));
    defparam i10_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1520 (.I0(\data_in_frame[2]_c [5]), .I1(\data_in_frame[0][3] ), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26188));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1520.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_4_lut_adj_1521 (.I0(n66857), .I1(n66692), .I2(n66216), 
            .I3(n61328), .O(n22_adj_5641));
    defparam i8_4_lut_adj_1521.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1522 (.I0(n66763), .I1(n24_adj_5640), .I2(n18_adj_5622), 
            .I3(n66568), .O(n26_adj_5642));
    defparam i12_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1523 (.I0(\data_in_frame[9] [7]), .I1(n26_adj_5642), 
            .I2(n22_adj_5641), .I3(n27071), .O(n61528));
    defparam i13_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1524 (.I0(n26362), .I1(n66401), .I2(GND_net), 
            .I3(GND_net), .O(n26843));
    defparam i1_2_lut_adj_1524.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13]_c [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5623));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_in_frame[13][7] ), .I1(n66734), 
            .I2(GND_net), .I3(GND_net), .O(n66597));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1527 (.I0(\data_in_frame[11] [6]), .I1(n24268), 
            .I2(n26098), .I3(n26846), .O(n66401));
    defparam i3_4_lut_adj_1527.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1528 (.I0(\data_in_frame[10]_c [1]), .I1(\data_in_frame[10]_c [4]), 
            .I2(\data_in_frame[11] [4]), .I3(\data_in_frame[12] [1]), .O(n70977));
    defparam i1_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 n78645_bdd_4_lut (.I0(n78645), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[1]), 
            .O(n78648));
    defparam n78645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1529 (.I0(n70977), .I1(n66315), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[11] [0]), .O(n70985));
    defparam i1_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1530 (.I0(n70985), .I1(n66815), .I2(n70987), 
            .I3(n70983), .O(n70993));
    defparam i1_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1531 (.I0(Kp_23__N_993), .I1(Kp_23__N_974), .I2(n24272), 
            .I3(n70993), .O(n70999));
    defparam i1_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1532 (.I0(n66565), .I1(n66860), .I2(n66322), 
            .I3(n70999), .O(n71005));
    defparam i1_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1533 (.I0(n66854), .I1(n61577), .I2(n66625), 
            .I3(n71005), .O(n61308));
    defparam i1_4_lut_adj_1533.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(\data_in_frame[13] [1]), .I1(n61308), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5643));
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1535 (.I0(n26416), .I1(\data_in_frame[13] [2]), 
            .I2(n66555), .I3(n6_adj_5643), .O(n66734));
    defparam i4_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1536 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[16] [0]), .I3(\data_in_frame[16] [1]), .O(n18_adj_5644));
    defparam i7_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1537 (.I0(n66401), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[13][6] ), .I3(\data_in_frame[13] [3]), .O(n19_adj_5645));
    defparam i8_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1538 (.I0(n19_adj_5645), .I1(n61601), .I2(n18_adj_5644), 
            .I3(n12_adj_5471), .O(n60723));
    defparam i10_4_lut_adj_1538.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1539 (.I0(n26843), .I1(n61528), .I2(\data_in_frame[14] [0]), 
            .I3(\data_in_frame[16] [2]), .O(n10_adj_5624));
    defparam i4_4_lut_adj_1539.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26794));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1541 (.I0(n66163), .I1(\data_in_frame[16] [3]), 
            .I2(n60723), .I3(GND_net), .O(n60628));
    defparam i2_3_lut_adj_1541.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1542 (.I0(n69038), .I1(n26957), .I2(GND_net), 
            .I3(GND_net), .O(n61599));
    defparam i1_2_lut_adj_1542.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1543 (.I0(n26343), .I1(n26362), .I2(GND_net), 
            .I3(GND_net), .O(n66432));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1543.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1544 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [7]), 
            .I2(\control_mode[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1544.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1545 (.I0(n26685), .I1(n26846), .I2(GND_net), 
            .I3(GND_net), .O(n27115));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1546 (.I0(n26244), .I1(n26329), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1546.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(n60607), .I1(n66312), .I2(GND_net), 
            .I3(GND_net), .O(n71177));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1548 (.I0(n71177), .I1(n26244), .I2(n25467), 
            .I3(\data_in_frame[9] [0]), .O(n61180));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1549 (.I0(n71165), .I1(n66860), .I2(n26673), 
            .I3(n7_adj_15), .O(n71171));
    defparam i1_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1550 (.I0(n66352), .I1(n66754), .I2(n66827), 
            .I3(n71171), .O(n25467));
    defparam i1_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26098));
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1552 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [6]), 
            .I2(\control_mode[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1552.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1553 (.I0(\data_in_frame[10][7] ), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66695));
    defparam i1_2_lut_adj_1553.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1554 (.I0(n26098), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [3]), .I3(n66301), .O(n66312));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1555 (.I0(n25467), .I1(n61180), .I2(n60607), 
            .I3(n71181), .O(n69038));
    defparam i1_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1556 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [5]), 
            .I2(\control_mode[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1556.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(GND_net), .I3(GND_net), .O(n27071));
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1558 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66315));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1558.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62988 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n78861));
    defparam byte_transmit_counter_0__bdd_4_lut_62988.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1559 (.I0(n26321), .I1(n66219), .I2(n66666), 
            .I3(n6_adj_5619), .O(n26343));
    defparam i4_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1560 (.I0(n66212), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66660));
    defparam i1_2_lut_adj_1560.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1561 (.I0(n26343), .I1(n26957), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_5634));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1561.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1562 (.I0(\data_in_frame[20][2] ), .I1(n30_adj_5634), 
            .I2(n66660), .I3(\data_in_frame[13]_c [4]), .O(n66863));
    defparam i3_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1563 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n71265));
    defparam i1_2_lut_adj_1563.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1564 (.I0(n68099), .I1(n61599), .I2(n71265), 
            .I3(\data_in_frame[13] [3]), .O(n68633));
    defparam i1_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i15983_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n30195));
    defparam i15983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [1]), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1566 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n66830));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1566.LUT_INIT = 16'h6666;
    SB_LUT4 i15986_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n30198));
    defparam i15986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(n66680), .I1(n66701), .I2(n66481), 
            .I3(n71295), .O(n26873));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(\data_in_frame[12] [5]), .I1(n26873), 
            .I2(GND_net), .I3(GND_net), .O(n66369));
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(n26873), .I1(n61123), .I2(GND_net), 
            .I3(GND_net), .O(n61577));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 n78861_bdd_4_lut (.I0(n78861), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n78864));
    defparam n78861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15989_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n30201));
    defparam i15989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1570 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[12] [6]), .I3(GND_net), .O(n66244));
    defparam i2_3_lut_adj_1570.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n71802), .I2(n71803), .I3(byte_transmit_counter[2]), .O(n78633));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i15992_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n30204));
    defparam i15992_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1571 (.I0(n60607), .I1(n27223), .I2(GND_net), 
            .I3(GND_net), .O(n66565));
    defparam i1_2_lut_adj_1571.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1572 (.I0(\data_in_frame[10][5] ), .I1(n26816), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n66322));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1572.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1573 (.I0(\data_in_frame[15] [0]), .I1(n26329), 
            .I2(\data_in_frame[14][7] ), .I3(n66322), .O(n66677));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(\data_in_frame[10]_c [1]), .I1(n26280), 
            .I2(n66565), .I3(\data_in_frame[9] [7]), .O(n27241));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'h9669;
    SB_LUT4 i15995_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n30207));
    defparam i15995_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15998_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n30210));
    defparam i15998_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16001_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n30213));
    defparam i16001_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1575 (.I0(\data_in_frame[8] [1]), .I1(n69075), 
            .I2(GND_net), .I3(GND_net), .O(n66854));
    defparam i1_2_lut_adj_1575.LUT_INIT = 16'h9999;
    SB_LUT4 i16005_3_lut_4_lut (.I0(n45146), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n30217));
    defparam i16005_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(n26777), .I1(n66701), .I2(n66318), 
            .I3(\data_in_frame[8] [0]), .O(n26280));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1577 (.I0(n26280), .I1(n66854), .I2(GND_net), 
            .I3(GND_net), .O(n66754));
    defparam i1_2_lut_adj_1577.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n61449), .I1(n66754), .I2(n24272), 
            .I3(\data_in_frame[10]_c [2]), .O(n61123));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1579 (.I0(n27241), .I1(n66677), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5647));
    defparam i1_2_lut_adj_1579.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1580 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[14][5] ), 
            .I2(n66244), .I3(n6_adj_5647), .O(n25505));
    defparam i4_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1581 (.I0(\data_in_frame[14][6] ), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5648));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1581.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1582 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[16] [6]), 
            .I2(n61589), .I3(n6_adj_5648), .O(n66500));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1582.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1583 (.I0(n66500), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5649));
    defparam i2_2_lut_adj_1583.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1584 (.I0(\data_in_frame[19] [2]), .I1(n26758), 
            .I2(n6_adj_5649), .I3(n25505), .O(n66558));
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16132_3_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n30344));
    defparam i16132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16128_3_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n30340));
    defparam i16128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1585 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[2][0] ), 
            .I2(n66264), .I3(n26750), .O(n66362));   // verilog/coms.v(76[16:42])
    defparam i3_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 n78633_bdd_4_lut (.I0(n78633), .I1(n71869), .I2(n71868), .I3(byte_transmit_counter[2]), 
            .O(n78636));
    defparam n78633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_2036_i7_2_lut (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_15));   // verilog/coms.v(239[9:81])
    defparam equal_2036_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1586 (.I0(\data_in_frame[8] [5]), .I1(n66362), 
            .I2(\data_in_frame[6] [3]), .I3(Kp_23__N_872), .O(n26244));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1587 (.I0(n26294), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_869), .I3(Kp_23__N_872), .O(n26329));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1587.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1588 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[2][6] ), .I3(GND_net), .O(n14_adj_5650));
    defparam i5_3_lut_adj_1588.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1589 (.I0(n66420), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[2]_c [5]), .I3(n66359), .O(n15_adj_5651));
    defparam i6_4_lut_adj_1589.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1590 (.I0(n15_adj_5651), .I1(\data_in_frame[2] [7]), 
            .I2(n14_adj_5650), .I3(\data_in_frame[4] [6]), .O(n26846));
    defparam i8_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66209));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1592 (.I0(n26306), .I1(\data_in_frame[1] [7]), 
            .I2(n66209), .I3(n6_adj_5402), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1592.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1593 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n66372));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1593.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1594 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n66456));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1594.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1595 (.I0(\data_in_frame[1] [7]), .I1(n66286), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [4]), .O(n66686));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i16125_3_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n30337));
    defparam i16125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1596 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[7] [5]), .I3(n26583), .O(n12_adj_5652));
    defparam i5_4_lut_adj_1596.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1597 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_5652), 
            .I2(n66276), .I3(\data_in_frame[5] [3]), .O(n60607));
    defparam i6_4_lut_adj_1597.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1598 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_869), 
            .I2(\data_in_frame[6] [2]), .I3(n26315), .O(n26816));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1599 (.I0(n26719), .I1(n66456), .I2(n26722), 
            .I3(n27050), .O(n26685));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1600 (.I0(\data_in_frame[8] [7]), .I1(Kp_23__N_993), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5653));
    defparam i2_2_lut_adj_1600.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(n26583), .I1(n66397), .I2(n66470), 
            .I3(\data_in_frame[7] [4]), .O(n66763));
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1602 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [6]), .O(n34));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1602.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1603 (.I0(n26137), .I1(\data_in_frame[7] [6]), 
            .I2(n26297), .I3(GND_net), .O(n24272));
    defparam i2_3_lut_adj_1603.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1604 (.I0(n27046), .I1(n66763), .I2(GND_net), 
            .I3(GND_net), .O(n24268));
    defparam i1_2_lut_adj_1604.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1605 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[12] [3]), .I3(GND_net), .O(n66851));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1605.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1606 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0][6] ), 
            .I2(\data_in_frame[1][0] ), .I3(\data_in_frame[3] [2]), .O(n66470));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1607 (.I0(\data_in_frame[5] [4]), .I1(n66470), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n26137));
    defparam i1_3_lut_adj_1607.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1608 (.I0(\data_in_frame[6] [7]), .I1(n26188), 
            .I2(GND_net), .I3(GND_net), .O(n27050));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1608.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1609 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n66622), .I3(n1516), .O(n27157));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1609.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1610 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n66219));
    defparam i1_2_lut_adj_1610.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1611 (.I0(\data_out_frame[8] [4]), .I1(n27192), 
            .I2(\data_out_frame[9] [0]), .I3(n10_adj_5586), .O(n1720));
    defparam i5_3_lut_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1612 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26306));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1612.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1613 (.I0(\data_out_frame[8] [4]), .I1(n27192), 
            .I2(n68749), .I3(\data_out_frame[12] [7]), .O(n14));
    defparam i5_3_lut_4_lut_adj_1613.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1614 (.I0(\data_out_frame[11] [5]), .I1(n60445), 
            .I2(n26781), .I3(GND_net), .O(n66608));
    defparam i1_2_lut_3_lut_adj_1614.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1615 (.I0(\data_in_frame[5] [6]), .I1(n26297), 
            .I2(GND_net), .I3(GND_net), .O(n66481));
    defparam i1_2_lut_adj_1615.LUT_INIT = 16'h6666;
    SB_LUT4 i16112_3_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n30324));
    defparam i16112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1616 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26777));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1616.LUT_INIT = 16'h6666;
    SB_LUT4 i16109_3_lut_4_lut (.I0(n28670), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n30321));
    defparam i16109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1617 (.I0(\data_out_frame[11] [5]), .I1(n60445), 
            .I2(n27182), .I3(n27087), .O(n60640));
    defparam i2_3_lut_4_lut_adj_1617.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1618 (.I0(n26777), .I1(n66481), .I2(n66254), 
            .I3(\data_in_frame[1] [4]), .O(n27223));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[16] [1]), .I1(n66474), .I2(\data_out_frame[16] [4]), 
            .I3(n27157), .O(n6_adj_5614));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1619 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26321));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_adj_1619.LUT_INIT = 16'h6666;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5610));
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_adj_1620 (.I0(\data_in_frame[6] [0]), .I1(n66365), 
            .I2(GND_net), .I3(GND_net), .O(n66722));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1620.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(Kp_23__N_799), .I1(n61328), .I2(n66722), 
            .I3(n70901), .O(n61665));
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1622 (.I0(\data_out_frame[16] [1]), .I1(n66474), 
            .I2(\data_out_frame[16] [4]), .I3(n60646), .O(n6_adj_5615));
    defparam i1_2_lut_4_lut_adj_1622.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(\data_in_frame[5] [5]), .I1(n26284), 
            .I2(n66175), .I3(\data_in_frame[0][7] ), .O(n66394));
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 i31069_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n45146));
    defparam i31069_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_adj_1624 (.I0(n66394), .I1(n61665), .I2(\data_in_frame[7] [7]), 
            .I3(GND_net), .O(n61449));
    defparam i1_3_lut_adj_1624.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62958 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n78849));
    defparam byte_transmit_counter_0__bdd_4_lut_62958.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1625 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5655));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1625.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1626 (.I0(n26188), .I1(Kp_23__N_767), .I2(\data_in_frame[0][7] ), 
            .I3(n26583), .O(n69112));   // verilog/coms.v(74[16:69])
    defparam i3_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1627 (.I0(n69112), .I1(n27046), .I2(n66404), 
            .I3(n6_adj_5655), .O(n60664));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1628 (.I0(n26315), .I1(n27223), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_adj_5621));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1628.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1629 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26294));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1629.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_772));   // verilog/coms.v(81[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(\data_in_frame[1] [4]), .I1(Kp_23__N_772), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[1] [3]), .O(n66276));
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1631 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26284));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1631.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1632 (.I0(\data_in_frame[1][0] ), .I1(Kp_23__N_767), 
            .I2(GND_net), .I3(GND_net), .O(n26266));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1632.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1633 (.I0(\data_in_frame[0][6] ), .I1(\data_in_frame[3] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n66420));
    defparam i1_2_lut_adj_1633.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1634 (.I0(\data_in_frame[5] [0]), .I1(Kp_23__N_799), 
            .I2(GND_net), .I3(GND_net), .O(n26716));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1634.LUT_INIT = 16'h6666;
    SB_LUT4 i60968_4_lut (.I0(n78636), .I1(n78840), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n76803));
    defparam i60968_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i55771_3_lut (.I0(n78540), .I1(n76803), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i55771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(n66420), .I1(n26266), .I2(\data_in_frame[5] [2]), 
            .I3(\data_in_frame[5] [3]), .O(n66397));
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1636 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n26297));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1637 (.I0(n26297), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n66175));
    defparam i1_2_lut_adj_1637.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1638 (.I0(\data_in_frame[0][0] ), .I1(\data_in_frame[2][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n66286));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1638.LUT_INIT = 16'h6666;
    SB_LUT4 i15625_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29837));
    defparam i15625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n66657));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'h6666;
    SB_LUT4 i15622_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29834));
    defparam i15622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1640 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [1]), 
            .I2(\data_in_frame[4] [7]), .I3(GND_net), .O(n66404));   // verilog/coms.v(88[17:70])
    defparam i1_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1641 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n66318));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1641.LUT_INIT = 16'h6666;
    SB_LUT4 i15619_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29831));
    defparam i15619_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[3] [5]), .O(n71027));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'h6996;
    SB_LUT4 i15616_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29828));
    defparam i15616_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[2][4] ), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[4] [0]), .O(n71025));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1644 (.I0(\data_in_frame[2]_c [2]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [6]), .I3(GND_net), .O(n71023));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_adj_1644.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1645 (.I0(n66404), .I1(n71025), .I2(n71027), 
            .I3(GND_net), .O(n71037));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_adj_1645.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n71023), .I1(Kp_23__N_753), .I2(\data_in_frame[2][0] ), 
            .I3(\data_in_frame[2][6] ), .O(n71035));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i15613_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29825));
    defparam i15613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n71035), .I1(n71037), .I2(n66657), 
            .I3(n66286), .O(n71041));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n66175), .I1(n26722), .I2(n71041), 
            .I3(n26188), .O(n71049));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1649 (.I0(n71049), .I1(n26137), .I2(n66264), 
            .I3(GND_net), .O(n71051));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_adj_1649.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n26583), .I1(n66397), .I2(n26716), 
            .I3(n71051), .O(n61328));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 i15610_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29822));
    defparam i15610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(\data_in_frame[6] [4]), .I1(n26294), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[6] [1]), .O(n66365));   // verilog/coms.v(88[17:28])
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1652 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n66254));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1652.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1653 (.I0(n66365), .I1(n61328), .I2(n26722), 
            .I3(n66318), .O(n15_adj_5656));
    defparam i6_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i15607_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29819));
    defparam i15607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1654 (.I0(n15_adj_5656), .I1(n70901), .I2(n14_adj_5627), 
            .I3(\data_in_frame[3] [6]), .O(n69110));
    defparam i8_4_lut_adj_1654.LUT_INIT = 16'h6996;
    SB_LUT4 i4_3_lut (.I0(n26673), .I1(n69075), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n21_adj_5657));
    defparam i4_3_lut.LUT_INIT = 16'h4141;
    SB_LUT4 i10_4_lut_adj_1655 (.I0(n69189), .I1(n24268), .I2(n24272), 
            .I3(n69110), .O(n27_adj_5658));
    defparam i10_4_lut_adj_1655.LUT_INIT = 16'h0040;
    SB_LUT4 i9_3_lut (.I0(n4_adj_5621), .I1(n60664), .I2(n61449), .I3(GND_net), 
            .O(n26_adj_5659));
    defparam i9_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i55542_2_lut (.I0(n26846), .I1(n26329), .I2(GND_net), .I3(GND_net), 
            .O(n71362));
    defparam i55542_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i55660_4_lut (.I0(n7_adj_5653), .I1(n26685), .I2(n26816), 
            .I3(n60607), .O(n71486));
    defparam i55660_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15604_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66099), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29816));
    defparam i15604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1656 (.I0(n27_adj_5658), .I1(n21_adj_5657), .I2(n26244), 
            .I3(n7_adj_15), .O(n31_adj_5660));
    defparam i14_4_lut_adj_1656.LUT_INIT = 16'h0008;
    SB_LUT4 i16_4_lut_adj_1657 (.I0(n31_adj_5660), .I1(n71486), .I2(n71362), 
            .I3(n26_adj_5659), .O(LED_N_3408));
    defparam i16_4_lut_adj_1657.LUT_INIT = 16'h0200;
    SB_LUT4 i5_4_lut_adj_1658 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[22] [1]), .I3(\data_in_frame[21] [7]), .O(n12_adj_5661));
    defparam i5_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1659 (.I0(\data_in_frame[21] [3]), .I1(n66558), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5662));
    defparam i1_2_lut_adj_1659.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1660 (.I0(\data_in_frame[20][3] ), .I1(\data_in_frame[18] [2]), 
            .I2(n66584), .I3(GND_net), .O(n8_adj_5663));
    defparam i3_3_lut_adj_1660.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1661 (.I0(\data_in_frame[20][4] ), .I1(n66574), 
            .I2(n60628), .I3(\data_in_frame[22] [6]), .O(n68484));
    defparam i3_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n60723), .I1(n68484), .I2(n8_adj_5663), 
            .I3(\data_in_frame[22] [4]), .O(n70941));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1663 (.I0(\data_in_frame[22] [5]), .I1(n66429), 
            .I2(GND_net), .I3(GND_net), .O(n66430));
    defparam i1_2_lut_adj_1663.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62770 (.I0(byte_transmit_counter[1]), 
            .I1(n71916), .I2(n71917), .I3(byte_transmit_counter[2]), .O(n78621));
    defparam byte_transmit_counter_1__bdd_4_lut_62770.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1664 (.I0(\data_in_frame[23] [4]), .I1(\data_in_frame[21] [2]), 
            .I2(n66193), .I3(n6_adj_5662), .O(n68439));
    defparam i4_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1665 (.I0(\data_in_frame[20][0] ), .I1(n12_adj_5661), 
            .I2(n66488), .I3(\data_in_frame[19] [5]), .O(n68725));
    defparam i6_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i6772_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1949), 
            .I2(n68081), .I3(n4452), .O(n20632));   // verilog/coms.v(148[4] 304[11])
    defparam i6772_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i3_4_lut_adj_1666 (.I0(n68427), .I1(n68131), .I2(\data_in_frame[21] [7]), 
            .I3(\data_in_frame[21] [6]), .O(n8_adj_5664));
    defparam i3_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(n68725), .I1(n68439), .I2(n66430), 
            .I3(n70941), .O(n70947));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'h0800;
    SB_LUT4 i2_3_lut_adj_1668 (.I0(n26522), .I1(\data_in_frame[21] [4]), 
            .I2(\data_in_frame[21] [3]), .I3(GND_net), .O(n66261));
    defparam i2_3_lut_adj_1668.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(\data_in_frame[22] [0]), .I1(n70947), 
            .I2(n8_adj_5664), .I3(\data_in_frame[19] [6]), .O(n70949));
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_adj_1670 (.I0(n68427), .I1(\data_in_frame[21] [4]), 
            .I2(n66558), .I3(GND_net), .O(n6_adj_5665));
    defparam i2_3_lut_adj_1670.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(\data_in_frame[23] [5]), .I1(n70949), 
            .I2(n66261), .I3(n68895), .O(n70951));
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'h4884;
    SB_LUT4 i1_4_lut_adj_1672 (.I0(n20632), .I1(n1949), .I2(n23015), .I3(n4), 
            .O(n27430));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1672.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_3_lut_adj_1673 (.I0(\data_in_frame[21] [2]), .I1(\data_in_frame[23] [3]), 
            .I2(\data_in_frame[21] [1]), .I3(GND_net), .O(n71153));
    defparam i1_3_lut_adj_1673.LUT_INIT = 16'h9696;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2058));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n26522), .I1(Kp_23__N_1607), .I2(n71153), 
            .I3(n66193), .O(n68677));
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(n66538), .I1(n60628), .I2(\data_in_frame[17] [6]), 
            .I3(\data_in_frame[22] [2]), .O(n71149));
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n66584), .I1(n66497), .I2(\data_in_frame[20][1] ), 
            .I3(\data_in_frame[22] [3]), .O(n71123));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1677 (.I0(\data_in_frame[21] [6]), .I1(n66336), 
            .I2(n68895), .I3(\data_in_frame[23] [7]), .O(n67899));
    defparam i3_4_lut_adj_1677.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(\data_in_frame[23] [6]), .I1(n70951), 
            .I2(n6_adj_5665), .I3(\data_in_frame[21] [5]), .O(n70953));
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'h4884;
    SB_LUT4 i1_3_lut_adj_1679 (.I0(n66384), .I1(Kp_23__N_1607), .I2(\data_in_frame[23] [1]), 
            .I3(GND_net), .O(n68042));
    defparam i1_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n71149), .I1(n68677), .I2(n66713), 
            .I3(n61678), .O(n70959));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'h4884;
    SB_LUT4 n78621_bdd_4_lut (.I0(n78621), .I1(n71914), .I2(n71913), .I3(byte_transmit_counter[2]), 
            .O(n78624));
    defparam n78621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n70959), .I1(n68042), .I2(n70953), 
            .I3(n67899), .O(n70961));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'h0080;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(\data_in_frame[19] [7]), .I1(n66713), 
            .I2(n71123), .I3(n60628), .O(n68851));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1683 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n71127));
    defparam i1_2_lut_adj_1683.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n71127), .I1(n68851), .I2(n70961), 
            .I3(n68740), .O(n70965));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'h2010;
    SB_LUT4 i55491_4_lut (.I0(n1949), .I1(n1952), .I2(n3303), .I3(n1955), 
            .O(n71310));   // verilog/coms.v(139[4] 141[7])
    defparam i55491_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n66833), .I1(n68740), .I2(n70933), 
            .I3(n66384), .O(n68441));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1686 (.I0(\data_in_frame[23] [0]), .I1(n68740), 
            .I2(n66384), .I3(GND_net), .O(n66732));
    defparam i1_3_lut_adj_1686.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n69189), .I1(n66732), .I2(n68441), 
            .I3(n70965), .O(Kp_23__N_612));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1952), 
            .I2(n71310), .I3(n67901), .O(n65018));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'hb3a0;
    SB_LUT4 i6777_4_lut (.I0(n1953), .I1(\FRAME_MATCHER.state[3] ), .I2(n1955), 
            .I3(n25857), .O(n20637));   // verilog/coms.v(148[4] 304[11])
    defparam i6777_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2047));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2046));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16158_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[7]), 
            .I3(\data_in_frame[13][7] ), .O(n30370));
    defparam i16158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1689 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n66491));
    defparam i1_2_lut_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1690 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n6_adj_5564));
    defparam i1_2_lut_3_lut_adj_1690.LUT_INIT = 16'h9696;
    SB_LUT4 i16154_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[6]), 
            .I3(\data_in_frame[13][6] ), .O(n30366));
    defparam i16154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16151_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n30363));
    defparam i16151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16148_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[4]), 
            .I3(\data_in_frame[13]_c [4]), .O(n30360));
    defparam i16148_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16145_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n30357));
    defparam i16145_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16141_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n30353));
    defparam i16141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n78849_bdd_4_lut (.I0(n78849), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n78852));
    defparam n78849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30605_4_lut (.I0(n5_adj_5385), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i30605_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i16138_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n30350));
    defparam i16138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16135_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66103), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n30347));
    defparam i16135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1691 (.I0(\FRAME_MATCHER.i[4] ), .I1(n25877), .I2(GND_net), 
            .I3(GND_net), .O(n25747));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1691.LUT_INIT = 16'heeee;
    SB_LUT4 i30609_4_lut (.I0(n8_adj_9), .I1(\FRAME_MATCHER.i [31]), .I2(n25747), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i30609_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut_adj_1692 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n23015));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1692.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1693 (.I0(Kp_23__N_612), .I1(Kp_23__N_1748), .I2(GND_net), 
            .I3(GND_net), .O(n28088));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'h8888;
    SB_LUT4 i61893_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_612), 
            .I2(LED_N_3408), .I3(Kp_23__N_1748), .O(n28129));
    defparam i61893_4_lut.LUT_INIT = 16'hc4a0;
    SB_LUT4 i3_2_lut (.I0(n25857), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27992));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1694 (.I0(n4452), .I1(n27992), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n23015), .O(n68490));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1694.LUT_INIT = 16'hffdc;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62756 (.I0(byte_transmit_counter[1]), 
            .I1(n71775), .I2(n71776), .I3(byte_transmit_counter[2]), .O(n78603));
    defparam byte_transmit_counter_1__bdd_4_lut_62756.LUT_INIT = 16'he4aa;
    SB_LUT4 n78603_bdd_4_lut (.I0(n78603), .I1(n71875), .I2(n71874), .I3(byte_transmit_counter[2]), 
            .O(n78606));
    defparam n78603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i58932_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74435));   // verilog/coms.v(158[12:15])
    defparam i58932_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n25866), .I1(n1955), .I2(n1953), .I3(n68490), 
            .O(n27427));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hbaaa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62746 (.I0(byte_transmit_counter[1]), 
            .I1(n71856), .I2(n71857), .I3(byte_transmit_counter[2]), .O(n78597));
    defparam byte_transmit_counter_1__bdd_4_lut_62746.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_adj_1696 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5666));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_adj_1696.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1697 (.I0(\data_in[1] [7]), .I1(\data_in[3] [4]), 
            .I2(\data_in[0] [0]), .I3(\data_in[1] [1]), .O(n68362));
    defparam i3_4_lut_adj_1697.LUT_INIT = 16'hfff7;
    SB_LUT4 i6_4_lut_adj_1698 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n14_adj_5667));   // verilog/coms.v(157[7:23])
    defparam i6_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1699 (.I0(\FRAME_MATCHER.i [15]), .I1(n14_adj_5667), 
            .I2(n10_adj_5666), .I3(\FRAME_MATCHER.i [22]), .O(n68038));   // verilog/coms.v(157[7:23])
    defparam i7_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1700 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(\FRAME_MATCHER.i [19]), .O(n14_adj_5668));   // verilog/coms.v(157[7:23])
    defparam i6_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1701 (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [23]), .O(n13_adj_5669));   // verilog/coms.v(157[7:23])
    defparam i5_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1702 (.I0(\FRAME_MATCHER.i [20]), .I1(n68038), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [11]), .O(n20_adj_5670));   // verilog/coms.v(157[7:23])
    defparam i8_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1703 (.I0(\FRAME_MATCHER.i [13]), .I1(n13_adj_5669), 
            .I2(n14_adj_5668), .I3(GND_net), .O(n13_adj_5671));   // verilog/coms.v(157[7:23])
    defparam i1_3_lut_adj_1703.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5672));   // verilog/coms.v(157[7:23])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1704 (.I0(n13_adj_5671), .I1(n20_adj_5670), .I2(\FRAME_MATCHER.i [28]), 
            .I3(\FRAME_MATCHER.i [16]), .O(n22_adj_5673));   // verilog/coms.v(157[7:23])
    defparam i10_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1705 (.I0(\data_in[2] [7]), .I1(\data_in[0] [4]), 
            .I2(n68362), .I3(GND_net), .O(n25913));
    defparam i2_3_lut_adj_1705.LUT_INIT = 16'hf7f7;
    SB_LUT4 i16184_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[7]), 
            .I3(\data_in_frame[14][7] ), .O(n30396));
    defparam i16184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1706 (.I0(\FRAME_MATCHER.i [7]), .I1(n22_adj_5673), 
            .I2(n18_adj_5672), .I3(\FRAME_MATCHER.i [12]), .O(n25877));   // verilog/coms.v(157[7:23])
    defparam i11_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i30610_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25877), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i30610_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i6_4_lut_adj_1707 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5674));
    defparam i6_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i16181_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[6]), 
            .I3(\data_in_frame[14][6] ), .O(n30393));
    defparam i16181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16178_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[5]), 
            .I3(\data_in_frame[14][5] ), .O(n30390));
    defparam i16178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2066));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1708 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5675));
    defparam i7_4_lut_adj_1708.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_4_lut_adj_1709 (.I0(n61607), .I1(n10_adj_5513), .I2(\data_out_frame[18] [2]), 
            .I3(\data_out_frame[20] [4]), .O(n60687));
    defparam i1_2_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 i16174_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[4]), 
            .I3(\data_in_frame[14][4] ), .O(n30386));
    defparam i16174_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1710 (.I0(n61607), .I1(n10_adj_5513), .I2(\data_out_frame[18] [2]), 
            .I3(n68344), .O(n66745));
    defparam i1_2_lut_4_lut_adj_1710.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1711 (.I0(n17_adj_5675), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5674), .I3(\data_in[2] [6]), .O(n25954));
    defparam i9_4_lut_adj_1711.LUT_INIT = 16'hfbff;
    SB_LUT4 i16171_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[3]), 
            .I3(\data_in_frame[14]_c [3]), .O(n30383));
    defparam i16171_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15934_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n30146));
    defparam i15934_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15937_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n30149));
    defparam i15937_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15940_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n30152));
    defparam i15940_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1712 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5676));
    defparam i2_2_lut_adj_1712.LUT_INIT = 16'heeee;
    SB_LUT4 i15943_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n30155));
    defparam i15943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n78597_bdd_4_lut (.I0(n78597), .I1(n71848), .I2(n71847), .I3(byte_transmit_counter[2]), 
            .O(n78600));
    defparam n78597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15946_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n30158));
    defparam i15946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15949_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n30161));
    defparam i15949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i58948_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74439));   // verilog/coms.v(158[12:15])
    defparam i58948_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1713 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5677));
    defparam i6_4_lut_adj_1713.LUT_INIT = 16'hfeff;
    SB_LUT4 i15952_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n30164));
    defparam i15952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1714 (.I0(\data_in[3] [6]), .I1(n14_adj_5677), 
            .I2(n10_adj_5676), .I3(\data_in[2] [1]), .O(n25907));
    defparam i7_4_lut_adj_1714.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1715 (.I0(n25907), .I1(\data_in[2] [0]), .I2(\data_in[2] [6]), 
            .I3(\data_in[0] [5]), .O(n20_adj_5678));
    defparam i8_4_lut_adj_1715.LUT_INIT = 16'hfbff;
    SB_LUT4 i16168_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n30380));
    defparam i16168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16164_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n30376));
    defparam i16164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15955_3_lut_4_lut (.I0(n8_adj_5632), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n30167));
    defparam i15955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1716 (.I0(n25777), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_adj_5679));
    defparam i7_4_lut_adj_1716.LUT_INIT = 16'hfeff;
    SB_LUT4 i16161_3_lut_4_lut (.I0(n8_adj_5610), .I1(n66103), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n30373));
    defparam i16161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i55664_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[3] [2]), .I2(\data_in[1] [3]), 
            .I3(\data_in[1] [2]), .O(n71490));
    defparam i55664_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62741 (.I0(byte_transmit_counter[1]), 
            .I1(n71835), .I2(n71836), .I3(byte_transmit_counter[2]), .O(n78591));
    defparam byte_transmit_counter_1__bdd_4_lut_62741.LUT_INIT = 16'he4aa;
    SB_LUT4 equal_308_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5632));   // verilog/coms.v(157[7:23])
    defparam equal_308_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i11_3_lut_adj_1717 (.I0(n71490), .I1(n19_adj_5679), .I2(n20_adj_5678), 
            .I3(GND_net), .O(n1949));
    defparam i11_3_lut_adj_1717.LUT_INIT = 16'hfdfd;
    SB_LUT4 n78591_bdd_4_lut (.I0(n78591), .I1(n71827), .I2(n71826), .I3(byte_transmit_counter[2]), 
            .O(n78594));
    defparam n78591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1718 (.I0(\data_out_frame[20] [2]), .I1(n61643), 
            .I2(\data_out_frame[22] [3]), .I3(n66562), .O(n25456));
    defparam i2_3_lut_4_lut_adj_1718.LUT_INIT = 16'h9669;
    SB_LUT4 i55567_2_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n71389));
    defparam i55567_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1719 (.I0(\data_in[3] [0]), .I1(\data_in[1] [5]), 
            .I2(n25913), .I3(n25907), .O(n18_adj_5680));
    defparam i7_4_lut_adj_1719.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1720 (.I0(n25954), .I1(\data_in[0] [3]), .I2(\data_in[1] [0]), 
            .I3(\data_in[2] [2]), .O(n19_adj_5681));
    defparam i8_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1721 (.I0(n19_adj_5681), .I1(\data_in[0] [6]), 
            .I2(n18_adj_5680), .I3(n71389), .O(n1952));
    defparam i10_4_lut_adj_1721.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_1722 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5682));
    defparam i5_3_lut_adj_1722.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1723 (.I0(\data_in[0] [6]), .I1(n25913), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5683));
    defparam i6_4_lut_adj_1723.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1724 (.I0(n15_adj_5683), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5682), .I3(\data_in[0] [3]), .O(n25777));
    defparam i8_4_lut_adj_1724.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_4_lut_adj_1725 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n10_adj_5507), .I3(n61760), .O(n66562));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_4_lut_adj_1725.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1726 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n25777), .O(n16_adj_5684));
    defparam i6_4_lut_adj_1726.LUT_INIT = 16'hffef;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n66704), .I3(\data_out_frame[19] [5]), .O(n20_adj_5479));   // verilog/coms.v(74[16:27])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1727 (.I0(n25954), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5685));
    defparam i7_4_lut_adj_1727.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1728 (.I0(n17_adj_5685), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5684), .I3(\data_in[3] [3]), .O(n1955));
    defparam i9_4_lut_adj_1728.LUT_INIT = 16'hfbff;
    SB_LUT4 i366_2_lut (.I0(n1952), .I1(n1949), .I2(GND_net), .I3(GND_net), 
            .O(n1953));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1729 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(GND_net), .I3(GND_net), .O(n66134));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1730 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5686));   // verilog/coms.v(217[11:56])
    defparam i1_2_lut_adj_1730.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5687));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'ha8a0;
    SB_LUT4 i31193_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5687), .I3(n4_adj_5686), .O(n45273));
    defparam i31193_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i2_4_lut_adj_1732 (.I0(n66134), .I1(n1953), .I2(n1955), .I3(\FRAME_MATCHER.i_31__N_2507 ), 
            .O(n6_adj_5688));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1732.LUT_INIT = 16'heaaa;
    SB_LUT4 i14495_3_lut_4_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n82), .I2(n66108), 
            .I3(reset), .O(n66998));   // verilog/coms.v(156[9:50])
    defparam i14495_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1733 (.I0(\FRAME_MATCHER.i[5] ), .I1(n82), 
            .I2(n3474), .I3(GND_net), .O(n41543));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_adj_1733.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_4_lut_adj_1734 (.I0(\data_out_frame[20] [4]), .I1(n66248), 
            .I2(\data_out_frame[20] [5]), .I3(n66435), .O(n68344));
    defparam i2_3_lut_4_lut_adj_1734.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1735 (.I0(n68152), .I1(n6_adj_5688), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n79076));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1735.LUT_INIT = 16'hefee;
    SB_LUT4 i16211_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n30423));
    defparam i16211_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1736 (.I0(\data_out_frame[20] [4]), .I1(n66248), 
            .I2(\data_out_frame[22] [7]), .I3(n68344), .O(n66413));
    defparam i2_3_lut_4_lut_adj_1736.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1737 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n66248));
    defparam i1_2_lut_3_lut_adj_1737.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1738 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(n68217), .I3(n61306), .O(n24043));
    defparam i2_3_lut_4_lut_adj_1738.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1739 (.I0(\data_out_frame[23] [5]), .I1(n66616), 
            .I2(n61583), .I3(\data_out_frame[24] [0]), .O(n66824));
    defparam i2_3_lut_4_lut_adj_1739.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1740 (.I0(\data_out_frame[23] [5]), .I1(n66616), 
            .I2(\data_out_frame[23] [3]), .I3(n26898), .O(n66444));
    defparam i1_2_lut_3_lut_4_lut_adj_1740.LUT_INIT = 16'h6996;
    SB_LUT4 i16208_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n30420));
    defparam i16208_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16204_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n30416));
    defparam i16204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i23_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(\data_in_frame[15] [4]), 
            .I3(rx_data[4]), .O(n15));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16198_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n30410));
    defparam i16198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [3]), 
            .I2(encoder0_position[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62736 (.I0(byte_transmit_counter[1]), 
            .I1(n71898), .I2(n71899), .I3(byte_transmit_counter[2]), .O(n78585));
    defparam byte_transmit_counter_1__bdd_4_lut_62736.LUT_INIT = 16'he4aa;
    SB_LUT4 i16194_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n30406));
    defparam i16194_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15549_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29761));
    defparam i15549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16191_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n30403));
    defparam i16191_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i58925_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74440));   // verilog/coms.v(158[12:15])
    defparam i58925_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15545_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29757));
    defparam i15545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16188_3_lut_4_lut (.I0(n45146), .I1(n66103), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n30400));
    defparam i16188_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15542_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29754));
    defparam i15542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15538_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29750));
    defparam i15538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15535_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29747));
    defparam i15535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15532_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29744));
    defparam i15532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15529_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29741));
    defparam i15529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15526_3_lut_4_lut (.I0(n8_adj_5608), .I1(n66099), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29738));
    defparam i15526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n78585_bdd_4_lut (.I0(n78585), .I1(n71830), .I2(n71829), .I3(byte_transmit_counter[2]), 
            .O(n78588));
    defparam n78585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62948 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n78837));
    defparam byte_transmit_counter_0__bdd_4_lut_62948.LUT_INIT = 16'he4aa;
    SB_LUT4 n78837_bdd_4_lut (.I0(n78837), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n78840));
    defparam n78837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15717_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[2][6] ), .O(n29929));
    defparam i15717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15714_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[2]_c [5]), .O(n29926));
    defparam i15714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15711_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[2][4] ), .O(n29923));
    defparam i15711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5558));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5557));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5556));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62938 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n78831));
    defparam byte_transmit_counter_0__bdd_4_lut_62938.LUT_INIT = 16'he4aa;
    SB_LUT4 select_789_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5555));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i15708_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[2][3] ), .O(n29920));
    defparam i15708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15705_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[2]_c [2]), .O(n29917));
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5554));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5551));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i15702_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[1]), 
            .I3(\data_in_frame[2][1] ), .O(n29914));
    defparam i15702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_adj_5550));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1742 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n66131));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i15697_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[0]), 
            .I3(\data_in_frame[2][0] ), .O(n29909));
    defparam i15697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_789_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5549));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 n78831_bdd_4_lut (.I0(n78831), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n78834));
    defparam n78831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15739_3_lut_4_lut (.I0(n8_adj_13), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29951));
    defparam i15739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[23] [3]), .I3(n26898), .O(n6_c));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_4_lut_adj_1743 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n61587), .I3(n10_adj_5384), .O(n26526));
    defparam i5_3_lut_4_lut_adj_1743.LUT_INIT = 16'h6996;
    SB_LUT4 equal_311_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_13));   // verilog/coms.v(157[7:23])
    defparam equal_311_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62780 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(byte_transmit_counter[1]), .O(n78561));
    defparam byte_transmit_counter_0__bdd_4_lut_62780.LUT_INIT = 16'he4aa;
    SB_LUT4 n78561_bdd_4_lut (.I0(n78561), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(byte_transmit_counter[1]), 
            .O(n78564));
    defparam n78561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59191_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74446));   // verilog/coms.v(158[12:15])
    defparam i59191_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i58982_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74447));   // verilog/coms.v(158[12:15])
    defparam i58982_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 equal_310_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5608));   // verilog/coms.v(157[7:23])
    defparam equal_310_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62933 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n78825));
    defparam byte_transmit_counter_0__bdd_4_lut_62933.LUT_INIT = 16'he4aa;
    SB_LUT4 i58983_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74448));   // verilog/coms.v(158[12:15])
    defparam i58983_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i59039_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74463));   // verilog/coms.v(158[12:15])
    defparam i59039_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i59093_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74465));   // verilog/coms.v(158[12:15])
    defparam i59093_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n78825_bdd_4_lut (.I0(n78825), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n78828));
    defparam n78825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i59029_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74467));   // verilog/coms.v(158[12:15])
    defparam i59029_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i59028_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74468));   // verilog/coms.v(158[12:15])
    defparam i59028_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i19852_3_lut_4_lut (.I0(deadband[19]), .I1(\data_in_frame[14]_c [3]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30075));
    defparam i19852_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62928 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n78819));
    defparam byte_transmit_counter_0__bdd_4_lut_62928.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_62731 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[21] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[0]), .O(n78543));
    defparam byte_transmit_counter_1__bdd_4_lut_62731.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5488));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n78543_bdd_4_lut (.I0(n78543), .I1(\data_out_frame[22] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(byte_transmit_counter[0]), 
            .O(n78546));
    defparam n78543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [1]), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_62722 (.I0(byte_transmit_counter[2]), 
            .I1(n71867), .I2(n71834), .I3(byte_transmit_counter[3]), .O(n78537));
    defparam byte_transmit_counter_2__bdd_4_lut_62722.LUT_INIT = 16'he4aa;
    SB_LUT4 n78537_bdd_4_lut (.I0(n78537), .I1(n71761), .I2(n71760), .I3(byte_transmit_counter[3]), 
            .O(n78540));
    defparam n78537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62712 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n78525));
    defparam byte_transmit_counter_0__bdd_4_lut_62712.LUT_INIT = 16'he4aa;
    SB_LUT4 n78525_bdd_4_lut (.I0(n78525), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n78528));
    defparam n78525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n78819_bdd_4_lut (.I0(n78819), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n78822));
    defparam n78819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62685 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n78501));
    defparam byte_transmit_counter_0__bdd_4_lut_62685.LUT_INIT = 16'he4aa;
    SB_LUT4 n78501_bdd_4_lut (.I0(n78501), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n78504));
    defparam n78501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15693_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29905));
    defparam i15693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i59008_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74469));   // verilog/coms.v(158[12:15])
    defparam i59008_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i19656_3_lut_4_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13]_c [4]), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30067));
    defparam i19656_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15689_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[6]), 
            .I3(\data_in_frame[1][6] ), .O(n29901));
    defparam i15689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i59788_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n74486));   // verilog/coms.v(158[12:15])
    defparam i59788_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14438_1_lut (.I0(n3474), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28649));   // verilog/coms.v(148[4] 304[11])
    defparam i14438_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_62665 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n78495));
    defparam byte_transmit_counter_0__bdd_4_lut_62665.LUT_INIT = 16'he4aa;
    SB_LUT4 i15686_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29898));
    defparam i15686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n78495_bdd_4_lut (.I0(n78495), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n78498));
    defparam n78495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5486));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15683_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29895));
    defparam i15683_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15680_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29892));
    defparam i15680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1745 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[3][7] ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5485));
    defparam i1_3_lut_adj_1745.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_3_lut_adj_1746 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[3][6] ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5484));
    defparam i1_3_lut_adj_1746.LUT_INIT = 16'ha8a8;
    SB_LUT4 select_787_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15677_3_lut_4_lut (.I0(n8), .I1(n66156), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29889));
    defparam i15677_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.clk16MHz(clk16MHz), .tx_o(tx_o), .tx_data({tx_data[7:4], 
            \tx_data[3] , tx_data[2:0]}), .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), 
            .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), .GND_net(GND_net), 
            .n29954(n29954), .tx_active(tx_active), .r_Clock_Count({r_Clock_Count}), 
            .VCC_net(VCC_net), .n67642(n67642), .n6(n6_adj_16), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29(n29), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n23(n23), .n5218(n5218), .n67002(n67002), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.baudrate({baudrate}), .GND_net(GND_net), .n28238(n28238), 
            .clk16MHz(clk16MHz), .n67079(n67079), .\r_SM_Main[2] (\r_SM_Main[2]_adj_17 ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .n33(n33), .n34(n34_adj_18), 
            .n29935(n29935), .rx_data({rx_data}), .n29934(n29934), .n29932(n29932), 
            .n29913(n29913), .n29912(n29912), .n29908(n29908), .n29904(n29904), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n5215(n5215), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n29(n29), .n23(n23), .\r_SM_Main[1] (\r_SM_Main[1]_adj_19 ), 
            .n27(n27), .n28115(n28115), .r_Clock_Count({r_Clock_Count_adj_28}), 
            .VCC_net(VCC_net), .n30760(n30760), .n61786(n61786), .rx_data_ready(rx_data_ready), 
            .n30756(n30756), .\r_Bit_Index[0] (\r_Bit_Index[0] ), .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), 
            .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), 
            .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n69006(n69006), .n69649(n69649), .n69585(n69585), .n69665(n69665), 
            .n69633(n69633), .n69601(n69601), .n69617(n69617), .n69697(n69697), 
            .n69681(n69681), .n69523(n69523)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk16MHz, tx_o, tx_data, r_SM_Main, \r_SM_Main_2__N_3536[1] , 
            \r_SM_Main_2__N_3545[0] , GND_net, n29954, tx_active, r_Clock_Count, 
            VCC_net, n67642, n6, \o_Rx_DV_N_3488[24] , n27, n29, 
            \o_Rx_DV_N_3488[12] , n23, n5218, n67002, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output tx_o;
    input [7:0]tx_data;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    input \r_SM_Main_2__N_3545[0] ;
    input GND_net;
    input n29954;
    output tx_active;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n67642;
    output n6;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    input n29;
    input \o_Rx_DV_N_3488[12] ;
    input n23;
    input n5218;
    input n67002;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n460;
    
    wire n67121;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n29496, n3, n40335, n25368;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n61818, n71922, n71923, n71614, n71613, n79052, n74485, 
        n67613, n61816;
    wire [8:0]n41;
    
    wire n40307, n3_adj_5307, n59588, n59587, n59586, n59585, n59584, 
        n59583, n59582, n59581, n14, n15, n69541, n69547, n66052, 
        n74474, n74471, n9, n78558, n78555;
    
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n67121), 
            .D(n460[1]), .R(n29496));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n67121), 
            .D(n460[2]), .R(n29496));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40335), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n61818), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i62630_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n67121));
    defparam i62630_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n25368));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i56087_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n71922));
    defparam i56087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i56088_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n71923));
    defparam i56088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55779_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n71614));
    defparam i55779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i55778_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n71613));
    defparam i55778_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n79052));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29954));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i12_4_lut (.I0(n74485), .I1(n67121), .I2(r_Bit_Index[0]), 
            .I3(n67613), .O(n61816));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_DFFESR r_Clock_Count_2056__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40335), .D(n41[0]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40335), .D(n41[1]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40335), .D(n41[2]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40335), .D(n41[3]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40335), .D(n41[4]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40335), .D(n41[5]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40335), .D(n41[6]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40335), .D(n41[7]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40335), .D(n41[8]), .R(n40307));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n61816));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5307), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25368), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_2056_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n59588), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2056_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n59587), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_9 (.CI(n59587), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n59588));
    SB_LUT4 r_Clock_Count_2056_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n59586), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_8 (.CI(n59586), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n59587));
    SB_LUT4 r_Clock_Count_2056_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n59585), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_7 (.CI(n59585), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n59586));
    SB_LUT4 r_Clock_Count_2056_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n59584), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_6 (.CI(n59584), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n59585));
    SB_LUT4 r_Clock_Count_2056_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n59583), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_5 (.CI(n59583), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n59584));
    SB_LUT4 r_Clock_Count_2056_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n59582), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_4 (.CI(n59582), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n59583));
    SB_LUT4 r_Clock_Count_2056_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n59581), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_3 (.CI(n59581), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n59582));
    SB_LUT4 r_Clock_Count_2056_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n59581));
    SB_LUT4 i62484_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40307));
    defparam i62484_4_lut.LUT_INIT = 16'h1113;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n67642), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5218), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40335), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n79052));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i59786_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n74485));   // verilog/uart_tx.v(32[16:25])
    defparam i59786_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut (.I0(n5218), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n69541));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), .I3(n69541), 
            .O(n69547));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i10_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n69547), .O(n3_adj_5307));   // verilog/uart_tx.v(32[16:25])
    defparam i10_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i59747_3_lut (.I0(n66052), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5218), 
            .I3(GND_net), .O(n74474));   // verilog/uart_tx.v(32[16:25])
    defparam i59747_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i59744_4_lut (.I0(n74474), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n74471));   // verilog/uart_tx.v(32[16:25])
    defparam i59744_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i23_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n74471), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n61818));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40335));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n78558), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i26191_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i26191_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n66052));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i51108_rep_30_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n67613));
    defparam i51108_rep_30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1069 (.I0(n67002), .I1(n67613), .I2(r_SM_Main[1]), 
            .I3(n66052), .O(n29496));
    defparam i1_4_lut_adj_1069.LUT_INIT = 16'h1101;
    SB_LUT4 i16_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n71613), 
            .I2(n71614), .I3(r_Bit_Index[1]), .O(n78555));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n78555_bdd_4_lut (.I0(n78555), .I1(n71923), .I2(n71922), .I3(r_Bit_Index[1]), 
            .O(n78558));
    defparam n78555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (baudrate, GND_net, n28238, clk16MHz, n67079, \r_SM_Main[2] , 
            r_Rx_Data, RX_N_2, n33, n34, n29935, rx_data, n29934, 
            n29932, n29913, n29912, n29908, n29904, \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[12] , n5215, \o_Rx_DV_N_3488[24] , n29, 
            n23, \r_SM_Main[1] , n27, n28115, r_Clock_Count, VCC_net, 
            n30760, n61786, rx_data_ready, n30756, \r_Bit_Index[0] , 
            \r_SM_Main_2__N_3446[1] , \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            n69006, n69649, n69585, n69665, n69633, n69601, n69617, 
            n69697, n69681, n69523) /* synthesis syn_module_defined=1 */ ;
    input [31:0]baudrate;
    input GND_net;
    output n28238;
    input clk16MHz;
    output n67079;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input RX_N_2;
    output n33;
    output n34;
    input n29935;
    output [7:0]rx_data;
    input n29934;
    input n29932;
    input n29913;
    input n29912;
    input n29908;
    input n29904;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[12] ;
    input n5215;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output \r_SM_Main[1] ;
    output n27;
    output n28115;
    output [7:0]r_Clock_Count;
    input VCC_net;
    input n30760;
    input n61786;
    output rx_data_ready;
    input n30756;
    output \r_Bit_Index[0] ;
    input \r_SM_Main_2__N_3446[1] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n69006;
    output n69649;
    output n69585;
    output n69665;
    output n69633;
    output n69601;
    output n69617;
    output n69697;
    output n69681;
    input n69523;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n67224, n961, n42, n960, n77086, n959, n77087, n66912, 
        n48, n71570, n48_adj_5023, n962;
    wire [23:0]n294;
    
    wire n1115;
    wire [23:0]n8291;
    
    wire n1265, n1267, n36, n38, n41, n40, n74972, n77459, n1263, 
        n77460, n1262, n77288, n1261, n48_adj_5024;
    wire [23:0]n8317;
    
    wire n1414, n34_c, n41_adj_5025, n77078, n43, n77079, n39, 
        n74957, n75910, n36_adj_5026, n38_adj_5027, n45, n44, n76584, 
        n1408, n48_adj_5028, n69391, n1415;
    wire [23:0]n8343;
    
    wire n1559, n32, n39_adj_5029, n77076, n41_adj_5030, n77077, 
        n37, n74934, n75900, n34_adj_5031, n76586, n43_adj_5032, 
        n76949, n77074, n1553, n77075, n1552, n48_adj_5033, n25974, 
        n67167, n71554;
    wire [23:0]n8369;
    
    wire n1702;
    wire [23:0]n8395;
    
    wire n1840, n29_c, n35, n33_c, n31, n74859, n32_adj_5034, 
        n43_adj_5035, n40_adj_5036, n1841, n28, n77068, n37_adj_5037, 
        n77069, n41_adj_5038, n39_adj_5039, n74841, n30, n74834, 
        n77066, n76957, n77526, n1832, n77527, n1831, n48_adj_5040, 
        n1701, n1839;
    wire [23:0]n8421;
    
    wire n1974, n1975, n29_adj_5041, n31_adj_5042, n1973, n33_adj_5043, 
        n1976, n27_c, n74822, n71542, n67195, n30_adj_5044, n41_adj_5045, 
        n38_adj_5046, n26, n77235, n35_adj_5047, n77236, n39_adj_5048, 
        n37_adj_5049, n74815, n28_adj_5050, n74813, n77461, n76961, 
        n77625, n1968, n77626, n1967, n77604, n1966, n48_adj_5051;
    wire [23:0]n8447;
    
    wire n2108, n70773, n9, n14, n70643, n26008, n27_adj_5052, 
        n33_adj_5053, n31_adj_5054, n29_adj_5055, n74799, n30_adj_5056, 
        n41_adj_5057, n38_adj_5058, n67198, n2109, n26_adj_5059, n77062, 
        n35_adj_5060, n77063, n39_adj_5061, n37_adj_5062, n74795, 
        n28_adj_5063, n74790, n77463, n76967, n77627, n2100, n77628, 
        n2099, n77602, n2098, n48_adj_5064, n1977;
    wire [23:0]n8473;
    
    wire n2238, n2237, n25, n27_adj_5065, n2236, n29_adj_5066, n70817, 
        n70805, n71538, n71510, n71430, n2239, n23_c, n74758, 
        n35_adj_5067, n33_adj_5068, n31_adj_5069, n74754, n2240, n22, 
        n28_adj_5070, n30_adj_5071, n26_adj_5072, n37_adj_5073, n34_adj_5074, 
        n24, n74752, n77465, n39_adj_5075, n77466, n41_adj_5076, 
        n77278, n76872, n74756, n77052, n43_adj_5077, n42_adj_5078, 
        n77309, n2228, n77310, n2107;
    wire [23:0]n8499;
    
    wire n2362, n2234, n2360, n29_adj_5079, n2361, n31_adj_5080, 
        n33_adj_5081, n2366, n70793, n70769, n26014, n21, n27_adj_5082, 
        n25_adj_5083, n23_adj_5084, n74735, n74731, n2367, n20, 
        n26_adj_5085, n28_adj_5086, n24_adj_5087, n35_adj_5088, n32_adj_5089, 
        n22_adj_5090, n74729, n77467, n37_adj_5091, n77468, n39_adj_5092, 
        n77276, n76870, n74733, n77469, n41_adj_5093, n77244;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n77534, n2355, n77535, n2354, n77474, n2365;
    wire [23:0]n8525;
    
    wire n2488;
    wire [23:0]n8551;
    
    wire n2608, n23_adj_5094, n2607, n25_adj_5095, n2611, n17, n21_adj_5096, 
        n19, n75650, n29_adj_5097, n27_adj_5098, n75641, n35_adj_5099, 
        n33_adj_5100, n31_adj_5101, n77185, n2612, n16, n39_adj_5102, 
        n77014, n41_adj_5103, n77015, n75643, n76477, n22_adj_5104, 
        n76988, n43_adj_5105, n75941, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire r_Rx_Data_R, n20_adj_5106, n28_adj_5107, n18, n75639, n77261, 
        n77262, n77260, n37_adj_5108, n76479, n77010, n75939, n77543, 
        n2597, n77544, n2481, n2601;
    wire [23:0]n8577;
    
    wire n2718, n2609, n2726, n21_adj_5109, n2725, n23_adj_5110, 
        n2724, n25_adj_5111, n37_adj_5112, n69941, n70809, n70799, 
        n25965, n75539, n19_adj_5113, n17_adj_5114, n2729, n76465, 
        n76836, n31_adj_5115, n29_adj_5116, n27_adj_5117, n76834, 
        n35_adj_5118, n33_adj_5119, n75541, n2730, n14_adj_5120, n77004, 
        n39_adj_5121, n77005, n22_adj_5122, n45_adj_5123, n40_adj_5124, 
        n43_adj_5125, n41_adj_5126, n75534, n20_adj_5127, n75532, 
        n76990, n75951, n18_adj_5128, n26_adj_5129, n16_adj_5130, 
        n75575, n77263, n77264, n77256, n77179, n77430, n75949, 
        n77432;
    wire [23:0]n8603;
    
    wire n2839, n2727, n2841, n19_adj_5131, n2840, n21_adj_5132, 
        n23_adj_5133, n2833, n35_adj_5134, n70767, n70803, n25968, 
        n75491, n17_adj_5135, n15, n2844, n76423, n76818, n29_adj_5136, 
        n27_adj_5137, n25_adj_5138, n76816, n33_adj_5139, n31_adj_5140, 
        n75493, n2845, n12, n76964, n20_adj_5141, n43_adj_5142, 
        n38_adj_5143, n37_adj_5144, n76965, n41_adj_5145, n39_adj_5146, 
        n75481, n18_adj_5147, n75468, n77267, n75957, n16_adj_5148, 
        n24_adj_5149, n14_adj_5150, n75507, n77269, n77270, n77252, 
        n77171, n77599, n75955, n77633, n2828, n77634;
    wire [23:0]n8629;
    
    wire n2951, n2842, n2953, n17_adj_5151, n2952, n19_adj_5152, 
        n21_adj_5153, n70819, n70821, n25971, n33_adj_5154, n75434, 
        n15_adj_5155, n13, n2956, n76377, n76796, n1558, n27_adj_5156, 
        n25_adj_5157, n23_adj_5158, n76792, n31_adj_5159, n29_adj_5160, 
        n75436, n2957, n10, n76936, n35_adj_5161, n76937, n18_adj_5162, 
        n41_adj_5163, n36_adj_5164, n39_adj_5165, n37_adj_5166, n75425, 
        n16_adj_5167, n75419, n77291, n75963, n14_adj_5168, n22_adj_5169, 
        n12_adj_5170, n75448, n77289, n77290, n77232, n77161, n77524, 
        n75961, n77645, n2940, n77646, n2939, n77640, n2827, n2938;
    wire [23:0]n8655;
    
    wire n3046, n3186;
    wire [23:0]n8681;
    
    wire n3151, n26017, n67187, n67213, n71496, n76603, n66910, 
        n48_adj_5171, n25989, n74877, n44_adj_5172, n67171, n74573, 
        n71544, n71574, n45239, n69833, n48_adj_5173, n26020, n74882, 
        n805, n21177, n71578, n11690, n71498, n28_adj_5174, n2489, 
        n20_adj_5175, n2484, n74698, n22_adj_5176, n2486, n24_adj_5177, 
        n2487, n74703, n25935, n24_adj_5178, n22_adj_5179, n23_adj_5180;
    wire [23:0]n8707;
    
    wire n59407, n3152, n3082, n59406, n3153, n3188, n59405, n3154, 
        n3084, n59404, n69971, n3064, n10_adj_5181, n3061, n14_adj_5182, 
        n3051, n3060, n75356, n3155, n2977, n59403, n3156, n2867, 
        n59402, n3157, n2754, n59401, n16_adj_5183, n3059, n12_adj_5184, 
        n3158, n2638, n59400, n3159, n2519, n59399, n70801, n3160, 
        n2397, n59398, n3161, n2272, n59397, n3063, n75382, n70811, 
        n44716, n70745, n3162, n2144, n59396, n3163, n2013, n59395, 
        n66050, n74514, n74511, n79053;
    wire [7:0]n1;
    
    wire n28159, n29421, n3164, n1879, n59394, n3165, n1742, n59393, 
        n3166, n1602, n59392, n3167, n1459, n59391, n3168, n1460, 
        n59390, n3169, n1011, n59389, n3170, n856, n59388, n3171, 
        n698, n59387, n3172, n858, n59386, n69413, n538, n59385, 
        n67163, n59384, n3047, n59383, n3048, n59382, n3049, n59381, 
        n3050, n59380, n59379, n3052, n59378, n3053, n59377, n3054, 
        n59376, n3055, n59375, n3056, n59374, n3057, n59373, n3058, 
        n59372, n59371, n59370, n59369, n3062, n59368, n59367, 
        n59366, n3065, n59365, n3066, n59364, n69411, n59363, 
        n59362, n59361, n2941, n59360, n2942, n59359, n2943, n59358, 
        n2944, n59357, n2945, n59356, n2946, n59355, n25977, n2947, 
        n59354, n2948, n59353, n2949, n59352, n2950, n59351, n59350, 
        n59349, n41_adj_5198, n39_adj_5199, n37_adj_5200, n59348, 
        n23_adj_5201, n25_adj_5202, n2954, n59347, n29_adj_5203, n2955, 
        n59346, n31_adj_5204, n7, n59345, n45_adj_5205, n59344, 
        n43_adj_5206, n9_adj_5207, n17_adj_5208, n19_adj_5209, n69409, 
        n21_adj_5210, n35_adj_5211, n33_adj_5212, n11, n59343, n59342, 
        n13_adj_5213, n15_adj_5214, n27_adj_5215, n2829, n59341, n2830, 
        n59340, n75241, n2831, n59339, n2832, n59338, n12_adj_5216, 
        n75231, n10_adj_5217, n59337, n2834, n59336, n30_adj_5218, 
        n75259, n2835, n59335, n16_adj_5219, n2836, n59334, n75205, 
        n2837, n59333, n2838, n59332, n8, n24_adj_5220, n3274, 
        n59331, n75281, n76213, n76207, n77345, n59330, n76700, 
        n59329, n77491, n59328, n2843, n59327, n59326, n6, n76894, 
        n59325, n76895, n48_adj_5221, n4, n76892, n69407, n67175, 
        n76893, n2713, n59324, n2714, n59323, n75233, n2715, n59322, 
        n2716, n59321, n77375, n76001, n77585, n77586, n77513, 
        n75211, n2717, n59320, n77000, n59319, n75999, n75213, 
        n2719, n59318, n77433, n3_adj_5222, n76007, n3253, n77435, 
        n2720, n59317, n69339, n68384, n2721, n59316, n2722, n59315, 
        n2723, n59314, n33_adj_5223, n31_adj_5224, n59313, n59312, 
        n37_adj_5225, n35_adj_5226, n25_adj_5227, n27_adj_5228, n21_adj_5229, 
        n23_adj_5230, n59311, n9_adj_5231, n59310, n11_adj_5232, n19_adj_5233, 
        n13_adj_5234, n15_adj_5235, n17_adj_5236, n29_adj_5237, n75309, 
        n76273, n2728, n59309, n76738, n76736, n75313, n6_adj_5238, 
        n59308, n76920, n14_adj_5239, n32_adj_5240, n76921, n75299, 
        n12_adj_5241, n75295, n77295, n75987, n59307, n8_adj_5242, 
        n76922, n76923, n69405, n67179, n75324, n76255, n10_adj_5243, 
        n76998, n2596, n59306, n59305, n75985, n2598, n59304, 
        n2599, n59303, n77139, n2600, n59302, n77574, n59301, 
        n77213, n77647, n2602, n59300, n77648, n77636, n2603, 
        n59299, n77407, n2604, n59298, n2605, n59297, n2606, n59296, 
        n77408, n59295, n59294, n59293, n2610, n59292, n59291, 
        n59290, n69403, n67183, n2476, n59289, n2477, n59288, 
        n2478, n59287, n2479, n59286, n2480, n59285, n59284, n2482, 
        n59283, n2483, n59282, n59281, n2485, n59280, n59279, 
        n59278, n59277, n59276, n2490, n59275, n2491, n59274, 
        n69401, n2353, n59273, n59272, n59271, n2356, n59270, 
        n2357, n59269, n2358, n59268, n2359, n59267, n59266, n59265, 
        n59264, n2363, n59263, n2364, n59262, n59261, n59260, 
        n59259, n71560, n67221, n69399, n67191, n2227, n59258, 
        n59257, n58290, n2229, n59256, n2230, n59255, n2231, n59254, 
        n58289, n69351, n2232, n59253, n2233, n59252, n59251, 
        n2235, n59250, n58288, n69453, n59249, n59248, n65798, 
        n74542, n74539, n59247, n59246, n58287;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n74536, n59245, n69477, n69483, n69397, n59244, n59243, 
        n59242, n58286, n69451, n2101, n59241, n2102, n59240, 
        n58285, n69449, n2103, n59239, n2104, n59238, n2105, n59237, 
        n2106, n59236, n59235, n59234, n59233, n58284, n2110, 
        n59232, n59231, n59230, n1969, n59229, n1970, n59228, 
        n1971, n59227, n1972, n59226, n58283, n69447, n59225, 
        n59224, n59223, n58282, n69445, n59222, n59221, n58281, 
        n69349, n59220, n59219, n1833, n59218, n58280, n69443, 
        n1834, n59217, n1835, n59216, n1836, n59215, n1837, n59214, 
        n58279, n1838, n59213, n58278, n59212, n59211, n59210, 
        n69395, n67204, n58277, n1693, n59209, n1694, n59208, 
        n1695, n59207, n58276, n1696, n59206, n1697, n59205, n1698, 
        n59204, n1699, n59203, n1700, n59202, n59201, n58275, 
        n59200, n59199, n1554, n59198, n58274, n1555, n59197, 
        n21187, n44_adj_5244, n1556, n59196, n1557, n59195, n59194, 
        n58273, n59193, n1560, n59192, n59191, n1409, n59190, 
        n1410, n59189, n1411, n59188, n1412, n59187, n1413, n59186, 
        n59185, n59184, n69393, n59183, n59182, n59181, n1264, 
        n59180, n59179, n804, n44_adj_5245, n1266, n59178, n59177, 
        n67217, n1111, n59176, n1112, n59175, n58272, n1113, n59174, 
        n1114, n59173, n59172, n1116, n59171, n69389, n58271, 
        n58270, n58269, n58268, n58267, n59549, n59548, n59547, 
        n59546, n59545, n59544, n59543, n14_adj_5246, n15_adj_5247, 
        n4_adj_5248, n69875, n6_adj_5249, n42_adj_5250, n21179, n67659, 
        n42_adj_5251, n21189, n67643, n77085, n40_adj_5252, n74978, 
        n74903, n34_adj_5253, n77428, n77041, n35_adj_5254, n39_adj_5255, 
        n33_adj_5256, n37_adj_5257, n23_adj_5258, n25_adj_5259, n74551, 
        n27_adj_5260, n29_adj_5261, n74557, n74548, n74554, n11_adj_5262, 
        n31_adj_5263, n13_adj_5264, n21_adj_5265, n15_adj_5266, n17_adj_5267, 
        n19_adj_5268, n75366, n76329, n76768, n76764, n75368, n8_adj_5269, 
        n76930, n76931, n34_adj_5270, n75360, n77293, n75975, n76932, 
        n76933, n76305, n20_adj_5271, n75973, n77151, n77562, n76994, 
        n77631, n77632, n77040, n39_adj_5272, n45_adj_5273, n41_adj_5274, 
        n43_adj_5275, n33_adj_5276, n35_adj_5277, n37_adj_5278, n21_adj_5279, 
        n23_adj_5280, n29_adj_5281, n31_adj_5282, n25_adj_5283, n27_adj_5284, 
        n19_adj_5285, n74705, n74700, n76868, n18_adj_5286, n77042, 
        n77043, n75675, n26_adj_5287, n76985, n30_adj_5288, n77471, 
        n77472, n77272, n75679, n76986, n77250, n69945, n3_adj_5289, 
        n69949, n5, n69953, n8_adj_5290, n71462, n71534, n2, n69923, 
        n11915, n43_adj_5291, n37_adj_5292, n39_adj_5293, n41_adj_5294, 
        n67207, n32_adj_5295, n77072, n70749, n77073, n75884, n76588, 
        n76953, n77070, n77071, n48_adj_5296, n70747, n26027, n46, 
        n43_adj_5297, n38_adj_5298, n42_adj_5299, n77084, n40_adj_5300, 
        n26033, n803, n46_adj_5301, n44718, n67667, n644, n46_adj_5302, 
        n66908, n71500, n71516, n48_adj_5303, n25986, n67691, n5_adj_5304, 
        n69765, n71520, n71506, n69807, n71432, n71530, n71532, 
        n69873, n69877, n46_adj_5305, n42_adj_5306, n76602, n70649;
    
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n67224), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61251_3_lut (.I0(n42), .I1(baudrate[3]), .I2(n960), .I3(GND_net), 
            .O(n77086));   // verilog/uart_rx.v(119[33:55])
    defparam i61251_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61252_3_lut (.I0(n77086), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n77087));   // verilog/uart_rx.v(119[33:55])
    defparam i61252_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61104_3_lut (.I0(n77087), .I1(baudrate[5]), .I2(n66912), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i61104_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_3_lut (.I0(n71570), .I1(n48_adj_5023), .I2(baudrate[0]), 
            .I3(GND_net), .O(n962));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i59720_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i59720_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8291[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38), .I1(baudrate[4]), .I2(n41), 
            .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61624_4_lut (.I0(n40), .I1(n36), .I2(n41), .I3(n74972), 
            .O(n77459));   // verilog/uart_rx.v(119[33:55])
    defparam i61624_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61625_3_lut (.I0(n77459), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n77460));   // verilog/uart_rx.v(119[33:55])
    defparam i61625_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61453_3_lut (.I0(n77460), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n77288));   // verilog/uart_rx.v(119[33:55])
    defparam i61453_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61399_3_lut (.I0(n77288), .I1(baudrate[7]), .I2(n1261), .I3(GND_net), 
            .O(n48_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam i61399_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8317[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61243_3_lut (.I0(n34_c), .I1(baudrate[5]), .I2(n41_adj_5025), 
            .I3(GND_net), .O(n77078));   // verilog/uart_rx.v(119[33:55])
    defparam i61243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61244_3_lut (.I0(n77078), .I1(baudrate[6]), .I2(n43), .I3(GND_net), 
            .O(n77079));   // verilog/uart_rx.v(119[33:55])
    defparam i61244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60075_4_lut (.I0(n43), .I1(n41_adj_5025), .I2(n39), .I3(n74957), 
            .O(n75910));
    defparam i60075_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5026), .I1(baudrate[4]), 
            .I2(n39), .I3(GND_net), .O(n38_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61112_3_lut (.I0(n77079), .I1(baudrate[7]), .I2(n45), .I3(GND_net), 
            .O(n44));   // verilog/uart_rx.v(119[33:55])
    defparam i61112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60749_4_lut (.I0(n44), .I1(n38_adj_5027), .I2(n45), .I3(n75910), 
            .O(n76584));   // verilog/uart_rx.v(119[33:55])
    defparam i60749_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60750_3_lut (.I0(n76584), .I1(baudrate[8]), .I2(n1408), .I3(GND_net), 
            .O(n48_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam i60750_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut (.I0(n69391), .I1(n48_adj_5024), .I2(GND_net), .I3(GND_net), 
            .O(n1415));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8343[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61241_3_lut (.I0(n32), .I1(baudrate[5]), .I2(n39_adj_5029), 
            .I3(GND_net), .O(n77076));   // verilog/uart_rx.v(119[33:55])
    defparam i61241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61242_3_lut (.I0(n77076), .I1(baudrate[6]), .I2(n41_adj_5030), 
            .I3(GND_net), .O(n77077));   // verilog/uart_rx.v(119[33:55])
    defparam i61242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60065_4_lut (.I0(n41_adj_5030), .I1(n39_adj_5029), .I2(n37), 
            .I3(n74934), .O(n75900));
    defparam i60065_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60751_3_lut (.I0(n34_adj_5031), .I1(baudrate[4]), .I2(n37), 
            .I3(GND_net), .O(n76586));   // verilog/uart_rx.v(119[33:55])
    defparam i60751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61114_3_lut (.I0(n77077), .I1(baudrate[7]), .I2(n43_adj_5032), 
            .I3(GND_net), .O(n76949));   // verilog/uart_rx.v(119[33:55])
    defparam i61114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61239_4_lut (.I0(n76949), .I1(n76586), .I2(n43_adj_5032), 
            .I3(n75900), .O(n77074));   // verilog/uart_rx.v(119[33:55])
    defparam i61239_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61240_3_lut (.I0(n77074), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n77075));   // verilog/uart_rx.v(119[33:55])
    defparam i61240_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61116_3_lut (.I0(n77075), .I1(baudrate[9]), .I2(n1552), .I3(GND_net), 
            .O(n48_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam i61116_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51380_1_lut (.I0(n25974), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67167));
    defparam i51380_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_989 (.I0(n71554), .I1(n48_adj_5033), .I2(n8369[14]), 
            .I3(GND_net), .O(n1702));
    defparam i1_3_lut_adj_989.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8395[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59024_4_lut (.I0(n35), .I1(n33_c), .I2(n31), .I3(n29_c), 
            .O(n74859));
    defparam i59024_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5034), .I1(baudrate[9]), 
            .I2(n43_adj_5035), .I3(GND_net), .O(n40_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61233_3_lut (.I0(n28), .I1(baudrate[5]), .I2(n35), .I3(GND_net), 
            .O(n77068));   // verilog/uart_rx.v(119[33:55])
    defparam i61233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61234_3_lut (.I0(n77068), .I1(baudrate[6]), .I2(n37_adj_5037), 
            .I3(GND_net), .O(n77069));   // verilog/uart_rx.v(119[33:55])
    defparam i61234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59006_4_lut (.I0(n41_adj_5038), .I1(n39_adj_5039), .I2(n37_adj_5037), 
            .I3(n74859), .O(n74841));
    defparam i59006_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61231_4_lut (.I0(n40_adj_5036), .I1(n30), .I2(n43_adj_5035), 
            .I3(n74834), .O(n77066));   // verilog/uart_rx.v(119[33:55])
    defparam i61231_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61122_3_lut (.I0(n77069), .I1(baudrate[7]), .I2(n39_adj_5039), 
            .I3(GND_net), .O(n76957));   // verilog/uart_rx.v(119[33:55])
    defparam i61122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61691_4_lut (.I0(n76957), .I1(n77066), .I2(n43_adj_5035), 
            .I3(n74841), .O(n77526));   // verilog/uart_rx.v(119[33:55])
    defparam i61691_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61692_3_lut (.I0(n77526), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n77527));   // verilog/uart_rx.v(119[33:55])
    defparam i61692_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61592_3_lut (.I0(n77527), .I1(baudrate[11]), .I2(n1831), 
            .I3(GND_net), .O(n48_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam i61592_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8395[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8421[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8421[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58987_4_lut (.I0(n33_adj_5043), .I1(n31_adj_5042), .I2(n29_adj_5041), 
            .I3(n27_c), .O(n74822));
    defparam i58987_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i55717_1_lut (.I0(n71542), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67195));
    defparam i55717_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5044), .I1(baudrate[9]), 
            .I2(n41_adj_5045), .I3(GND_net), .O(n38_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61400_3_lut (.I0(n26), .I1(baudrate[5]), .I2(n33_adj_5043), 
            .I3(GND_net), .O(n77235));   // verilog/uart_rx.v(119[33:55])
    defparam i61400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61401_3_lut (.I0(n77235), .I1(baudrate[6]), .I2(n35_adj_5047), 
            .I3(GND_net), .O(n77236));   // verilog/uart_rx.v(119[33:55])
    defparam i61401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i58980_4_lut (.I0(n39_adj_5048), .I1(n37_adj_5049), .I2(n35_adj_5047), 
            .I3(n74822), .O(n74815));
    defparam i58980_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61626_4_lut (.I0(n38_adj_5046), .I1(n28_adj_5050), .I2(n41_adj_5045), 
            .I3(n74813), .O(n77461));   // verilog/uart_rx.v(119[33:55])
    defparam i61626_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61126_3_lut (.I0(n77236), .I1(baudrate[7]), .I2(n37_adj_5049), 
            .I3(GND_net), .O(n76961));   // verilog/uart_rx.v(119[33:55])
    defparam i61126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61790_4_lut (.I0(n76961), .I1(n77461), .I2(n41_adj_5045), 
            .I3(n74815), .O(n77625));   // verilog/uart_rx.v(119[33:55])
    defparam i61790_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61791_3_lut (.I0(n77625), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n77626));   // verilog/uart_rx.v(119[33:55])
    defparam i61791_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61769_3_lut (.I0(n77626), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n77604));   // verilog/uart_rx.v(119[33:55])
    defparam i61769_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61702_3_lut (.I0(n77604), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam i61702_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8421[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8447[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n70773), .I1(n9), .I2(n14), .I3(n70643), .O(n26008));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58964_4_lut (.I0(n33_adj_5053), .I1(n31_adj_5054), .I2(n29_adj_5055), 
            .I3(n27_adj_5052), .O(n74799));
    defparam i58964_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5056), .I1(baudrate[10]), 
            .I2(n41_adj_5057), .I3(GND_net), .O(n38_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30681_rep_4_2_lut (.I0(n8447[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n67198));   // verilog/uart_rx.v(119[33:55])
    defparam i30681_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n67198), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61227_3_lut (.I0(n26_adj_5059), .I1(baudrate[6]), .I2(n33_adj_5053), 
            .I3(GND_net), .O(n77062));   // verilog/uart_rx.v(119[33:55])
    defparam i61227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61228_3_lut (.I0(n77062), .I1(baudrate[7]), .I2(n35_adj_5060), 
            .I3(GND_net), .O(n77063));   // verilog/uart_rx.v(119[33:55])
    defparam i61228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i58960_4_lut (.I0(n39_adj_5061), .I1(n37_adj_5062), .I2(n35_adj_5060), 
            .I3(n74799), .O(n74795));
    defparam i58960_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61628_4_lut (.I0(n38_adj_5058), .I1(n28_adj_5063), .I2(n41_adj_5057), 
            .I3(n74790), .O(n77463));   // verilog/uart_rx.v(119[33:55])
    defparam i61628_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61132_3_lut (.I0(n77063), .I1(baudrate[8]), .I2(n37_adj_5062), 
            .I3(GND_net), .O(n76967));   // verilog/uart_rx.v(119[33:55])
    defparam i61132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61792_4_lut (.I0(n76967), .I1(n77463), .I2(n41_adj_5057), 
            .I3(n74795), .O(n77627));   // verilog/uart_rx.v(119[33:55])
    defparam i61792_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61793_3_lut (.I0(n77627), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n77628));   // verilog/uart_rx.v(119[33:55])
    defparam i61793_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61767_3_lut (.I0(n77628), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n77602));   // verilog/uart_rx.v(119[33:55])
    defparam i61767_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61704_3_lut (.I0(n77602), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam i61704_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8447[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8473[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8473[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i55712_4_lut (.I0(n70817), .I1(n9), .I2(n70805), .I3(baudrate[17]), 
            .O(n71538));
    defparam i55712_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i55716_4_lut (.I0(n71510), .I1(n71538), .I2(n14), .I3(n71430), 
            .O(n71542));
    defparam i55716_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58923_4_lut (.I0(n29_adj_5066), .I1(n27_adj_5065), .I2(n25), 
            .I3(n23_c), .O(n74758));
    defparam i58923_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i58919_4_lut (.I0(n35_adj_5067), .I1(n33_adj_5068), .I2(n31_adj_5069), 
            .I3(n74758), .O(n74754));
    defparam i58919_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5070), .I1(baudrate[7]), 
            .I2(n33_adj_5068), .I3(GND_net), .O(n30_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5072), .I1(baudrate[9]), 
            .I2(n37_adj_5073), .I3(GND_net), .O(n34_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61630_4_lut (.I0(n34_adj_5074), .I1(n24), .I2(n37_adj_5073), 
            .I3(n74752), .O(n77465));   // verilog/uart_rx.v(119[33:55])
    defparam i61630_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61631_3_lut (.I0(n77465), .I1(baudrate[10]), .I2(n39_adj_5075), 
            .I3(GND_net), .O(n77466));   // verilog/uart_rx.v(119[33:55])
    defparam i61631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61443_3_lut (.I0(n77466), .I1(baudrate[11]), .I2(n41_adj_5076), 
            .I3(GND_net), .O(n77278));   // verilog/uart_rx.v(119[33:55])
    defparam i61443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61037_4_lut (.I0(n41_adj_5076), .I1(n39_adj_5075), .I2(n37_adj_5073), 
            .I3(n74754), .O(n76872));
    defparam i61037_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61217_4_lut (.I0(n30_adj_5071), .I1(n22), .I2(n33_adj_5068), 
            .I3(n74756), .O(n77052));   // verilog/uart_rx.v(119[33:55])
    defparam i61217_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61407_3_lut (.I0(n77278), .I1(baudrate[12]), .I2(n43_adj_5077), 
            .I3(GND_net), .O(n42_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam i61407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61474_4_lut (.I0(n42_adj_5078), .I1(n77052), .I2(n43_adj_5077), 
            .I3(n76872), .O(n77309));   // verilog/uart_rx.v(119[33:55])
    defparam i61474_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61475_3_lut (.I0(n77309), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n77310));   // verilog/uart_rx.v(119[33:55])
    defparam i61475_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8473[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8499[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8499[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8499[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_990 (.I0(n14), .I1(n9), .I2(n70793), .I3(n70769), 
            .O(n26014));
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58900_4_lut (.I0(n27_adj_5082), .I1(n25_adj_5083), .I2(n23_adj_5084), 
            .I3(n21), .O(n74735));
    defparam i58900_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i58896_4_lut (.I0(n33_adj_5081), .I1(n31_adj_5080), .I2(n29_adj_5079), 
            .I3(n74735), .O(n74731));
    defparam i58896_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5085), .I1(baudrate[7]), 
            .I2(n31_adj_5080), .I3(GND_net), .O(n28_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5087), .I1(baudrate[9]), 
            .I2(n35_adj_5088), .I3(GND_net), .O(n32_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61632_4_lut (.I0(n32_adj_5089), .I1(n22_adj_5090), .I2(n35_adj_5088), 
            .I3(n74729), .O(n77467));   // verilog/uart_rx.v(119[33:55])
    defparam i61632_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61633_3_lut (.I0(n77467), .I1(baudrate[10]), .I2(n37_adj_5091), 
            .I3(GND_net), .O(n77468));   // verilog/uart_rx.v(119[33:55])
    defparam i61633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61441_3_lut (.I0(n77468), .I1(baudrate[11]), .I2(n39_adj_5092), 
            .I3(GND_net), .O(n77276));   // verilog/uart_rx.v(119[33:55])
    defparam i61441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61035_4_lut (.I0(n39_adj_5092), .I1(n37_adj_5091), .I2(n35_adj_5088), 
            .I3(n74731), .O(n76870));
    defparam i61035_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61634_4_lut (.I0(n28_adj_5086), .I1(n20), .I2(n31_adj_5080), 
            .I3(n74733), .O(n77469));   // verilog/uart_rx.v(119[33:55])
    defparam i61634_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61409_3_lut (.I0(n77276), .I1(baudrate[12]), .I2(n41_adj_5093), 
            .I3(GND_net), .O(n77244));   // verilog/uart_rx.v(119[33:55])
    defparam i61409_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n28238), 
            .D(n479[1]), .R(n67079));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i61699_4_lut (.I0(n77244), .I1(n77469), .I2(n41_adj_5093), 
            .I3(n76870), .O(n77534));   // verilog/uart_rx.v(119[33:55])
    defparam i61699_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61700_3_lut (.I0(n77534), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n77535));   // verilog/uart_rx.v(119[33:55])
    defparam i61700_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61639_3_lut (.I0(n77535), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n77474));   // verilog/uart_rx.v(119[33:55])
    defparam i61639_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8499[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8525[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8551[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n28238), 
            .D(n479[2]), .R(n67079));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59815_4_lut (.I0(n23_adj_5094), .I1(n21_adj_5096), .I2(n19), 
            .I3(n17), .O(n75650));
    defparam i59815_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59806_4_lut (.I0(n29_adj_5097), .I1(n27_adj_5098), .I2(n25_adj_5095), 
            .I3(n75650), .O(n75641));
    defparam i59806_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61350_4_lut (.I0(n35_adj_5099), .I1(n33_adj_5100), .I2(n31_adj_5101), 
            .I3(n75641), .O(n77185));
    defparam i61350_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61179_3_lut (.I0(n16), .I1(baudrate[13]), .I2(n39_adj_5102), 
            .I3(GND_net), .O(n77014));   // verilog/uart_rx.v(119[33:55])
    defparam i61179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61180_3_lut (.I0(n77014), .I1(baudrate[14]), .I2(n41_adj_5103), 
            .I3(GND_net), .O(n77015));   // verilog/uart_rx.v(119[33:55])
    defparam i61180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60642_4_lut (.I0(n41_adj_5103), .I1(n39_adj_5102), .I2(n27_adj_5098), 
            .I3(n75643), .O(n76477));
    defparam i60642_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61153_3_lut (.I0(n22_adj_5104), .I1(baudrate[7]), .I2(n27_adj_5098), 
            .I3(GND_net), .O(n76988));   // verilog/uart_rx.v(119[33:55])
    defparam i61153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60106_3_lut (.I0(n77015), .I1(baudrate[15]), .I2(n43_adj_5105), 
            .I3(GND_net), .O(n75941));   // verilog/uart_rx.v(119[33:55])
    defparam i60106_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5106), .I1(baudrate[9]), 
            .I2(n31_adj_5101), .I3(GND_net), .O(n28_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61426_4_lut (.I0(n28_adj_5107), .I1(n18), .I2(n31_adj_5101), 
            .I3(n75639), .O(n77261));   // verilog/uart_rx.v(119[33:55])
    defparam i61426_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61427_3_lut (.I0(n77261), .I1(baudrate[10]), .I2(n33_adj_5100), 
            .I3(GND_net), .O(n77262));   // verilog/uart_rx.v(119[33:55])
    defparam i61427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61425_3_lut (.I0(n77262), .I1(baudrate[11]), .I2(n35_adj_5099), 
            .I3(GND_net), .O(n77260));   // verilog/uart_rx.v(119[33:55])
    defparam i61425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60644_4_lut (.I0(n41_adj_5103), .I1(n39_adj_5102), .I2(n37_adj_5108), 
            .I3(n77185), .O(n76479));
    defparam i60644_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61175_4_lut (.I0(n75941), .I1(n76988), .I2(n43_adj_5105), 
            .I3(n76477), .O(n77010));   // verilog/uart_rx.v(119[33:55])
    defparam i61175_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60104_3_lut (.I0(n77260), .I1(baudrate[12]), .I2(n37_adj_5108), 
            .I3(GND_net), .O(n75939));   // verilog/uart_rx.v(119[33:55])
    defparam i60104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61708_4_lut (.I0(n75939), .I1(n77010), .I2(n43_adj_5105), 
            .I3(n76479), .O(n77543));   // verilog/uart_rx.v(119[33:55])
    defparam i61708_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61709_3_lut (.I0(n77543), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n77544));   // verilog/uart_rx.v(119[33:55])
    defparam i61709_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8551[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8577[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8577[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_991 (.I0(n69941), .I1(n70809), .I2(n70799), .I3(baudrate[19]), 
            .O(n25965));
    defparam i1_4_lut_adj_991.LUT_INIT = 16'hfffe;
    SB_LUT4 i59704_4_lut (.I0(n37_adj_5112), .I1(n25_adj_5111), .I2(n23_adj_5110), 
            .I3(n21_adj_5109), .O(n75539));
    defparam i59704_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60630_4_lut (.I0(n19_adj_5113), .I1(n17_adj_5114), .I2(n2729), 
            .I3(baudrate[2]), .O(n76465));
    defparam i60630_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i61001_4_lut (.I0(n25_adj_5111), .I1(n23_adj_5110), .I2(n21_adj_5109), 
            .I3(n76465), .O(n76836));
    defparam i61001_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60999_4_lut (.I0(n31_adj_5115), .I1(n29_adj_5116), .I2(n27_adj_5117), 
            .I3(n76836), .O(n76834));
    defparam i60999_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59706_4_lut (.I0(n37_adj_5112), .I1(n35_adj_5118), .I2(n33_adj_5119), 
            .I3(n76834), .O(n75541));
    defparam i59706_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61169_3_lut (.I0(n14_adj_5120), .I1(baudrate[13]), .I2(n37_adj_5112), 
            .I3(GND_net), .O(n77004));   // verilog/uart_rx.v(119[33:55])
    defparam i61169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61170_3_lut (.I0(n77004), .I1(baudrate[14]), .I2(n39_adj_5121), 
            .I3(GND_net), .O(n77005));   // verilog/uart_rx.v(119[33:55])
    defparam i61170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_5122), .I1(baudrate[17]), 
            .I2(n45_adj_5123), .I3(GND_net), .O(n40_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59699_4_lut (.I0(n43_adj_5125), .I1(n41_adj_5126), .I2(n39_adj_5121), 
            .I3(n75539), .O(n75534));
    defparam i59699_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61155_4_lut (.I0(n40_adj_5124), .I1(n20_adj_5127), .I2(n45_adj_5123), 
            .I3(n75532), .O(n76990));   // verilog/uart_rx.v(119[33:55])
    defparam i61155_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60116_3_lut (.I0(n77005), .I1(baudrate[15]), .I2(n41_adj_5126), 
            .I3(GND_net), .O(n75951));   // verilog/uart_rx.v(119[33:55])
    defparam i60116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5128), .I1(baudrate[9]), 
            .I2(n29_adj_5116), .I3(GND_net), .O(n26_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61428_4_lut (.I0(n26_adj_5129), .I1(n16_adj_5130), .I2(n29_adj_5116), 
            .I3(n75575), .O(n77263));   // verilog/uart_rx.v(119[33:55])
    defparam i61428_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61429_3_lut (.I0(n77263), .I1(baudrate[10]), .I2(n31_adj_5115), 
            .I3(GND_net), .O(n77264));   // verilog/uart_rx.v(119[33:55])
    defparam i61429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61421_3_lut (.I0(n77264), .I1(baudrate[11]), .I2(n33_adj_5119), 
            .I3(GND_net), .O(n77256));   // verilog/uart_rx.v(119[33:55])
    defparam i61421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61344_4_lut (.I0(n43_adj_5125), .I1(n41_adj_5126), .I2(n39_adj_5121), 
            .I3(n75541), .O(n77179));
    defparam i61344_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61595_4_lut (.I0(n75951), .I1(n76990), .I2(n45_adj_5123), 
            .I3(n75534), .O(n77430));   // verilog/uart_rx.v(119[33:55])
    defparam i61595_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60114_3_lut (.I0(n77256), .I1(baudrate[12]), .I2(n35_adj_5118), 
            .I3(GND_net), .O(n75949));   // verilog/uart_rx.v(119[33:55])
    defparam i60114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61597_4_lut (.I0(n75949), .I1(n77430), .I2(n45_adj_5123), 
            .I3(n77179), .O(n77432));   // verilog/uart_rx.v(119[33:55])
    defparam i61597_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8577[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8603[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8603[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_992 (.I0(n70767), .I1(n14), .I2(n9), .I3(n70803), 
            .O(n25968));
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i59656_4_lut (.I0(n35_adj_5134), .I1(n23_adj_5133), .I2(n21_adj_5132), 
            .I3(n19_adj_5131), .O(n75491));
    defparam i59656_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60588_4_lut (.I0(n17_adj_5135), .I1(n15), .I2(n2844), .I3(baudrate[2]), 
            .O(n76423));
    defparam i60588_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i60983_4_lut (.I0(n23_adj_5133), .I1(n21_adj_5132), .I2(n19_adj_5131), 
            .I3(n76423), .O(n76818));
    defparam i60983_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60981_4_lut (.I0(n29_adj_5136), .I1(n27_adj_5137), .I2(n25_adj_5138), 
            .I3(n76818), .O(n76816));
    defparam i60981_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59658_4_lut (.I0(n35_adj_5134), .I1(n33_adj_5139), .I2(n31_adj_5140), 
            .I3(n76816), .O(n75493));
    defparam i59658_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61129_3_lut (.I0(n12), .I1(baudrate[13]), .I2(n35_adj_5134), 
            .I3(GND_net), .O(n76964));   // verilog/uart_rx.v(119[33:55])
    defparam i61129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5141), .I1(baudrate[17]), 
            .I2(n43_adj_5142), .I3(GND_net), .O(n38_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61130_3_lut (.I0(n76964), .I1(baudrate[14]), .I2(n37_adj_5144), 
            .I3(GND_net), .O(n76965));   // verilog/uart_rx.v(119[33:55])
    defparam i61130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59646_4_lut (.I0(n41_adj_5145), .I1(n39_adj_5146), .I2(n37_adj_5144), 
            .I3(n75491), .O(n75481));
    defparam i59646_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61432_4_lut (.I0(n38_adj_5143), .I1(n18_adj_5147), .I2(n43_adj_5142), 
            .I3(n75468), .O(n77267));   // verilog/uart_rx.v(119[33:55])
    defparam i61432_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60122_3_lut (.I0(n76965), .I1(baudrate[15]), .I2(n39_adj_5146), 
            .I3(GND_net), .O(n75957));   // verilog/uart_rx.v(119[33:55])
    defparam i60122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5148), .I1(baudrate[9]), 
            .I2(n27_adj_5137), .I3(GND_net), .O(n24_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61434_4_lut (.I0(n24_adj_5149), .I1(n14_adj_5150), .I2(n27_adj_5137), 
            .I3(n75507), .O(n77269));   // verilog/uart_rx.v(119[33:55])
    defparam i61434_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61435_3_lut (.I0(n77269), .I1(baudrate[10]), .I2(n29_adj_5136), 
            .I3(GND_net), .O(n77270));   // verilog/uart_rx.v(119[33:55])
    defparam i61435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61417_3_lut (.I0(n77270), .I1(baudrate[11]), .I2(n31_adj_5140), 
            .I3(GND_net), .O(n77252));   // verilog/uart_rx.v(119[33:55])
    defparam i61417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61336_4_lut (.I0(n41_adj_5145), .I1(n39_adj_5146), .I2(n37_adj_5144), 
            .I3(n75493), .O(n77171));
    defparam i61336_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61764_4_lut (.I0(n75957), .I1(n77267), .I2(n43_adj_5142), 
            .I3(n75481), .O(n77599));   // verilog/uart_rx.v(119[33:55])
    defparam i61764_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60120_3_lut (.I0(n77252), .I1(baudrate[12]), .I2(n33_adj_5139), 
            .I3(GND_net), .O(n75955));   // verilog/uart_rx.v(119[33:55])
    defparam i60120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61798_4_lut (.I0(n75955), .I1(n77599), .I2(n43_adj_5142), 
            .I3(n77171), .O(n77633));   // verilog/uart_rx.v(119[33:55])
    defparam i61798_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61799_3_lut (.I0(n77633), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n77634));   // verilog/uart_rx.v(119[33:55])
    defparam i61799_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8603[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8629[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8629[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_993 (.I0(baudrate[31]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n70817));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_994 (.I0(baudrate[30]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n70819));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_995 (.I0(n70821), .I1(n14), .I2(n9), .I3(n70819), 
            .O(n25971));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'hfffe;
    SB_LUT4 i59599_4_lut (.I0(n33_adj_5154), .I1(n21_adj_5153), .I2(n19_adj_5152), 
            .I3(n17_adj_5151), .O(n75434));
    defparam i59599_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60542_4_lut (.I0(n15_adj_5155), .I1(n13), .I2(n2956), .I3(baudrate[2]), 
            .O(n76377));
    defparam i60542_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i60961_4_lut (.I0(n21_adj_5153), .I1(n19_adj_5152), .I2(n17_adj_5151), 
            .I3(n76377), .O(n76796));
    defparam i60961_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59099_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n74934));   // verilog/uart_rx.v(119[33:55])
    defparam i59099_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i60957_4_lut (.I0(n27_adj_5156), .I1(n25_adj_5157), .I2(n23_adj_5158), 
            .I3(n76796), .O(n76792));
    defparam i60957_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59601_4_lut (.I0(n33_adj_5154), .I1(n31_adj_5159), .I2(n29_adj_5160), 
            .I3(n76792), .O(n75436));
    defparam i59601_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61101_3_lut (.I0(n10), .I1(baudrate[13]), .I2(n33_adj_5154), 
            .I3(GND_net), .O(n76936));   // verilog/uart_rx.v(119[33:55])
    defparam i61101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61102_3_lut (.I0(n76936), .I1(baudrate[14]), .I2(n35_adj_5161), 
            .I3(GND_net), .O(n76937));   // verilog/uart_rx.v(119[33:55])
    defparam i61102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5162), .I1(baudrate[17]), 
            .I2(n41_adj_5163), .I3(GND_net), .O(n36_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59590_4_lut (.I0(n39_adj_5165), .I1(n37_adj_5166), .I2(n35_adj_5161), 
            .I3(n75434), .O(n75425));
    defparam i59590_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61456_4_lut (.I0(n36_adj_5164), .I1(n16_adj_5167), .I2(n41_adj_5163), 
            .I3(n75419), .O(n77291));   // verilog/uart_rx.v(119[33:55])
    defparam i61456_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60128_3_lut (.I0(n76937), .I1(baudrate[15]), .I2(n37_adj_5166), 
            .I3(GND_net), .O(n75963));   // verilog/uart_rx.v(119[33:55])
    defparam i60128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5168), .I1(baudrate[9]), 
            .I2(n25_adj_5157), .I3(GND_net), .O(n22_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61454_4_lut (.I0(n22_adj_5169), .I1(n12_adj_5170), .I2(n25_adj_5157), 
            .I3(n75448), .O(n77289));   // verilog/uart_rx.v(119[33:55])
    defparam i61454_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61455_3_lut (.I0(n77289), .I1(baudrate[10]), .I2(n27_adj_5156), 
            .I3(GND_net), .O(n77290));   // verilog/uart_rx.v(119[33:55])
    defparam i61455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61397_3_lut (.I0(n77290), .I1(baudrate[11]), .I2(n29_adj_5160), 
            .I3(GND_net), .O(n77232));   // verilog/uart_rx.v(119[33:55])
    defparam i61397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61326_4_lut (.I0(n39_adj_5165), .I1(n37_adj_5166), .I2(n35_adj_5161), 
            .I3(n75436), .O(n77161));
    defparam i61326_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61689_4_lut (.I0(n75963), .I1(n77291), .I2(n41_adj_5163), 
            .I3(n75425), .O(n77524));   // verilog/uart_rx.v(119[33:55])
    defparam i61689_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60126_3_lut (.I0(n77232), .I1(baudrate[12]), .I2(n31_adj_5159), 
            .I3(GND_net), .O(n75961));   // verilog/uart_rx.v(119[33:55])
    defparam i60126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61810_4_lut (.I0(n75961), .I1(n77524), .I2(n41_adj_5163), 
            .I3(n77161), .O(n77645));   // verilog/uart_rx.v(119[33:55])
    defparam i61810_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61811_3_lut (.I0(n77645), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n77646));   // verilog/uart_rx.v(119[33:55])
    defparam i61811_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61805_3_lut (.I0(n77646), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n77640));   // verilog/uart_rx.v(119[33:55])
    defparam i61805_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8629[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8655[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8681[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51400_1_lut (.I0(n26017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67187));
    defparam i51400_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i55731_1_lut_2_lut (.I0(baudrate[9]), .I1(n71554), .I2(GND_net), 
            .I3(GND_net), .O(n67213));
    defparam i55731_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i55670_2_lut_4_lut (.I0(baudrate[6]), .I1(baudrate[7]), .I2(baudrate[8]), 
            .I3(baudrate[9]), .O(n71496));
    defparam i55670_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[27]), .I2(n14), 
            .I3(n70767), .O(n25974));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i62481_2_lut_4_lut (.I0(n76603), .I1(baudrate[4]), .I2(n66910), 
            .I3(n71570), .O(n294[19]));
    defparam i62481_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i59042_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5171), .I2(n25989), 
            .I3(GND_net), .O(n74877));   // verilog/uart_rx.v(119[33:55])
    defparam i59042_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_996 (.I0(n25989), .I1(n48_adj_5171), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5172));
    defparam i1_3_lut_4_lut_adj_996.LUT_INIT = 16'hefff;
    SB_LUT4 i51384_1_lut_4_lut (.I0(n70821), .I1(n14), .I2(n9), .I3(n70819), 
            .O(n67171));
    defparam i51384_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i59718_2_lut_3_lut (.I0(n25989), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n74573));   // verilog/uart_rx.v(119[33:55])
    defparam i59718_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i55728_2_lut_3_lut_4_lut (.I0(baudrate[12]), .I1(n71544), .I2(baudrate[10]), 
            .I3(baudrate[11]), .O(n71554));
    defparam i55728_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), .I2(n71574), 
            .I3(GND_net), .O(n45239));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_997 (.I0(baudrate[14]), .I1(baudrate[2]), 
            .I2(baudrate[1]), .I3(baudrate[0]), .O(n69833));
    defparam i1_3_lut_4_lut_adj_997.LUT_INIT = 16'h1000;
    SB_LUT4 i59047_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5173), .I2(n26020), 
            .I3(GND_net), .O(n74882));   // verilog/uart_rx.v(119[33:55])
    defparam i59047_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i7309_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21177));   // verilog/uart_rx.v(119[33:55])
    defparam i7309_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i62403_3_lut_4_lut_3_lut (.I0(n71574), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n71578));
    defparam i62403_3_lut_4_lut_3_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5828_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11690));   // verilog/uart_rx.v(119[33:55])
    defparam i5828_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i62601_2_lut_4_lut (.I0(n77075), .I1(baudrate[9]), .I2(n1552), 
            .I3(n71554), .O(n294[14]));
    defparam i62601_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i55672_2_lut_3_lut_4_lut (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[10]), .I3(baudrate[11]), .O(n71498));
    defparam i55672_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n28_adj_5174));
    defparam i10_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58863_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n74698));
    defparam i58863_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i62592_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n71554), .I2(n48_adj_5024), 
            .I3(baudrate[8]), .O(n294[16]));
    defparam i62592_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58868_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n74703));
    defparam i58868_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n14), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(n70773), .O(n25935));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5178));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_2_lut (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5179));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_2_lut (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5180));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i62595_2_lut_3_lut (.I0(baudrate[9]), .I1(n71554), .I2(n48_adj_5028), 
            .I3(GND_net), .O(n294[15]));
    defparam i62595_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_2903_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n59407), 
            .O(n8707[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2903_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n59406), 
            .O(n8707[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_24 (.CI(n59406), .I0(n3152), .I1(n3082), .CO(n59407));
    SB_LUT4 add_2903_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n59405), 
            .O(n8707[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_23 (.CI(n59405), .I0(n3153), .I1(n3188), .CO(n59406));
    SB_LUT4 add_2903_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n59404), 
            .O(n8707[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n69971));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_CARRY add_2903_22 (.CI(n59404), .I0(n3154), .I1(n3084), .CO(n59405));
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59521_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n75356));
    defparam i59521_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2903_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n59403), 
            .O(n8707[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_21 (.CI(n59403), .I0(n3155), .I1(n2977), .CO(n59404));
    SB_LUT4 add_2903_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n59402), 
            .O(n8707[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_20 (.CI(n59402), .I0(n3156), .I1(n2867), .CO(n59403));
    SB_LUT4 add_2903_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n59401), 
            .O(n8707[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2903_19 (.CI(n59401), .I0(n3157), .I1(n2754), .CO(n59402));
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2903_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n59400), 
            .O(n8707[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_18 (.CI(n59400), .I0(n3158), .I1(n2638), .CO(n59401));
    SB_LUT4 add_2903_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n59399), 
            .O(n8707[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut (.I0(n69971), .I1(n23_adj_5180), .I2(n22_adj_5179), 
            .I3(n24_adj_5178), .O(n33));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_999 (.I0(baudrate[31]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n70801));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n70803));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'heeee;
    SB_CARRY add_2903_17 (.CI(n59399), .I0(n3159), .I1(n2519), .CO(n59400));
    SB_LUT4 add_2903_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n59398), 
            .O(n8707[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'heeee;
    SB_CARRY add_2903_16 (.CI(n59398), .I0(n3160), .I1(n2397), .CO(n59399));
    SB_LUT4 add_2903_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n59397), 
            .O(n8707[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1002 (.I0(baudrate[24]), .I1(baudrate[26]), .I2(baudrate[25]), 
            .I3(baudrate[29]), .O(n14));
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_CARRY add_2903_15 (.CI(n59397), .I0(n3161), .I1(n2272), .CO(n59398));
    SB_LUT4 i1_2_lut_adj_1003 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n70805));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'heeee;
    SB_LUT4 i59547_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n75382));
    defparam i59547_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n70799));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1005 (.I0(n70799), .I1(n70805), .I2(baudrate[17]), 
            .I3(GND_net), .O(n70811));
    defparam i1_3_lut_adj_1005.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(n14), .I1(n9), .I2(n70811), .I3(n70809), 
            .O(n26017));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'hfffe;
    SB_LUT4 i30642_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44716));
    defparam i30642_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut (.I0(n70745), .I1(baudrate[16]), .I2(n28_adj_5174), 
            .I3(n26017), .O(n34));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2903_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n59396), 
            .O(n8707[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_14 (.CI(n59396), .I0(n3162), .I1(n2144), .CO(n59397));
    SB_LUT4 add_2903_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n59395), 
            .O(n8707[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29935));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29934));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29932));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29913));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29912));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29908));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29904));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i59736_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5215), .I3(n66050), .O(n74514));
    defparam i59736_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i59733_4_lut (.I0(n74514), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n74511));
    defparam i59733_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n74511), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n28115));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n79053));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Clock_Count_2053__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n28159), .D(n1[0]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n28159), .D(n1[1]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n28159), .D(n1[2]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n28159), .D(n1[3]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n28159), .D(n1[4]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n28159), .D(n1[5]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n28159), .D(n1[6]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n28159), .D(n1[7]), .R(n29421));   // verilog/uart_rx.v(121[34:51])
    SB_CARRY add_2903_13 (.CI(n59395), .I0(n3163), .I1(n2013), .CO(n59396));
    SB_LUT4 add_2903_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n59394), 
            .O(n8707[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_12 (.CI(n59394), .I0(n3164), .I1(n1879), .CO(n59395));
    SB_LUT4 add_2903_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n59393), 
            .O(n8707[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_11 (.CI(n59393), .I0(n3165), .I1(n1742), .CO(n59394));
    SB_LUT4 add_2903_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n59392), 
            .O(n8707[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_10 (.CI(n59392), .I0(n3166), .I1(n1602), .CO(n59393));
    SB_LUT4 add_2903_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n59391), 
            .O(n8707[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_9 (.CI(n59391), .I0(n3167), .I1(n1459), .CO(n59392));
    SB_LUT4 add_2903_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n59390), 
            .O(n8707[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_8 (.CI(n59390), .I0(n3168), .I1(n1460), .CO(n59391));
    SB_LUT4 add_2903_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n59389), 
            .O(n8707[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_7 (.CI(n59389), .I0(n3169), .I1(n1011), .CO(n59390));
    SB_LUT4 add_2903_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n59388), 
            .O(n8707[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_6 (.CI(n59388), .I0(n3170), .I1(n856), .CO(n59389));
    SB_LUT4 add_2903_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n59387), 
            .O(n8707[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_5 (.CI(n59387), .I0(n3171), .I1(n698), .CO(n59388));
    SB_LUT4 add_2903_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n59386), 
            .O(n8707[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2903_4 (.CI(n59386), .I0(n3172), .I1(n858), .CO(n59387));
    SB_LUT4 add_2903_3_lut (.I0(n67163), .I1(GND_net), .I2(n538), .I3(n59385), 
            .O(n69413)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2903_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2903_3 (.CI(n59385), .I0(GND_net), .I1(n538), .CO(n59386));
    SB_CARRY add_2903_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n59385));
    SB_LUT4 add_2902_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n59384), 
            .O(n8681[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2902_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n59383), 
            .O(n8681[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_22 (.CI(n59383), .I0(n3047), .I1(n3188), .CO(n59384));
    SB_LUT4 add_2902_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n59382), 
            .O(n8681[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_21 (.CI(n59382), .I0(n3048), .I1(n3084), .CO(n59383));
    SB_LUT4 add_2902_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n59381), 
            .O(n8681[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_20 (.CI(n59381), .I0(n3049), .I1(n2977), .CO(n59382));
    SB_LUT4 add_2902_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n59380), 
            .O(n8681[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_19 (.CI(n59380), .I0(n3050), .I1(n2867), .CO(n59381));
    SB_LUT4 add_2902_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n59379), 
            .O(n8681[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_18 (.CI(n59379), .I0(n3051), .I1(n2754), .CO(n59380));
    SB_LUT4 add_2902_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n59378), 
            .O(n8681[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_17 (.CI(n59378), .I0(n3052), .I1(n2638), .CO(n59379));
    SB_LUT4 add_2902_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n59377), 
            .O(n8681[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_16 (.CI(n59377), .I0(n3053), .I1(n2519), .CO(n59378));
    SB_LUT4 add_2902_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n59376), 
            .O(n8681[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30760));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n61786));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30756));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2902_15 (.CI(n59376), .I0(n3054), .I1(n2397), .CO(n59377));
    SB_LUT4 add_2902_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n59375), 
            .O(n8681[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_14 (.CI(n59375), .I0(n3055), .I1(n2272), .CO(n59376));
    SB_LUT4 add_2902_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n59374), 
            .O(n8681[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_13 (.CI(n59374), .I0(n3056), .I1(n2144), .CO(n59375));
    SB_LUT4 add_2902_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n59373), 
            .O(n8681[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_12 (.CI(n59373), .I0(n3057), .I1(n2013), .CO(n59374));
    SB_LUT4 add_2902_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n59372), 
            .O(n8681[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_11 (.CI(n59372), .I0(n3058), .I1(n1879), .CO(n59373));
    SB_LUT4 add_2902_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n59371), 
            .O(n8681[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_10 (.CI(n59371), .I0(n3059), .I1(n1742), .CO(n59372));
    SB_LUT4 add_2902_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n59370), 
            .O(n8681[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_9 (.CI(n59370), .I0(n3060), .I1(n1602), .CO(n59371));
    SB_LUT4 add_2902_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n59369), 
            .O(n8681[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_8 (.CI(n59369), .I0(n3061), .I1(n1459), .CO(n59370));
    SB_LUT4 add_2902_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n59368), 
            .O(n8681[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_7 (.CI(n59368), .I0(n3062), .I1(n1460), .CO(n59369));
    SB_LUT4 add_2902_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n59367), 
            .O(n8681[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_6 (.CI(n59367), .I0(n3063), .I1(n1011), .CO(n59368));
    SB_LUT4 add_2902_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n59366), 
            .O(n8681[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_5 (.CI(n59366), .I0(n3064), .I1(n856), .CO(n59367));
    SB_LUT4 add_2902_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n59365), 
            .O(n8681[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_4 (.CI(n59365), .I0(n3065), .I1(n698), .CO(n59366));
    SB_LUT4 add_2902_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n59364), 
            .O(n8681[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2902_3 (.CI(n59364), .I0(n3066), .I1(n858), .CO(n59365));
    SB_LUT4 add_2902_2_lut (.I0(n67167), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69411)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2902_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2902_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59364));
    SB_LUT4 add_2901_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n59363), 
            .O(n8655[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2901_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n59362), 
            .O(n8655[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_21 (.CI(n59362), .I0(n2939), .I1(n3084), .CO(n59363));
    SB_LUT4 add_2901_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n59361), 
            .O(n8655[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_20 (.CI(n59361), .I0(n2940), .I1(n2977), .CO(n59362));
    SB_LUT4 add_2901_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n59360), 
            .O(n8655[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_19 (.CI(n59360), .I0(n2941), .I1(n2867), .CO(n59361));
    SB_LUT4 add_2901_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n59359), 
            .O(n8655[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_18 (.CI(n59359), .I0(n2942), .I1(n2754), .CO(n59360));
    SB_LUT4 add_2901_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n59358), 
            .O(n8655[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_17 (.CI(n59358), .I0(n2943), .I1(n2638), .CO(n59359));
    SB_LUT4 add_2901_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n59357), 
            .O(n8655[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_16 (.CI(n59357), .I0(n2944), .I1(n2519), .CO(n59358));
    SB_LUT4 add_2901_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n59356), 
            .O(n8655[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_15 (.CI(n59356), .I0(n2945), .I1(n2397), .CO(n59357));
    SB_LUT4 add_2901_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n59355), 
            .O(n8655[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_14 (.CI(n59355), .I0(n2946), .I1(n2272), .CO(n59356));
    SB_LUT4 i1_4_lut_adj_1007 (.I0(n9), .I1(n14), .I2(n70817), .I3(baudrate[30]), 
            .O(n25977));
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2901_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n59354), 
            .O(n8655[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_13 (.CI(n59354), .I0(n2947), .I1(n2144), .CO(n59355));
    SB_LUT4 add_2901_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n59353), 
            .O(n8655[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_12 (.CI(n59353), .I0(n2948), .I1(n2013), .CO(n59354));
    SB_LUT4 add_2901_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n59352), 
            .O(n8655[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_11 (.CI(n59352), .I0(n2949), .I1(n1879), .CO(n59353));
    SB_LUT4 add_2901_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n59351), 
            .O(n8655[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_10 (.CI(n59351), .I0(n2950), .I1(n1742), .CO(n59352));
    SB_LUT4 add_2901_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n59350), 
            .O(n8655[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_9 (.CI(n59350), .I0(n2951), .I1(n1602), .CO(n59351));
    SB_LUT4 add_2901_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n59349), 
            .O(n8655[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_8 (.CI(n59349), .I0(n2952), .I1(n1459), .CO(n59350));
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8707[20]), .I3(n294[1]), .O(n41_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8707[19]), .I3(n294[1]), .O(n39_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8707[18]), .I3(n294[1]), .O(n37_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n59348), 
            .O(n8655[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_7 (.CI(n59348), .I0(n2953), .I1(n1460), .CO(n59349));
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8707[11]), .I3(n294[1]), .O(n23_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8707[12]), .I3(n294[1]), .O(n25_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n59347), 
            .O(n8655[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_6 (.CI(n59347), .I0(n2954), .I1(n1011), .CO(n59348));
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8707[14]), .I3(n294[1]), .O(n29_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n59346), 
            .O(n8655[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8707[15]), .I3(n294[1]), .O(n31_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2901_5 (.CI(n59346), .I0(n2955), .I1(n856), .CO(n59347));
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8707[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n59345), 
            .O(n8655[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2901_4 (.CI(n59345), .I0(n2956), .I1(n698), .CO(n59346));
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8707[22]), .I3(n294[1]), .O(n45_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n59344), 
            .O(n8655[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8707[21]), .I3(n294[1]), .O(n43_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2901_3 (.CI(n59344), .I0(n2957), .I1(n858), .CO(n59345));
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8707[4]), .I3(n294[1]), .O(n9_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8707[8]), .I3(n294[1]), .O(n17_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8707[9]), .I3(n294[1]), .O(n19_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2901_2_lut (.I0(n67171), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69409)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2901_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2901_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59344));
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8707[10]), .I3(n294[1]), .O(n21_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8707[17]), .I3(n294[1]), .O(n35_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8707[16]), .I3(n294[1]), .O(n33_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8707[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2900_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n59343), 
            .O(n8629[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2900_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n59342), 
            .O(n8629[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8707[6]), .I3(n294[1]), .O(n13_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8707[7]), .I3(n294[1]), .O(n15_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8707[13]), .I3(n294[1]), .O(n27_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2900_20 (.CI(n59342), .I0(n2828), .I1(n2977), .CO(n59343));
    SB_LUT4 add_2900_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n59341), 
            .O(n8629[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_19 (.CI(n59341), .I0(n2829), .I1(n2867), .CO(n59342));
    SB_LUT4 add_2900_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n59340), 
            .O(n8629[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59406_4_lut (.I0(n27_adj_5215), .I1(n15_adj_5214), .I2(n13_adj_5213), 
            .I3(n11), .O(n75241));
    defparam i59406_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2900_18 (.CI(n59340), .I0(n2830), .I1(n2754), .CO(n59341));
    SB_LUT4 add_2900_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n59339), 
            .O(n8629[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_17 (.CI(n59339), .I0(n2831), .I1(n2638), .CO(n59340));
    SB_LUT4 add_2900_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n59338), 
            .O(n8629[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5212), .I3(GND_net), .O(n12_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59396_2_lut (.I0(n33_adj_5212), .I1(n15_adj_5214), .I2(GND_net), 
            .I3(GND_net), .O(n75231));
    defparam i59396_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5213), .I3(GND_net), .O(n10_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_16 (.CI(n59338), .I0(n2832), .I1(n2519), .CO(n59339));
    SB_LUT4 add_2900_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n59337), 
            .O(n8629[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_15 (.CI(n59337), .I0(n2833), .I1(n2397), .CO(n59338));
    SB_LUT4 add_2900_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n59336), 
            .O(n8629[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5216), .I1(baudrate[17]), 
            .I2(n35_adj_5211), .I3(GND_net), .O(n30_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59424_4_lut (.I0(n21_adj_5210), .I1(n19_adj_5209), .I2(n17_adj_5208), 
            .I3(n9_adj_5207), .O(n75259));
    defparam i59424_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2900_14 (.CI(n59336), .I0(n2834), .I1(n2272), .CO(n59337));
    SB_LUT4 add_2900_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n59335), 
            .O(n8629[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5206), .I3(GND_net), .O(n16_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_13 (.CI(n59335), .I0(n2835), .I1(n2144), .CO(n59336));
    SB_LUT4 add_2900_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n59334), 
            .O(n8629[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59370_2_lut (.I0(n43_adj_5206), .I1(n19_adj_5209), .I2(GND_net), 
            .I3(GND_net), .O(n75205));
    defparam i59370_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2900_12 (.CI(n59334), .I0(n2836), .I1(n2013), .CO(n59335));
    SB_LUT4 add_2900_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n59333), 
            .O(n8629[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_11 (.CI(n59333), .I0(n2837), .I1(n1879), .CO(n59334));
    SB_LUT4 add_2900_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n59332), 
            .O(n8629[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5208), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5219), .I1(baudrate[22]), 
            .I2(n45_adj_5205), .I3(GND_net), .O(n24_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_10 (.CI(n59332), .I0(n2838), .I1(n1742), .CO(n59333));
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8707[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2900_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n59331), 
            .O(n8629[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59446_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n75281));
    defparam i59446_3_lut.LUT_INIT = 16'hbebe;
    SB_CARRY add_2900_9 (.CI(n59331), .I0(n2839), .I1(n1602), .CO(n59332));
    SB_LUT4 i60378_4_lut (.I0(n13_adj_5213), .I1(n11), .I2(n9_adj_5207), 
            .I3(n75281), .O(n76213));
    defparam i60378_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60372_4_lut (.I0(n19_adj_5209), .I1(n17_adj_5208), .I2(n15_adj_5214), 
            .I3(n76213), .O(n76207));
    defparam i60372_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61510_4_lut (.I0(n25_adj_5202), .I1(n23_adj_5201), .I2(n21_adj_5210), 
            .I3(n76207), .O(n77345));
    defparam i61510_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2900_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n59330), 
            .O(n8629[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60865_4_lut (.I0(n31_adj_5204), .I1(n29_adj_5203), .I2(n27_adj_5215), 
            .I3(n77345), .O(n76700));
    defparam i60865_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2900_8 (.CI(n59330), .I0(n2840), .I1(n1459), .CO(n59331));
    SB_LUT4 add_2900_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n59329), 
            .O(n8629[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61656_4_lut (.I0(n37_adj_5200), .I1(n35_adj_5211), .I2(n33_adj_5212), 
            .I3(n76700), .O(n77491));
    defparam i61656_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2900_7 (.CI(n59329), .I0(n2841), .I1(n1460), .CO(n59330));
    SB_LUT4 add_2900_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n59328), 
            .O(n8629[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_6 (.CI(n59328), .I0(n2842), .I1(n1011), .CO(n59329));
    SB_LUT4 add_2900_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n59327), 
            .O(n8629[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2900_5 (.CI(n59327), .I0(n2843), .I1(n856), .CO(n59328));
    SB_LUT4 add_2900_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n59326), 
            .O(n8629[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61059_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21_adj_5210), 
            .I3(GND_net), .O(n76894));   // verilog/uart_rx.v(119[33:55])
    defparam i61059_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_4 (.CI(n59326), .I0(n2844), .I1(n698), .CO(n59327));
    SB_LUT4 add_2900_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n59325), 
            .O(n8629[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i61060_3_lut (.I0(n76894), .I1(baudrate[11]), .I2(n23_adj_5201), 
            .I3(GND_net), .O(n76895));   // verilog/uart_rx.v(119[33:55])
    defparam i61060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n69413), .I3(n48_adj_5221), .O(n4));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i61057_3_lut (.I0(n4), .I1(baudrate[13]), .I2(n27_adj_5215), 
            .I3(GND_net), .O(n76892));   // verilog/uart_rx.v(119[33:55])
    defparam i61057_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_3 (.CI(n59325), .I0(n2845), .I1(n858), .CO(n59326));
    SB_LUT4 add_2900_2_lut (.I0(n67175), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69407)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2900_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i61058_3_lut (.I0(n76892), .I1(baudrate[14]), .I2(n29_adj_5203), 
            .I3(GND_net), .O(n76893));   // verilog/uart_rx.v(119[33:55])
    defparam i61058_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2900_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59325));
    SB_LUT4 add_2899_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n59324), 
            .O(n8603[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2899_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n59323), 
            .O(n8603[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_19 (.CI(n59323), .I0(n2714), .I1(n2867), .CO(n59324));
    SB_LUT4 i59398_4_lut (.I0(n33_adj_5212), .I1(n31_adj_5204), .I2(n29_adj_5203), 
            .I3(n75241), .O(n75233));
    defparam i59398_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2899_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n59322), 
            .O(n8603[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_18 (.CI(n59322), .I0(n2715), .I1(n2754), .CO(n59323));
    SB_LUT4 add_2899_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n59321), 
            .O(n8603[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61540_4_lut (.I0(n30_adj_5218), .I1(n10_adj_5217), .I2(n35_adj_5211), 
            .I3(n75231), .O(n77375));   // verilog/uart_rx.v(119[33:55])
    defparam i61540_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2899_17 (.CI(n59321), .I0(n2716), .I1(n2638), .CO(n59322));
    SB_LUT4 i60166_3_lut (.I0(n76893), .I1(baudrate[15]), .I2(n31_adj_5204), 
            .I3(GND_net), .O(n76001));   // verilog/uart_rx.v(119[33:55])
    defparam i60166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61750_4_lut (.I0(n76001), .I1(n77375), .I2(n35_adj_5211), 
            .I3(n75233), .O(n77585));   // verilog/uart_rx.v(119[33:55])
    defparam i61750_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61751_3_lut (.I0(n77585), .I1(baudrate[18]), .I2(n37_adj_5200), 
            .I3(GND_net), .O(n77586));   // verilog/uart_rx.v(119[33:55])
    defparam i61751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61678_3_lut (.I0(n77586), .I1(baudrate[19]), .I2(n39_adj_5199), 
            .I3(GND_net), .O(n77513));   // verilog/uart_rx.v(119[33:55])
    defparam i61678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8681[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59376_4_lut (.I0(n43_adj_5206), .I1(n25_adj_5202), .I2(n23_adj_5201), 
            .I3(n75259), .O(n75211));
    defparam i59376_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2899_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n59320), 
            .O(n8603[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_16 (.CI(n59320), .I0(n2717), .I1(n2519), .CO(n59321));
    SB_LUT4 i61165_4_lut (.I0(n24_adj_5220), .I1(n8), .I2(n45_adj_5205), 
            .I3(n75205), .O(n77000));   // verilog/uart_rx.v(119[33:55])
    defparam i61165_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2899_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n59319), 
            .O(n8603[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_15 (.CI(n59319), .I0(n2718), .I1(n2397), .CO(n59320));
    SB_LUT4 i60164_3_lut (.I0(n76895), .I1(baudrate[12]), .I2(n25_adj_5202), 
            .I3(GND_net), .O(n75999));   // verilog/uart_rx.v(119[33:55])
    defparam i60164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59378_4_lut (.I0(n43_adj_5206), .I1(n41_adj_5198), .I2(n39_adj_5199), 
            .I3(n77491), .O(n75213));
    defparam i59378_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2899_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n59318), 
            .O(n8603[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_14 (.CI(n59318), .I0(n2719), .I1(n2272), .CO(n59319));
    SB_LUT4 i61598_4_lut (.I0(n75999), .I1(n77000), .I2(n45_adj_5205), 
            .I3(n75211), .O(n77433));   // verilog/uart_rx.v(119[33:55])
    defparam i61598_4_lut.LUT_INIT = 16'hccca;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_5222), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i60172_3_lut (.I0(n77513), .I1(baudrate[20]), .I2(n41_adj_5198), 
            .I3(GND_net), .O(n76007));   // verilog/uart_rx.v(119[33:55])
    defparam i60172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8707[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61600_4_lut (.I0(n76007), .I1(n77433), .I2(n45_adj_5205), 
            .I3(n75213), .O(n77435));   // verilog/uart_rx.v(119[33:55])
    defparam i61600_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2899_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n59317), 
            .O(n8603[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_13 (.CI(n59317), .I0(n2720), .I1(n2144), .CO(n59318));
    SB_LUT4 i62242_4_lut (.I0(n69339), .I1(n77435), .I2(baudrate[23]), 
            .I3(n3253), .O(n68384));   // verilog/uart_rx.v(119[33:55])
    defparam i62242_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 add_2899_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n59316), 
            .O(n8603[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_12 (.CI(n59316), .I0(n2721), .I1(n2013), .CO(n59317));
    SB_LUT4 add_2899_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n59315), 
            .O(n8603[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8681[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2899_11 (.CI(n59315), .I0(n2722), .I1(n1879), .CO(n59316));
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2899_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n59314), 
            .O(n8603[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_10 (.CI(n59314), .I0(n2723), .I1(n1742), .CO(n59315));
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2899_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n59313), 
            .O(n8603[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_9 (.CI(n59313), .I0(n2724), .I1(n1602), .CO(n59314));
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8681[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2899_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n59312), 
            .O(n8603[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_8 (.CI(n59312), .I0(n2725), .I1(n1459), .CO(n59313));
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2899_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n59311), 
            .O(n8603[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2899_7 (.CI(n59311), .I0(n2726), .I1(n1460), .CO(n59312));
    SB_LUT4 add_2899_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n59310), 
            .O(n8603[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2899_6 (.CI(n59310), .I0(n2727), .I1(n1011), .CO(n59311));
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59474_4_lut (.I0(n29_adj_5237), .I1(n17_adj_5236), .I2(n15_adj_5235), 
            .I3(n13_adj_5234), .O(n75309));
    defparam i59474_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60438_4_lut (.I0(n11_adj_5232), .I1(n9_adj_5231), .I2(n3171), 
            .I3(baudrate[2]), .O(n76273));
    defparam i60438_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 add_2899_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n59309), 
            .O(n8603[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60903_4_lut (.I0(n17_adj_5236), .I1(n15_adj_5235), .I2(n13_adj_5234), 
            .I3(n76273), .O(n76738));
    defparam i60903_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60901_4_lut (.I0(n23_adj_5230), .I1(n21_adj_5229), .I2(n19_adj_5233), 
            .I3(n76738), .O(n76736));
    defparam i60901_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59478_4_lut (.I0(n29_adj_5237), .I1(n27_adj_5228), .I2(n25_adj_5227), 
            .I3(n76736), .O(n75313));
    defparam i59478_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2899_5 (.CI(n59309), .I0(n2728), .I1(n856), .CO(n59310));
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2899_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n59308), 
            .O(n8603[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61085_3_lut (.I0(n6_adj_5238), .I1(baudrate[13]), .I2(n29_adj_5237), 
            .I3(GND_net), .O(n76920));   // verilog/uart_rx.v(119[33:55])
    defparam i61085_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2899_4 (.CI(n59308), .I0(n2729), .I1(n698), .CO(n59309));
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5239), .I1(baudrate[17]), 
            .I2(n37_adj_5225), .I3(GND_net), .O(n32_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61086_3_lut (.I0(n76920), .I1(baudrate[14]), .I2(n31_adj_5224), 
            .I3(GND_net), .O(n76921));   // verilog/uart_rx.v(119[33:55])
    defparam i61086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59464_4_lut (.I0(n35_adj_5226), .I1(n33_adj_5223), .I2(n31_adj_5224), 
            .I3(n75309), .O(n75299));
    defparam i59464_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61460_4_lut (.I0(n32_adj_5240), .I1(n12_adj_5241), .I2(n37_adj_5225), 
            .I3(n75295), .O(n77295));   // verilog/uart_rx.v(119[33:55])
    defparam i61460_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60152_3_lut (.I0(n76921), .I1(baudrate[15]), .I2(n33_adj_5223), 
            .I3(GND_net), .O(n75987));   // verilog/uart_rx.v(119[33:55])
    defparam i60152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2899_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n59307), 
            .O(n8603[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2899_3 (.CI(n59307), .I0(n2730), .I1(n858), .CO(n59308));
    SB_LUT4 i61087_3_lut (.I0(n8_adj_5242), .I1(baudrate[10]), .I2(n23_adj_5230), 
            .I3(GND_net), .O(n76922));   // verilog/uart_rx.v(119[33:55])
    defparam i61087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61088_3_lut (.I0(n76922), .I1(baudrate[11]), .I2(n25_adj_5227), 
            .I3(GND_net), .O(n76923));   // verilog/uart_rx.v(119[33:55])
    defparam i61088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2899_2_lut (.I0(n67179), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69405)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2899_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i60420_4_lut (.I0(n25_adj_5227), .I1(n23_adj_5230), .I2(n21_adj_5229), 
            .I3(n75324), .O(n76255));
    defparam i60420_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2899_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59307));
    SB_LUT4 i61163_3_lut (.I0(n10_adj_5243), .I1(baudrate[9]), .I2(n21_adj_5229), 
            .I3(GND_net), .O(n76998));   // verilog/uart_rx.v(119[33:55])
    defparam i61163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2898_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n59306), 
            .O(n8577[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2898_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n59305), 
            .O(n8577[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60150_3_lut (.I0(n76923), .I1(baudrate[12]), .I2(n27_adj_5228), 
            .I3(GND_net), .O(n75985));   // verilog/uart_rx.v(119[33:55])
    defparam i60150_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2898_18 (.CI(n59305), .I0(n2597), .I1(n2754), .CO(n59306));
    SB_LUT4 add_2898_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n59304), 
            .O(n8577[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_17 (.CI(n59304), .I0(n2598), .I1(n2638), .CO(n59305));
    SB_LUT4 add_2898_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n59303), 
            .O(n8577[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61304_4_lut (.I0(n35_adj_5226), .I1(n33_adj_5223), .I2(n31_adj_5224), 
            .I3(n75313), .O(n77139));
    defparam i61304_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2898_16 (.CI(n59303), .I0(n2599), .I1(n2519), .CO(n59304));
    SB_LUT4 add_2898_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n59302), 
            .O(n8577[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61739_4_lut (.I0(n75987), .I1(n77295), .I2(n37_adj_5225), 
            .I3(n75299), .O(n77574));   // verilog/uart_rx.v(119[33:55])
    defparam i61739_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2898_15 (.CI(n59302), .I0(n2600), .I1(n2397), .CO(n59303));
    SB_LUT4 add_2898_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n59301), 
            .O(n8577[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61378_4_lut (.I0(n75985), .I1(n76998), .I2(n27_adj_5228), 
            .I3(n76255), .O(n77213));   // verilog/uart_rx.v(119[33:55])
    defparam i61378_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61812_4_lut (.I0(n77213), .I1(n77574), .I2(n37_adj_5225), 
            .I3(n77139), .O(n77647));   // verilog/uart_rx.v(119[33:55])
    defparam i61812_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2898_14 (.CI(n59301), .I0(n2601), .I1(n2272), .CO(n59302));
    SB_LUT4 add_2898_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n59300), 
            .O(n8577[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61813_3_lut (.I0(n77647), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n77648));   // verilog/uart_rx.v(119[33:55])
    defparam i61813_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2898_13 (.CI(n59300), .I0(n2602), .I1(n2144), .CO(n59301));
    SB_LUT4 i61801_3_lut (.I0(n77648), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n77636));   // verilog/uart_rx.v(119[33:55])
    defparam i61801_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2898_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n59299), 
            .O(n8577[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61572_3_lut (.I0(n77636), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n77407));   // verilog/uart_rx.v(119[33:55])
    defparam i61572_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2898_12 (.CI(n59299), .I0(n2603), .I1(n2013), .CO(n59300));
    SB_LUT4 add_2898_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n59298), 
            .O(n8577[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_11 (.CI(n59298), .I0(n2604), .I1(n1879), .CO(n59299));
    SB_LUT4 add_2898_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n59297), 
            .O(n8577[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_10 (.CI(n59297), .I0(n2605), .I1(n1742), .CO(n59298));
    SB_LUT4 add_2898_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n59296), 
            .O(n8577[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_9 (.CI(n59296), .I0(n2606), .I1(n1602), .CO(n59297));
    SB_LUT4 i61573_3_lut (.I0(n77407), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n77408));   // verilog/uart_rx.v(119[33:55])
    defparam i61573_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2898_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n59295), 
            .O(n8577[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60162_3_lut (.I0(n77408), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam i60162_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2898_8 (.CI(n59295), .I0(n2607), .I1(n1459), .CO(n59296));
    SB_LUT4 add_2898_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n59294), 
            .O(n8577[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_7 (.CI(n59294), .I0(n2608), .I1(n1460), .CO(n59295));
    SB_LUT4 add_2898_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n59293), 
            .O(n8577[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_6 (.CI(n59293), .I0(n2609), .I1(n1011), .CO(n59294));
    SB_LUT4 add_2898_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n59292), 
            .O(n8577[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_5 (.CI(n59292), .I0(n2610), .I1(n856), .CO(n59293));
    SB_LUT4 add_2898_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n59291), 
            .O(n8577[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8681[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2898_4 (.CI(n59291), .I0(n2611), .I1(n698), .CO(n59292));
    SB_LUT4 add_2898_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n59290), 
            .O(n8577[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2898_3 (.CI(n59290), .I0(n2612), .I1(n858), .CO(n59291));
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8681[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2898_2_lut (.I0(n67183), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69403)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2898_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2898_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59290));
    SB_LUT4 add_2897_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n59289), 
            .O(n8551[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2897_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n59288), 
            .O(n8551[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_17 (.CI(n59288), .I0(n2477), .I1(n2638), .CO(n59289));
    SB_LUT4 add_2897_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n59287), 
            .O(n8551[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_16 (.CI(n59287), .I0(n2478), .I1(n2519), .CO(n59288));
    SB_LUT4 add_2897_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n59286), 
            .O(n8551[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_15 (.CI(n59286), .I0(n2479), .I1(n2397), .CO(n59287));
    SB_LUT4 add_2897_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n59285), 
            .O(n8551[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_14 (.CI(n59285), .I0(n2480), .I1(n2272), .CO(n59286));
    SB_LUT4 add_2897_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n59284), 
            .O(n8551[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_13 (.CI(n59284), .I0(n2481), .I1(n2144), .CO(n59285));
    SB_LUT4 add_2897_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n59283), 
            .O(n8551[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8681[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2897_12 (.CI(n59283), .I0(n2482), .I1(n2013), .CO(n59284));
    SB_LUT4 add_2897_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n59282), 
            .O(n8551[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8681[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2897_11 (.CI(n59282), .I0(n2483), .I1(n1879), .CO(n59283));
    SB_LUT4 add_2897_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n59281), 
            .O(n8551[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_10 (.CI(n59281), .I0(n2484), .I1(n1742), .CO(n59282));
    SB_LUT4 add_2897_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n59280), 
            .O(n8551[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_9 (.CI(n59280), .I0(n2485), .I1(n1602), .CO(n59281));
    SB_LUT4 add_2897_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n59279), 
            .O(n8551[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_8 (.CI(n59279), .I0(n2486), .I1(n1459), .CO(n59280));
    SB_LUT4 add_2897_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n59278), 
            .O(n8551[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_7 (.CI(n59278), .I0(n2487), .I1(n1460), .CO(n59279));
    SB_LUT4 add_2897_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n59277), 
            .O(n8551[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_6 (.CI(n59277), .I0(n2488), .I1(n1011), .CO(n59278));
    SB_LUT4 add_2897_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n59276), 
            .O(n8551[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_5 (.CI(n59276), .I0(n2489), .I1(n856), .CO(n59277));
    SB_LUT4 add_2897_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n59275), 
            .O(n8551[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_4 (.CI(n59275), .I0(n2490), .I1(n698), .CO(n59276));
    SB_LUT4 add_2897_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n59274), 
            .O(n8551[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2897_3 (.CI(n59274), .I0(n2491), .I1(n858), .CO(n59275));
    SB_LUT4 add_2897_2_lut (.I0(n67187), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69401)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2897_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2897_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59274));
    SB_LUT4 add_2896_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n59273), 
            .O(n8525[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2896_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n59272), 
            .O(n8525[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_16 (.CI(n59272), .I0(n2354), .I1(n2519), .CO(n59273));
    SB_LUT4 add_2896_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n59271), 
            .O(n8525[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_15 (.CI(n59271), .I0(n2355), .I1(n2397), .CO(n59272));
    SB_LUT4 add_2896_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n59270), 
            .O(n8525[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_14 (.CI(n59270), .I0(n2356), .I1(n2272), .CO(n59271));
    SB_LUT4 add_2896_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n59269), 
            .O(n8525[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_13 (.CI(n59269), .I0(n2357), .I1(n2144), .CO(n59270));
    SB_LUT4 add_2896_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n59268), 
            .O(n8525[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_12 (.CI(n59268), .I0(n2358), .I1(n2013), .CO(n59269));
    SB_LUT4 add_2896_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n59267), 
            .O(n8525[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_11 (.CI(n59267), .I0(n2359), .I1(n1879), .CO(n59268));
    SB_LUT4 add_2896_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n59266), 
            .O(n8525[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_10 (.CI(n59266), .I0(n2360), .I1(n1742), .CO(n59267));
    SB_LUT4 add_2896_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n59265), 
            .O(n8525[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_9 (.CI(n59265), .I0(n2361), .I1(n1602), .CO(n59266));
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2896_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n59264), 
            .O(n8525[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_8 (.CI(n59264), .I0(n2362), .I1(n1459), .CO(n59265));
    SB_LUT4 add_2896_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n59263), 
            .O(n8525[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_7 (.CI(n59263), .I0(n2363), .I1(n1460), .CO(n59264));
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8681[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2896_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n59262), 
            .O(n8525[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_6 (.CI(n59262), .I0(n2364), .I1(n1011), .CO(n59263));
    SB_LUT4 add_2896_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n59261), 
            .O(n8525[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_5 (.CI(n59261), .I0(n2365), .I1(n856), .CO(n59262));
    SB_LUT4 add_2896_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n59260), 
            .O(n8525[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_4 (.CI(n59260), .I0(n2366), .I1(n698), .CO(n59261));
    SB_LUT4 add_2896_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n59259), 
            .O(n8525[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2896_3 (.CI(n59259), .I0(n2367), .I1(n858), .CO(n59260));
    SB_LUT4 i55735_1_lut (.I0(n71560), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67221));
    defparam i55735_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2896_2_lut (.I0(n67191), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69399)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2896_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2896_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59259));
    SB_LUT4 add_2895_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n59258), 
            .O(n8499[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2895_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n59257), 
            .O(n8499[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n58290), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_15 (.CI(n59257), .I0(n2228), .I1(n2397), .CO(n59258));
    SB_LUT4 add_2895_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n59256), 
            .O(n8499[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_14 (.CI(n59256), .I0(n2229), .I1(n2272), .CO(n59257));
    SB_LUT4 add_2895_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n59255), 
            .O(n8499[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_13 (.CI(n59255), .I0(n2230), .I1(n2144), .CO(n59256));
    SB_LUT4 add_2895_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n59254), 
            .O(n8499[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n69351), .I1(n294[23]), .I2(VCC_net), 
            .I3(n58289), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2895_12 (.CI(n59254), .I0(n2231), .I1(n2013), .CO(n59255));
    SB_LUT4 add_2895_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n59253), 
            .O(n8499[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_25 (.CI(n58289), .I0(n294[23]), .I1(VCC_net), 
            .CO(n58290));
    SB_CARRY add_2895_11 (.CI(n59253), .I0(n2232), .I1(n1879), .CO(n59254));
    SB_LUT4 add_2895_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n59252), 
            .O(n8499[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_10 (.CI(n59252), .I0(n2233), .I1(n1742), .CO(n59253));
    SB_LUT4 add_2895_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n59251), 
            .O(n8499[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_9 (.CI(n59251), .I0(n2234), .I1(n1602), .CO(n59252));
    SB_LUT4 add_2895_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n59250), 
            .O(n8499[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n69453), .I1(n71578), .I2(VCC_net), 
            .I3(n58288), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2895_8 (.CI(n59250), .I0(n2235), .I1(n1459), .CO(n59251));
    SB_LUT4 add_2895_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n59249), 
            .O(n8499[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_7 (.CI(n59249), .I0(n2236), .I1(n1460), .CO(n59250));
    SB_LUT4 add_2895_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n59248), 
            .O(n8499[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59784_2_lut (.I0(n65798), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n74542));
    defparam i59784_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2895_6 (.CI(n59248), .I0(n2237), .I1(n1011), .CO(n59249));
    SB_LUT4 i59773_4_lut (.I0(n74542), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n74539));
    defparam i59773_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2895_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n59247), 
            .O(n8499[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2895_5 (.CI(n59247), .I0(n2238), .I1(n856), .CO(n59248));
    SB_LUT4 add_2895_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n59246), 
            .O(n8499[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_24 (.CI(n58288), .I0(n71578), .I1(VCC_net), 
            .CO(n58289));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n58287), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i59087_4_lut (.I0(n74539), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n74536));
    defparam i59087_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i62326_4_lut (.I0(\r_SM_Main[2] ), .I1(n74536), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(\r_SM_Main[1] ), .O(n29421));
    defparam i62326_4_lut.LUT_INIT = 16'h0511;
    SB_CARRY sub_38_add_2_23 (.CI(n58287), .I0(n294[21]), .I1(VCC_net), 
            .CO(n58288));
    SB_CARRY add_2895_4 (.CI(n59246), .I0(n2239), .I1(n698), .CO(n59247));
    SB_LUT4 add_2895_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n59245), 
            .O(n8499[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(n65798), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n69477));
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n69477), .O(n69483));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'h0100;
    SB_CARRY add_2895_3 (.CI(n59245), .I0(n2240), .I1(n858), .CO(n59246));
    SB_LUT4 add_2895_2_lut (.I0(n67195), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69397)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2895_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2895_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59245));
    SB_LUT4 add_2894_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n59244), 
            .O(n8473[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61885_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n69483), .O(n28159));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i61885_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 add_2894_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n59243), 
            .O(n8473[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_13 (.CI(n59243), .I0(n2099), .I1(n2272), .CO(n59244));
    SB_LUT4 add_2894_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n59242), 
            .O(n8473[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_22_lut (.I0(n69451), .I1(n294[20]), .I2(VCC_net), 
            .I3(n58286), .O(n69453)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2894_12 (.CI(n59242), .I0(n2100), .I1(n2144), .CO(n59243));
    SB_CARRY sub_38_add_2_22 (.CI(n58286), .I0(n294[20]), .I1(VCC_net), 
            .CO(n58287));
    SB_LUT4 add_2894_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n59241), 
            .O(n8473[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_11 (.CI(n59241), .I0(n2101), .I1(n2013), .CO(n59242));
    SB_LUT4 add_2894_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n59240), 
            .O(n8473[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n69449), .I1(n294[19]), .I2(VCC_net), 
            .I3(n58285), .O(n69451)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2894_10 (.CI(n59240), .I0(n2102), .I1(n1879), .CO(n59241));
    SB_LUT4 add_2894_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n59239), 
            .O(n8473[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_21 (.CI(n58285), .I0(n294[19]), .I1(VCC_net), 
            .CO(n58286));
    SB_CARRY add_2894_9 (.CI(n59239), .I0(n2103), .I1(n1742), .CO(n59240));
    SB_LUT4 add_2894_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n59238), 
            .O(n8473[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_8 (.CI(n59238), .I0(n2104), .I1(n1602), .CO(n59239));
    SB_LUT4 add_2894_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n59237), 
            .O(n8473[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_7 (.CI(n59237), .I0(n2105), .I1(n1459), .CO(n59238));
    SB_LUT4 add_2894_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n59236), 
            .O(n8473[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_6 (.CI(n59236), .I0(n2106), .I1(n1460), .CO(n59237));
    SB_LUT4 add_2894_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n59235), 
            .O(n8473[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_5 (.CI(n59235), .I0(n2107), .I1(n1011), .CO(n59236));
    SB_LUT4 add_2894_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n59234), 
            .O(n8473[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_4 (.CI(n59234), .I0(n2108), .I1(n856), .CO(n59235));
    SB_LUT4 add_2894_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n59233), 
            .O(n8473[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n58284), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i55734_2_lut_3_lut_4_lut (.I0(baudrate[9]), .I1(n71554), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n71560));
    defparam i55734_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2894_3 (.CI(n59233), .I0(n2109), .I1(n698), .CO(n59234));
    SB_LUT4 add_2894_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8473[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2894_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2894_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n59233));
    SB_LUT4 add_2893_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n59232), 
            .O(n8447[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2893_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n59231), 
            .O(n8447[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_13 (.CI(n59231), .I0(n1967), .I1(n2144), .CO(n59232));
    SB_LUT4 add_2893_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n59230), 
            .O(n8447[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_12 (.CI(n59230), .I0(n1968), .I1(n2013), .CO(n59231));
    SB_LUT4 add_2893_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n59229), 
            .O(n8447[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_11 (.CI(n59229), .I0(n1969), .I1(n1879), .CO(n59230));
    SB_LUT4 add_2893_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n59228), 
            .O(n8447[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_10 (.CI(n59228), .I0(n1970), .I1(n1742), .CO(n59229));
    SB_LUT4 add_2893_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n59227), 
            .O(n8447[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_9 (.CI(n59227), .I0(n1971), .I1(n1602), .CO(n59228));
    SB_LUT4 add_2893_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n59226), 
            .O(n8447[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_8 (.CI(n59226), .I0(n1972), .I1(n1459), .CO(n59227));
    SB_CARRY sub_38_add_2_20 (.CI(n58284), .I0(n294[18]), .I1(VCC_net), 
            .CO(n58285));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n69447), .I1(n294[17]), .I2(VCC_net), 
            .I3(n58283), .O(n69449)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2893_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n59225), 
            .O(n8447[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_7 (.CI(n59225), .I0(n1973), .I1(n1460), .CO(n59226));
    SB_LUT4 add_2893_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n59224), 
            .O(n8447[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_6 (.CI(n59224), .I0(n1974), .I1(n1011), .CO(n59225));
    SB_CARRY sub_38_add_2_19 (.CI(n58283), .I0(n294[17]), .I1(VCC_net), 
            .CO(n58284));
    SB_LUT4 add_2893_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n59223), 
            .O(n8447[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_5 (.CI(n59223), .I0(n1975), .I1(n856), .CO(n59224));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n69445), .I1(n294[16]), .I2(VCC_net), 
            .I3(n58282), .O(n69447)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2893_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n59222), 
            .O(n8447[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_4 (.CI(n59222), .I0(n1976), .I1(n698), .CO(n59223));
    SB_LUT4 add_2893_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n59221), 
            .O(n8447[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2893_3 (.CI(n59221), .I0(n1977), .I1(n858), .CO(n59222));
    SB_LUT4 add_2893_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8447[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2893_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_18 (.CI(n58282), .I0(n294[16]), .I1(VCC_net), 
            .CO(n58283));
    SB_CARRY add_2893_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59221));
    SB_LUT4 sub_38_add_2_17_lut (.I0(n69349), .I1(n294[15]), .I2(VCC_net), 
            .I3(n58281), .O(n69351)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2892_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n59220), 
            .O(n8421[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2892_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n59219), 
            .O(n8421[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_12 (.CI(n59219), .I0(n1832), .I1(n2013), .CO(n59220));
    SB_LUT4 add_2892_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n59218), 
            .O(n8421[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_17 (.CI(n58281), .I0(n294[15]), .I1(VCC_net), 
            .CO(n58282));
    SB_CARRY add_2892_11 (.CI(n59218), .I0(n1833), .I1(n1879), .CO(n59219));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n69443), .I1(n294[14]), .I2(VCC_net), 
            .I3(n58280), .O(n69445)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n58280), .I0(n294[14]), .I1(VCC_net), 
            .CO(n58281));
    SB_LUT4 add_2892_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n59217), 
            .O(n8421[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_10 (.CI(n59217), .I0(n1834), .I1(n1742), .CO(n59218));
    SB_LUT4 add_2892_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n59216), 
            .O(n8421[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_9 (.CI(n59216), .I0(n1835), .I1(n1602), .CO(n59217));
    SB_LUT4 add_2892_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n59215), 
            .O(n8421[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_8 (.CI(n59215), .I0(n1836), .I1(n1459), .CO(n59216));
    SB_LUT4 add_2892_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n59214), 
            .O(n8421[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n58279), .O(n69443)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2892_7 (.CI(n59214), .I0(n1837), .I1(n1460), .CO(n59215));
    SB_CARRY sub_38_add_2_15 (.CI(n58279), .I0(n294[13]), .I1(VCC_net), 
            .CO(n58280));
    SB_LUT4 add_2892_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n59213), 
            .O(n8421[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n58278), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_6 (.CI(n59213), .I0(n1838), .I1(n1011), .CO(n59214));
    SB_LUT4 add_2892_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n59212), 
            .O(n8421[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_5 (.CI(n59212), .I0(n1839), .I1(n856), .CO(n59213));
    SB_LUT4 add_2892_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n59211), 
            .O(n8421[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_4 (.CI(n59211), .I0(n1840), .I1(n698), .CO(n59212));
    SB_CARRY sub_38_add_2_14 (.CI(n58278), .I0(n294[12]), .I1(VCC_net), 
            .CO(n58279));
    SB_LUT4 add_2892_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n59210), 
            .O(n8421[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2892_3 (.CI(n59210), .I0(n1841), .I1(n858), .CO(n59211));
    SB_LUT4 add_2892_2_lut (.I0(n67204), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69395)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2892_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n58277), .O(n69349)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2892_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59210));
    SB_LUT4 add_2891_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n59209), 
            .O(n8395[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2891_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n59208), 
            .O(n8395[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_13 (.CI(n58277), .I0(n294[11]), .I1(VCC_net), 
            .CO(n58278));
    SB_CARRY add_2891_10 (.CI(n59208), .I0(n1694), .I1(n1879), .CO(n59209));
    SB_LUT4 add_2891_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n59207), 
            .O(n8395[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n58276), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_9 (.CI(n59207), .I0(n1695), .I1(n1742), .CO(n59208));
    SB_LUT4 add_2891_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n59206), 
            .O(n8395[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_8 (.CI(n59206), .I0(n1696), .I1(n1602), .CO(n59207));
    SB_LUT4 add_2891_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n59205), 
            .O(n8395[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_7 (.CI(n59205), .I0(n1697), .I1(n1459), .CO(n59206));
    SB_LUT4 add_2891_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n59204), 
            .O(n8395[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_6 (.CI(n59204), .I0(n1698), .I1(n1460), .CO(n59205));
    SB_LUT4 add_2891_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n59203), 
            .O(n8395[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n58276), .I0(n294[10]), .I1(VCC_net), 
            .CO(n58277));
    SB_CARRY add_2891_5 (.CI(n59203), .I0(n1699), .I1(n1011), .CO(n59204));
    SB_LUT4 add_2891_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n59202), 
            .O(n8395[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_4 (.CI(n59202), .I0(n1700), .I1(n856), .CO(n59203));
    SB_LUT4 add_2891_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n59201), 
            .O(n8395[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_3 (.CI(n59201), .I0(n1701), .I1(n698), .CO(n59202));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n58275), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n58275), .I0(n294[9]), .I1(VCC_net), 
            .CO(n58276));
    SB_LUT4 add_2891_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8395[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2891_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2891_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n59201));
    SB_LUT4 add_2890_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n59200), 
            .O(n8369[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2890_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n59199), 
            .O(n8369[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_10 (.CI(n59199), .I0(n1553), .I1(n1742), .CO(n59200));
    SB_LUT4 add_2890_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n59198), 
            .O(n8369[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n58274), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_9 (.CI(n59198), .I0(n1554), .I1(n1602), .CO(n59199));
    SB_CARRY sub_38_add_2_10 (.CI(n58274), .I0(n294[8]), .I1(VCC_net), 
            .CO(n58275));
    SB_LUT4 add_2890_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n59197), 
            .O(n8369[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5837_2_lut_3_lut_4_lut (.I0(baudrate[3]), .I1(n21187), .I2(n11690), 
            .I3(n960), .O(n44_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam i5837_2_lut_3_lut_4_lut.LUT_INIT = 16'hfd54;
    SB_CARRY add_2890_8 (.CI(n59197), .I0(n1555), .I1(n1459), .CO(n59198));
    SB_LUT4 add_2890_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n59196), 
            .O(n8369[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_7 (.CI(n59196), .I0(n1556), .I1(n1460), .CO(n59197));
    SB_LUT4 add_2890_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n59195), 
            .O(n8369[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_6 (.CI(n59195), .I0(n1557), .I1(n1011), .CO(n59196));
    SB_LUT4 add_2890_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n59194), 
            .O(n8369[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_5 (.CI(n59194), .I0(n1558), .I1(n856), .CO(n59195));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n58273), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2890_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n59193), 
            .O(n8369[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_4 (.CI(n59193), .I0(n1559), .I1(n698), .CO(n59194));
    SB_LUT4 add_2890_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n59192), 
            .O(n8369[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_3 (.CI(n59192), .I0(n1560), .I1(n858), .CO(n59193));
    SB_LUT4 add_2890_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8369[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2890_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2890_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59192));
    SB_LUT4 add_2889_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n59191), 
            .O(n8343[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2889_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n59190), 
            .O(n8343[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_9 (.CI(n59190), .I0(n1409), .I1(n1602), .CO(n59191));
    SB_LUT4 add_2889_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n59189), 
            .O(n8343[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_8 (.CI(n59189), .I0(n1410), .I1(n1459), .CO(n59190));
    SB_LUT4 add_2889_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n59188), 
            .O(n8343[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_7 (.CI(n59188), .I0(n1411), .I1(n1460), .CO(n59189));
    SB_LUT4 add_2889_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n59187), 
            .O(n8343[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_6 (.CI(n59187), .I0(n1412), .I1(n1011), .CO(n59188));
    SB_LUT4 add_2889_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n59186), 
            .O(n8343[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_5 (.CI(n59186), .I0(n1413), .I1(n856), .CO(n59187));
    SB_LUT4 add_2889_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n59185), 
            .O(n8343[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_4 (.CI(n59185), .I0(n1414), .I1(n698), .CO(n59186));
    SB_LUT4 add_2889_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n59184), 
            .O(n8343[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2889_3 (.CI(n59184), .I0(n1415), .I1(n858), .CO(n59185));
    SB_LUT4 add_2889_2_lut (.I0(n67213), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69393)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2889_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2889_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59184));
    SB_LUT4 add_2888_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n59183), 
            .O(n8317[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2888_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n59182), 
            .O(n8317[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_8 (.CI(n59182), .I0(n1262), .I1(n1459), .CO(n59183));
    SB_LUT4 add_2888_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n59181), 
            .O(n8317[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_7 (.CI(n59181), .I0(n1263), .I1(n1460), .CO(n59182));
    SB_LUT4 add_2888_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n59180), 
            .O(n8317[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_6 (.CI(n59180), .I0(n1264), .I1(n1011), .CO(n59181));
    SB_LUT4 add_2888_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n59179), 
            .O(n8317[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5666_2_lut_3_lut_4_lut (.I0(baudrate[2]), .I1(n21177), .I2(n44716), 
            .I3(n804), .O(n44_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam i5666_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf45;
    SB_CARRY add_2888_5 (.CI(n59179), .I0(n1265), .I1(n856), .CO(n59180));
    SB_LUT4 add_2888_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n59178), 
            .O(n8317[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n58273), .I0(n294[7]), .I1(VCC_net), 
            .CO(n58274));
    SB_CARRY add_2888_4 (.CI(n59178), .I0(n1266), .I1(n698), .CO(n59179));
    SB_LUT4 add_2888_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n59177), 
            .O(n8317[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2888_3 (.CI(n59177), .I0(n1267), .I1(n858), .CO(n59178));
    SB_LUT4 add_2888_2_lut (.I0(n67217), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69391)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2888_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2888_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59177));
    SB_LUT4 add_2887_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n59176), 
            .O(n8291[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2887_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n59175), 
            .O(n8291[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_7 (.CI(n59175), .I0(n1112), .I1(n1460), .CO(n59176));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n58272), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2887_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n59174), 
            .O(n8291[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_6 (.CI(n59174), .I0(n1113), .I1(n1011), .CO(n59175));
    SB_CARRY sub_38_add_2_8 (.CI(n58272), .I0(n294[6]), .I1(VCC_net), 
            .CO(n58273));
    SB_LUT4 add_2887_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n59173), 
            .O(n8291[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_5 (.CI(n59173), .I0(n1114), .I1(n856), .CO(n59174));
    SB_LUT4 add_2887_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n59172), 
            .O(n8291[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_4 (.CI(n59172), .I0(n1115), .I1(n698), .CO(n59173));
    SB_LUT4 add_2887_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n59171), 
            .O(n8291[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2887_3 (.CI(n59171), .I0(n1116), .I1(n858), .CO(n59172));
    SB_LUT4 add_2887_2_lut (.I0(n67221), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n69389)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2887_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2887_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n59171));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n58271), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n58271), .I0(n294[5]), .I1(VCC_net), 
            .CO(n58272));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n58270), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n58270), .I0(n294[4]), .I1(VCC_net), 
            .CO(n58271));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n58269), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n58269), .I0(n294[3]), .I1(VCC_net), 
            .CO(n58270));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n58268), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n58268), .I0(n294[2]), .I1(VCC_net), 
            .CO(n58269));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n58267), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n58267), .I0(n294[1]), .I1(VCC_net), 
            .CO(n58268));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n68384), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n68384), .I1(GND_net), 
            .CO(n58267));
    SB_LUT4 i61882_2_lut_3_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n28238));
    defparam i61882_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 r_Clock_Count_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n59549), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n59548), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_8 (.CI(n59548), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n59549));
    SB_LUT4 r_Clock_Count_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n59547), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_7 (.CI(n59547), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n59548));
    SB_LUT4 r_Clock_Count_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n59546), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_6 (.CI(n59546), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n59547));
    SB_LUT4 r_Clock_Count_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n59545), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_5 (.CI(n59545), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n59546));
    SB_LUT4 r_Clock_Count_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n59544), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_4 (.CI(n59544), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n59545));
    SB_LUT4 r_Clock_Count_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n59543), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_3 (.CI(n59543), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n59544));
    SB_LUT4 r_Clock_Count_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n59543));
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\r_SM_Main[1] ), .I1(\r_SM_Main[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n66050));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5246));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5215), 
            .O(n15_adj_5247));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5247), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5246), 
            .I3(n66050), .O(n79053));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_adj_1011 (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[2] ), .I3(GND_net), .O(n4_adj_5248));
    defparam i1_2_lut_3_lut_adj_1011.LUT_INIT = 16'hfdfd;
    SB_LUT4 i55733_1_lut_2_lut_3_lut (.I0(baudrate[9]), .I1(n71554), .I2(baudrate[8]), 
            .I3(GND_net), .O(n67217));
    defparam i55733_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i59122_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n74957));   // verilog/uart_rx.v(119[33:55])
    defparam i59122_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i55744_2_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(n71560), 
            .I3(GND_net), .O(n71570));
    defparam i55744_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1012 (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(baudrate[4]), .I3(baudrate[3]), .O(n69875));
    defparam i1_2_lut_3_lut_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i62650_2_lut_4_lut (.I0(n77408), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25977), .O(n294[1]));
    defparam i62650_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i62397_4_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_5249), .I3(n69006), .O(n67079));
    defparam i62397_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i55748_3_lut_4_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(baudrate[2]), 
            .I3(n71570), .O(n71574));
    defparam i55748_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59460_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n75295));
    defparam i59460_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59489_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n75324));
    defparam i59489_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1013 (.I0(baudrate[28]), .I1(baudrate[27]), 
            .I2(n14), .I3(n70801), .O(n69339));
    defparam i1_3_lut_4_lut_adj_1013.LUT_INIT = 16'hfffe;
    SB_LUT4 i51376_1_lut_4_lut (.I0(n9), .I1(n14), .I2(n70817), .I3(baudrate[30]), 
            .O(n67163));
    defparam i51376_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_3_lut_4_lut_adj_1014 (.I0(baudrate[2]), .I1(n42_adj_5250), 
            .I2(baudrate[3]), .I3(n21179), .O(n67659));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1014.LUT_INIT = 16'hff4f;
    SB_LUT4 i1_3_lut_4_lut_adj_1015 (.I0(baudrate[3]), .I1(n42_adj_5251), 
            .I2(baudrate[4]), .I3(n21189), .O(n67643));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1015.LUT_INIT = 16'hff4f;
    SB_LUT4 i1_2_lut_4_lut (.I0(n77085), .I1(baudrate[6]), .I2(n1111), 
            .I3(n69389), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i62589_2_lut_4_lut (.I0(n77085), .I1(baudrate[6]), .I2(n1111), 
            .I3(n71560), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i62589_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59143_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n74978));   // verilog/uart_rx.v(119[33:55])
    defparam i59143_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i59068_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n74903));   // verilog/uart_rx.v(119[33:55])
    defparam i59068_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1016 (.I0(n77428), .I1(baudrate[16]), .I2(n2476), 
            .I3(n69401), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1016.LUT_INIT = 16'h7100;
    SB_LUT4 i62616_2_lut_4_lut (.I0(n77428), .I1(baudrate[16]), .I2(n2476), 
            .I3(n26017), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i62616_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8681[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8681[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1017 (.I0(n77041), .I1(baudrate[21]), .I2(n3046), 
            .I3(n69411), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1017.LUT_INIT = 16'h7100;
    SB_LUT4 i62647_2_lut_4_lut (.I0(n77041), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25974), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i62647_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1018 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[31]), .I3(baudrate[30]), .O(n70809));
    defparam i1_2_lut_4_lut_adj_1018.LUT_INIT = 16'hfffe;
    SB_LUT4 i51396_1_lut (.I0(n25935), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67183));
    defparam i51396_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8681[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8681[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8681[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8681[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51392_1_lut (.I0(n25965), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67179));
    defparam i51392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8681[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8681[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8681[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5659_2_lut_4_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam i5659_2_lut_4_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8681[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1019 (.I0(n77640), .I1(baudrate[20]), .I2(n2938), 
            .I3(n69409), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1019.LUT_INIT = 16'h7100;
    SB_LUT4 i62641_2_lut_4_lut (.I0(n77640), .I1(baudrate[20]), .I2(n2938), 
            .I3(n25971), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i62641_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8681[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59613_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n75448));
    defparam i59613_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8681[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8655[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8655[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8655[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8655[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8655[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8655[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8655[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59584_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n75419));
    defparam i59584_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8655[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8655[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8655[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8655[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1020 (.I0(baudrate[31]), .I1(baudrate[23]), 
            .I2(baudrate[21]), .I3(GND_net), .O(n70821));
    defparam i1_2_lut_3_lut_adj_1020.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8655[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59582_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5215), .I3(\o_Rx_DV_N_3488[8] ), .O(n74551));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i59582_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59714_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n65798), 
            .I3(r_SM_Main[0]), .O(n74557));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i59714_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i59579_4_lut (.I0(n74551), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n74548));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i59579_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i59589_4_lut (.I0(n74557), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n74554));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i59589_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n74554), .I1(n74548), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_5222));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8655[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8655[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8655[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8655[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8655[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8655[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8655[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59672_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n75507));
    defparam i59672_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59531_4_lut (.I0(n31_adj_5263), .I1(n19_adj_5268), .I2(n17_adj_5267), 
            .I3(n15_adj_5266), .O(n75366));
    defparam i59531_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60494_4_lut (.I0(n13_adj_5264), .I1(n11_adj_5262), .I2(n3065), 
            .I3(baudrate[2]), .O(n76329));
    defparam i60494_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60933_4_lut (.I0(n19_adj_5268), .I1(n17_adj_5267), .I2(n15_adj_5266), 
            .I3(n76329), .O(n76768));
    defparam i60933_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60929_4_lut (.I0(n25_adj_5259), .I1(n23_adj_5258), .I2(n21_adj_5265), 
            .I3(n76768), .O(n76764));
    defparam i60929_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59533_4_lut (.I0(n31_adj_5263), .I1(n29_adj_5261), .I2(n27_adj_5260), 
            .I3(n76764), .O(n75368));
    defparam i59533_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61095_3_lut (.I0(n8_adj_5269), .I1(baudrate[13]), .I2(n31_adj_5263), 
            .I3(GND_net), .O(n76930));   // verilog/uart_rx.v(119[33:55])
    defparam i61095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59633_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n75468));
    defparam i59633_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61096_3_lut (.I0(n76930), .I1(baudrate[14]), .I2(n33_adj_5256), 
            .I3(GND_net), .O(n76931));   // verilog/uart_rx.v(119[33:55])
    defparam i61096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1021 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69649));
    defparam i1_3_lut_4_lut_adj_1021.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_3_lut_4_lut_adj_1022 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69585));
    defparam i1_3_lut_4_lut_adj_1022.LUT_INIT = 16'hff7f;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5183), .I1(baudrate[17]), 
            .I2(n39_adj_5255), .I3(GND_net), .O(n34_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59525_4_lut (.I0(n37_adj_5257), .I1(n35_adj_5254), .I2(n33_adj_5256), 
            .I3(n75366), .O(n75360));
    defparam i59525_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61458_4_lut (.I0(n34_adj_5270), .I1(n14_adj_5182), .I2(n39_adj_5255), 
            .I3(n75356), .O(n77293));   // verilog/uart_rx.v(119[33:55])
    defparam i61458_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_adj_1023 (.I0(baudrate[22]), .I1(baudrate[23]), 
            .I2(baudrate[31]), .I3(baudrate[30]), .O(n70767));
    defparam i1_2_lut_4_lut_adj_1023.LUT_INIT = 16'hfffe;
    SB_LUT4 i60140_3_lut (.I0(n76931), .I1(baudrate[15]), .I2(n35_adj_5254), 
            .I3(GND_net), .O(n75975));   // verilog/uart_rx.v(119[33:55])
    defparam i60140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1024 (.I0(n77634), .I1(baudrate[19]), .I2(n2827), 
            .I3(n69407), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1024.LUT_INIT = 16'h7100;
    SB_LUT4 i1_3_lut_4_lut_adj_1025 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69665));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1025.LUT_INIT = 16'hffbf;
    SB_LUT4 i61097_3_lut (.I0(n10_adj_5181), .I1(baudrate[10]), .I2(n25_adj_5259), 
            .I3(GND_net), .O(n76932));   // verilog/uart_rx.v(119[33:55])
    defparam i61097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61098_3_lut (.I0(n76932), .I1(baudrate[11]), .I2(n27_adj_5260), 
            .I3(GND_net), .O(n76933));   // verilog/uart_rx.v(119[33:55])
    defparam i61098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1026 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69633));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1026.LUT_INIT = 16'hfffb;
    SB_LUT4 i60470_4_lut (.I0(n27_adj_5260), .I1(n25_adj_5259), .I2(n23_adj_5258), 
            .I3(n75382), .O(n76305));
    defparam i60470_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5184), .I1(baudrate[9]), 
            .I2(n23_adj_5258), .I3(GND_net), .O(n20_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1027 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69601));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1027.LUT_INIT = 16'hfffd;
    SB_LUT4 i62636_2_lut_4_lut (.I0(n77634), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25968), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i62636_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i60138_3_lut (.I0(n76933), .I1(baudrate[12]), .I2(n29_adj_5261), 
            .I3(GND_net), .O(n75973));   // verilog/uart_rx.v(119[33:55])
    defparam i60138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61316_4_lut (.I0(n37_adj_5257), .I1(n35_adj_5254), .I2(n33_adj_5256), 
            .I3(n75368), .O(n77151));
    defparam i61316_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61727_4_lut (.I0(n75975), .I1(n77293), .I2(n39_adj_5255), 
            .I3(n75360), .O(n77562));   // verilog/uart_rx.v(119[33:55])
    defparam i61727_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_4_lut_adj_1028 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69617));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1028.LUT_INIT = 16'hffdf;
    SB_LUT4 i61159_4_lut (.I0(n75973), .I1(n20_adj_5271), .I2(n29_adj_5261), 
            .I3(n76305), .O(n76994));   // verilog/uart_rx.v(119[33:55])
    defparam i61159_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61796_4_lut (.I0(n76994), .I1(n77562), .I2(n39_adj_5255), 
            .I3(n77151), .O(n77631));   // verilog/uart_rx.v(119[33:55])
    defparam i61796_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61797_3_lut (.I0(n77631), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n77632));   // verilog/uart_rx.v(119[33:55])
    defparam i61797_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61205_3_lut (.I0(n77632), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n77040));   // verilog/uart_rx.v(119[33:55])
    defparam i61205_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61206_3_lut (.I0(n77040), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n77041));   // verilog/uart_rx.v(119[33:55])
    defparam i61206_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1029 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69697));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1029.LUT_INIT = 16'hffef;
    SB_LUT4 i1_3_lut_4_lut_adj_1030 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4_adj_5248), .O(n69681));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8629[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59740_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n75575));
    defparam i59740_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8629[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8629[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8629[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59697_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n75532));
    defparam i59697_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8629[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8629[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8629[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8629[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8629[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51404_1_lut_4_lut (.I0(n14), .I1(n9), .I2(n70793), .I3(n70769), 
            .O(n67191));
    defparam i51404_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8629[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8629[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1031 (.I0(n14), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n69941));
    defparam i1_2_lut_3_lut_adj_1031.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8629[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8629[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8629[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8629[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8629[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8603[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8603[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8603[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8603[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8603[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8603[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8603[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8603[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51388_1_lut (.I0(n25968), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n67175));
    defparam i51388_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8603[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8603[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8603[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8603[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8603[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8603[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8603[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8577[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8577[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8577[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8577[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8577[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8577[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8577[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8577[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8577[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8577[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59804_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n75639));
    defparam i59804_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8577[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8577[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8577[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8577[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8551[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8551[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1032 (.I0(n77432), .I1(baudrate[18]), .I2(n2713), 
            .I3(n69405), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1032.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8551[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8551[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8551[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8551[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59808_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n75643));
    defparam i59808_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i62622_2_lut_4_lut (.I0(n77432), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25965), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i62622_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8551[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8551[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8551[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8551[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8551[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8551[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8551[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8551[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8525[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8525[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8525[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8525[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8525[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8525[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8525[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8525[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8525[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8525[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8525[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8525[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8525[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8525[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58870_4_lut (.I0(n25_adj_5283), .I1(n23_adj_5280), .I2(n21_adj_5279), 
            .I3(n19_adj_5285), .O(n74705));
    defparam i58870_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i58865_4_lut (.I0(n31_adj_5282), .I1(n29_adj_5281), .I2(n27_adj_5284), 
            .I3(n74705), .O(n74700));
    defparam i58865_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61033_4_lut (.I0(n37_adj_5278), .I1(n35_adj_5277), .I2(n33_adj_5276), 
            .I3(n74700), .O(n76868));
    defparam i61033_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2491), .I3(GND_net), .O(n18_adj_5286));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61207_3_lut (.I0(n18_adj_5286), .I1(baudrate[13]), .I2(n41_adj_5274), 
            .I3(GND_net), .O(n77042));   // verilog/uart_rx.v(119[33:55])
    defparam i61207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61208_3_lut (.I0(n77042), .I1(baudrate[14]), .I2(n43_adj_5275), 
            .I3(GND_net), .O(n77043));   // verilog/uart_rx.v(119[33:55])
    defparam i61208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59840_4_lut (.I0(n43_adj_5275), .I1(n41_adj_5274), .I2(n29_adj_5281), 
            .I3(n74703), .O(n75675));
    defparam i59840_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5177), .I1(baudrate[7]), 
            .I2(n29_adj_5281), .I3(GND_net), .O(n26_adj_5287));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61150_3_lut (.I0(n77043), .I1(baudrate[15]), .I2(n45_adj_5273), 
            .I3(GND_net), .O(n76985));   // verilog/uart_rx.v(119[33:55])
    defparam i61150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5176), .I1(baudrate[9]), 
            .I2(n33_adj_5276), .I3(GND_net), .O(n30_adj_5288));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61636_4_lut (.I0(n30_adj_5288), .I1(n20_adj_5175), .I2(n33_adj_5276), 
            .I3(n74698), .O(n77471));   // verilog/uart_rx.v(119[33:55])
    defparam i61636_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61637_3_lut (.I0(n77471), .I1(baudrate[10]), .I2(n35_adj_5277), 
            .I3(GND_net), .O(n77472));   // verilog/uart_rx.v(119[33:55])
    defparam i61637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61437_3_lut (.I0(n77472), .I1(baudrate[11]), .I2(n37_adj_5278), 
            .I3(GND_net), .O(n77272));   // verilog/uart_rx.v(119[33:55])
    defparam i61437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59844_4_lut (.I0(n43_adj_5275), .I1(n41_adj_5274), .I2(n39_adj_5272), 
            .I3(n76868), .O(n75679));
    defparam i59844_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61151_4_lut (.I0(n76985), .I1(n26_adj_5287), .I2(n45_adj_5273), 
            .I3(n75675), .O(n76986));   // verilog/uart_rx.v(119[33:55])
    defparam i61151_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61415_3_lut (.I0(n77272), .I1(baudrate[12]), .I2(n39_adj_5272), 
            .I3(GND_net), .O(n77250));   // verilog/uart_rx.v(119[33:55])
    defparam i61415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61593_4_lut (.I0(n77250), .I1(n76986), .I2(n45_adj_5273), 
            .I3(n75679), .O(n77428));   // verilog/uart_rx.v(119[33:55])
    defparam i61593_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8499[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8499[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8499[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8499[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8499[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8499[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8499[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8499[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8499[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8499[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8473[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8473[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58894_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n74729));
    defparam i58894_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8473[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8473[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1033 (.I0(n77544), .I1(baudrate[17]), .I2(n2596), 
            .I3(n69403), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1033.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8473[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8473[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1034 (.I0(n26008), .I1(n48_adj_5064), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1034.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8473[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8473[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8473[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1035 (.I0(n71544), .I1(n48_adj_5051), .I2(n8447[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_1035.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8473[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8447[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8447[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8447[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8447[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8447[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8447[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8447[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8447[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8447[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62619_2_lut_4_lut (.I0(n77544), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25935), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i62619_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8447[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n69945));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'h7bde;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8421[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5289));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8421[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8421[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(r_Clock_Count[3]), .I1(n3_adj_5289), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n69945), .O(n69949));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58898_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n74733));
    defparam i58898_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8421[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8421[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(n69395), .I1(n48_adj_5040), .I2(GND_net), 
            .I3(GND_net), .O(n1977));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8421[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n69949), .O(n69953));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hffde;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8421[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8421[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8395[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8395[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5290));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(r_Clock_Count[6]), .I1(n8_adj_5290), 
            .I2(n69953), .I3(\o_Rx_DV_N_3488[7] ), .O(n65798));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'hfdfe;
    SB_LUT4 i55637_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n65798), .I2(GND_net), 
            .I3(GND_net), .O(n71462));
    defparam i55637_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i55708_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n71462), .O(n71534));
    defparam i55708_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n69523), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i1_3_lut_4_lut_adj_1041 (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n69971), .I3(n71496), .O(n69923));
    defparam i1_3_lut_4_lut_adj_1041.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8395[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n71534), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11915));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11915), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8395[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8369[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5291));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8369[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1042 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[15]), .I3(baudrate[14]), .O(n70745));
    defparam i1_2_lut_3_lut_4_lut_adj_1042.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8369[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5292));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8369[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5293));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5294));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1043 (.I0(n77474), .I1(baudrate[15]), .I2(n2353), 
            .I3(n69399), .O(n2491));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1043.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8369[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62613_2_lut_4_lut (.I0(n77474), .I1(baudrate[15]), .I2(n2353), 
            .I3(n26014), .O(n294[8]));   // verilog/uart_rx.v(119[33:55])
    defparam i62613_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1044 (.I0(baudrate[18]), .I1(baudrate[19]), 
            .I2(baudrate[20]), .I3(baudrate[21]), .O(n70769));
    defparam i1_2_lut_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i30672_rep_5_2_lut (.I0(n8369[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n67207));   // verilog/uart_rx.v(119[33:55])
    defparam i30672_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n67207), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5295));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61237_3_lut (.I0(n32_adj_5295), .I1(baudrate[6]), .I2(n39_adj_5293), 
            .I3(GND_net), .O(n77072));   // verilog/uart_rx.v(119[33:55])
    defparam i61237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1045 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n70805), .I3(n70745), .O(n70749));
    defparam i1_3_lut_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 i61238_3_lut (.I0(n77072), .I1(baudrate[7]), .I2(n41_adj_5294), 
            .I3(GND_net), .O(n77073));   // verilog/uart_rx.v(119[33:55])
    defparam i61238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60049_4_lut (.I0(n41_adj_5294), .I1(n39_adj_5293), .I2(n37_adj_5292), 
            .I3(n74903), .O(n75884));
    defparam i60049_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60753_3_lut (.I0(n34_adj_5253), .I1(baudrate[5]), .I2(n37_adj_5292), 
            .I3(GND_net), .O(n76588));   // verilog/uart_rx.v(119[33:55])
    defparam i60753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61118_3_lut (.I0(n77073), .I1(baudrate[8]), .I2(n43_adj_5291), 
            .I3(GND_net), .O(n76953));   // verilog/uart_rx.v(119[33:55])
    defparam i61118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61235_4_lut (.I0(n76953), .I1(n76588), .I2(n43_adj_5291), 
            .I3(n75884), .O(n77070));   // verilog/uart_rx.v(119[33:55])
    defparam i61235_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61236_3_lut (.I0(n77070), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n77071));   // verilog/uart_rx.v(119[33:55])
    defparam i61236_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61120_3_lut (.I0(n77071), .I1(baudrate[10]), .I2(n1693), 
            .I3(GND_net), .O(n48_adj_5296));   // verilog/uart_rx.v(119[33:55])
    defparam i61120_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n70803), .I1(n70819), .I2(n70817), 
            .I3(baudrate[11]), .O(n70747));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1047 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n70767), .I3(GND_net), .O(n70793));
    defparam i1_2_lut_3_lut_adj_1047.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1048 (.I0(baudrate[14]), .I1(baudrate[15]), 
            .I2(baudrate[17]), .I3(baudrate[16]), .O(n70643));
    defparam i1_2_lut_3_lut_4_lut_adj_1048.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1049 (.I0(n77310), .I1(baudrate[14]), .I2(n2227), 
            .I3(n69397), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1049.LUT_INIT = 16'h7100;
    SB_LUT4 i1_3_lut_adj_1050 (.I0(n70749), .I1(n69941), .I2(n70747), 
            .I3(GND_net), .O(n26027));
    defparam i1_3_lut_adj_1050.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1051 (.I0(n26027), .I1(n48_adj_5296), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1051.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8369[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8395[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62610_2_lut_4_lut (.I0(n77310), .I1(baudrate[14]), .I2(n2227), 
            .I3(n71542), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i62610_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8369[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8395[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8369[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8369[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8395[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8395[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8343[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8343[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8343[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8343[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8343[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8343[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(n69393), .I1(n48_adj_5028), .I2(GND_net), 
            .I3(GND_net), .O(n1560));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8343[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8317[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8317[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8317[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8317[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8317[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8317[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8291[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5844_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n67643), .I3(n44_adj_5244), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i5844_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i742_4_lut (.I0(n66912), .I1(n294[18]), .I2(n46), .I3(baudrate[5]), 
            .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5297));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58917_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n74752));
    defparam i58917_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5298));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5252), .I1(baudrate[4]), 
            .I2(n43_adj_5297), .I3(GND_net), .O(n42_adj_5299));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61249_4_lut (.I0(n42_adj_5299), .I1(n38_adj_5298), .I2(n43_adj_5297), 
            .I3(n74978), .O(n77084));   // verilog/uart_rx.v(119[33:55])
    defparam i61249_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61250_3_lut (.I0(n77084), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n77085));   // verilog/uart_rx.v(119[33:55])
    defparam i61250_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58921_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n74756));
    defparam i58921_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7317_4_lut (.I0(n960), .I1(n11690), .I2(n21187), .I3(baudrate[3]), 
            .O(n21189));   // verilog/uart_rx.v(119[33:55])
    defparam i7317_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i55684_2_lut_4_lut (.I0(baudrate[20]), .I1(baudrate[21]), .I2(baudrate[30]), 
            .I3(baudrate[22]), .O(n71510));
    defparam i55684_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5244), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8291[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7316_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21187));   // verilog/uart_rx.v(119[33:55])
    defparam i7316_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i5830_2_lut (.I0(n21187), .I1(n11690), .I2(GND_net), .I3(GND_net), 
            .O(n42_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam i5830_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5251), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8291[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5822_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5300));   // verilog/uart_rx.v(119[33:55])
    defparam i5822_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5300), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8291[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1053 (.I0(n26033), .I1(n48), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1053.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8291[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i62194_2_lut_4_lut (.I0(n77602), .I1(baudrate[13]), .I2(n2098), 
            .I3(n26008), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i62194_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i5673_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n67659), .I3(n44_adj_5245), 
            .O(n46_adj_5301));   // verilog/uart_rx.v(119[33:55])
    defparam i5673_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i639_4_lut (.I0(n66910), .I1(n294[19]), .I2(n46_adj_5301), 
            .I3(baudrate[4]), .O(n66912));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5250), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i7310_4_lut (.I0(n804), .I1(n44716), .I2(n21177), .I3(baudrate[2]), 
            .O(n21179));   // verilog/uart_rx.v(119[33:55])
    defparam i7310_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i58955_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n74790));
    defparam i58955_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5245), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i1_4_lut_adj_1054 (.I0(n25989), .I1(n48_adj_5171), .I2(n44718), 
            .I3(baudrate[2]), .O(n67667));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'hefff;
    SB_LUT4 i5504_4_lut (.I0(n644), .I1(baudrate[2]), .I2(n67667), .I3(n44_adj_5172), 
            .O(n46_adj_5302));   // verilog/uart_rx.v(119[33:55])
    defparam i5504_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i534_4_lut (.I0(n66908), .I1(n294[20]), .I2(n46_adj_5302), 
            .I3(baudrate[3]), .O(n66910));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59727_4_lut (.I0(n25989), .I1(n74882), .I2(n48_adj_5171), 
            .I3(baudrate[0]), .O(n804));
    defparam i59727_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i55674_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), .I2(baudrate[12]), 
            .I3(baudrate[11]), .O(n71500));
    defparam i55674_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1055 (.I0(n26020), .I1(n48_adj_5173), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1055.LUT_INIT = 16'hefef;
    SB_LUT4 i62633_2_lut (.I0(n48_adj_5171), .I1(n25989), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i62633_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i55718_2_lut_3_lut (.I0(baudrate[13]), .I1(baudrate[14]), .I2(n71542), 
            .I3(GND_net), .O(n71544));
    defparam i55718_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i55690_4_lut (.I0(baudrate[1]), .I1(n71496), .I2(n69971), 
            .I3(baudrate[3]), .O(n71516));
    defparam i55690_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n71516), .I1(n71542), .I2(n71498), 
            .I3(n69833), .O(n48_adj_5303));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'h0100;
    SB_LUT4 i2314_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2314_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_2_lut_4_lut_adj_1057 (.I0(n70805), .I1(n70803), .I2(n70799), 
            .I3(n70801), .O(n70773));
    defparam i1_2_lut_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n69923), .I1(n25935), .I2(n71498), 
            .I3(n70643), .O(n25986));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 i62607_2_lut_4_lut (.I0(n77604), .I1(baudrate[12]), .I2(n1966), 
            .I3(n71544), .O(n294[11]));
    defparam i62607_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_adj_1059 (.I0(n25986), .I1(n48_adj_5303), .I2(n44718), 
            .I3(GND_net), .O(n67691));
    defparam i1_3_lut_adj_1059.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i427_4_lut (.I0(n5_adj_5304), .I1(n67691), .I2(n294[21]), 
            .I3(baudrate[2]), .O(n66908));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i62367_2_lut (.I0(baudrate[1]), .I1(n71574), .I2(GND_net), 
            .I3(GND_net), .O(n294[23]));
    defparam i62367_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n69395), .I3(n48_adj_5040), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(baudrate[23]), .I1(baudrate[1]), .I2(GND_net), 
            .I3(GND_net), .O(n69765));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h4444;
    SB_LUT4 i55694_4_lut (.I0(baudrate[19]), .I1(n69971), .I2(baudrate[3]), 
            .I3(baudrate[20]), .O(n71520));
    defparam i55694_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i55680_3_lut (.I0(baudrate[21]), .I1(baudrate[10]), .I2(baudrate[22]), 
            .I3(GND_net), .O(n71506));
    defparam i55680_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1061 (.I0(n71500), .I1(n71430), .I2(n70801), 
            .I3(n69765), .O(n69807));
    defparam i1_4_lut_adj_1061.LUT_INIT = 16'h0100;
    SB_LUT4 i55704_4_lut (.I0(n14), .I1(n71520), .I2(n71432), .I3(baudrate[2]), 
            .O(n71530));
    defparam i55704_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i55706_4_lut (.I0(n9), .I1(n23_adj_5180), .I2(n22_adj_5179), 
            .I3(n71506), .O(n71532));
    defparam i55706_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1062 (.I0(n45239), .I1(n71532), .I2(n71530), 
            .I3(n69807), .O(n5_adj_5304));   // verilog/uart_rx.v(119[33:55])
    defparam i1_4_lut_adj_1062.LUT_INIT = 16'habaa;
    SB_LUT4 div_37_LessThan_341_i48_4_lut (.I0(n71574), .I1(baudrate[2]), 
            .I2(n5_adj_5304), .I3(n44718), .O(n48_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_4_lut.LUT_INIT = 16'hd4c0;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58978_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n74813));
    defparam i58978_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i55721_1_lut_2_lut (.I0(baudrate[12]), .I1(n71544), .I2(GND_net), 
            .I3(GND_net), .O(n67204));
    defparam i55721_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5249));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i55607_2_lut (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n71432));
    defparam i55607_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i55605_2_lut (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n71430));
    defparam i55605_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30644_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n44718));
    defparam i30644_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1063 (.I0(baudrate[7]), .I1(baudrate[9]), .I2(baudrate[8]), 
            .I3(baudrate[10]), .O(n69873));
    defparam i1_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n69006));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_adj_1064 (.I0(n71500), .I1(n71430), .I2(n71432), 
            .I3(GND_net), .O(n69877));
    defparam i1_3_lut_adj_1064.LUT_INIT = 16'hfefe;
    SB_LUT4 i59137_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n74972));   // verilog/uart_rx.v(119[33:55])
    defparam i59137_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1065 (.I0(n69875), .I1(n25965), .I2(n69877), 
            .I3(n69873), .O(n25989));
    defparam i1_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 i2307_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2307_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i62604_2_lut_3_lut (.I0(baudrate[12]), .I1(n71544), .I2(n48_adj_5040), 
            .I3(GND_net), .O(n294[12]));
    defparam i62604_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_adj_1066 (.I0(n33), .I1(n25968), .I2(n70749), .I3(GND_net), 
            .O(n26020));
    defparam i1_3_lut_adj_1066.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n74573), .I1(baudrate[2]), 
            .I2(n644), .I3(n48_adj_5171), .O(n46_adj_5305));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5305), .I1(baudrate[3]), 
            .I2(n66908), .I3(GND_net), .O(n48_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i62096_2_lut (.I0(n48_adj_5173), .I1(n26020), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i62096_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i58999_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n74834));
    defparam i58999_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59730_4_lut (.I0(n25986), .I1(n74877), .I2(n48_adj_5303), 
            .I3(baudrate[0]), .O(n644));
    defparam i59730_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 div_37_i535_4_lut (.I0(n644), .I1(n44_adj_5172), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i62163_2_lut_4_lut (.I0(n77071), .I1(baudrate[10]), .I2(n1693), 
            .I3(n26027), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i62163_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n69393), .I3(n48_adj_5028), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5306));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60767_3_lut (.I0(n42_adj_5306), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n76602));   // verilog/uart_rx.v(119[33:55])
    defparam i60767_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60768_3_lut (.I0(n76602), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n76603));   // verilog/uart_rx.v(119[33:55])
    defparam i60768_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n76603), .I1(baudrate[4]), 
            .I2(n66910), .I3(GND_net), .O(n48_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_LessThan_965_i34_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n69391), .I3(n48_adj_5024), .O(n34_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(n70643), .I1(n70769), .I2(GND_net), 
            .I3(GND_net), .O(n70649));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(n71496), .I1(n25974), .I2(n70649), 
            .I3(n71498), .O(n26033));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'hfffe;
    SB_LUT4 i30649_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n67224));   // verilog/uart_rx.v(119[33:55])
    defparam i30649_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i62099_2_lut_4_lut (.I0(n77087), .I1(baudrate[5]), .I2(n66912), 
            .I3(n26033), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i62099_2_lut_4_lut.LUT_INIT = 16'h0017;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2872, pwm_out, clk32MHz, pwm_counter, GND_net, \pwm_counter[16] , 
            \pwm_counter[20] , \pwm_counter[19] , VCC_net, reset, \pwm_setpoint[2] , 
            \pwm_setpoint[3] , \pwm_setpoint[8] , \pwm_setpoint[4] , \pwm_setpoint[6] , 
            \pwm_setpoint[5] , \PWMLimit[6] , \data_in_frame[10][6] , 
            Kp_23__N_612, Kp_23__N_1748, n30764, \pwm_setpoint[22] , 
            \pwm_setpoint[21] , \pwm_setpoint[12] , \pwm_setpoint[10] , 
            \pwm_setpoint[11] , \pwm_setpoint[9] , \pwm_setpoint[7] , 
            n17, n13, \pwm_setpoint[1] , \pwm_setpoint[0] , \pwm_setpoint[13] , 
            \pwm_setpoint[14] , \pwm_setpoint[15] , n32, n34, \pwm_setpoint[20] , 
            n41, n39, \pwm_setpoint[19] , \pwm_setpoint[23] , \data_in_frame[12][7] , 
            \data_in_frame[12][0] , \data_in_frame[11][7] , n70983, \data_in_frame[10][5] , 
            n71189, \pwm_setpoint[18] , \pwm_setpoint[17] , n66769, 
            \data_in_frame[15][3] , n66751, n68353, n7, n69038, \data_in_frame[10][7] , 
            \data_in_frame[11][0] , n66791, n26329, n68099) /* synthesis syn_module_defined=1 */ ;
    input n2872;
    output pwm_out;
    input clk32MHz;
    output [23:0]pwm_counter;
    input GND_net;
    output \pwm_counter[16] ;
    output \pwm_counter[20] ;
    output \pwm_counter[19] ;
    input VCC_net;
    input reset;
    input \pwm_setpoint[2] ;
    input \pwm_setpoint[3] ;
    input \pwm_setpoint[8] ;
    input \pwm_setpoint[4] ;
    input \pwm_setpoint[6] ;
    input \pwm_setpoint[5] ;
    input \PWMLimit[6] ;
    input \data_in_frame[10][6] ;
    input Kp_23__N_612;
    input Kp_23__N_1748;
    output n30764;
    input \pwm_setpoint[22] ;
    input \pwm_setpoint[21] ;
    input \pwm_setpoint[12] ;
    input \pwm_setpoint[10] ;
    input \pwm_setpoint[11] ;
    input \pwm_setpoint[9] ;
    input \pwm_setpoint[7] ;
    input n17;
    input n13;
    input \pwm_setpoint[1] ;
    input \pwm_setpoint[0] ;
    input \pwm_setpoint[13] ;
    input \pwm_setpoint[14] ;
    input \pwm_setpoint[15] ;
    output n32;
    input n34;
    input \pwm_setpoint[20] ;
    input n41;
    input n39;
    input \pwm_setpoint[19] ;
    input \pwm_setpoint[23] ;
    input \data_in_frame[12][7] ;
    input \data_in_frame[12][0] ;
    input \data_in_frame[11][7] ;
    output n70983;
    input \data_in_frame[10][5] ;
    output n71189;
    input \pwm_setpoint[18] ;
    input \pwm_setpoint[17] ;
    input n66769;
    input \data_in_frame[15][3] ;
    input n66751;
    output n68353;
    input n7;
    input n69038;
    input \data_in_frame[10][7] ;
    input \data_in_frame[11][0] ;
    output n66791;
    input n26329;
    output n68099;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577;
    wire [23:0]pwm_counter_c;   // verilog/pwm.v(11[19:30])
    
    wire n69121, n22, n15, n20, n24, n19, n45, n64468, n59447, 
        n64508, n59446, n64540, n59445, n64580, n59444, n64620, 
        n59443, n64660, n59442, n64698, n59441, n64736, n59440, 
        n64766, n59439, n64806, n59438, n64838, n59437, n64876, 
        n59436, n64910, n59435, n64942, n59434, n64982, n59433, 
        n65032, n59432, n65076, n59431, n65136, n59430, n65258, 
        n59429, n65426, n59428, n65556, n59427, n65558, n59426, 
        n65560, n59425, n65550, n6, n75666, n8, n74692, n10, 
        n45_adj_5019, n43, n25, n21, n23, n19_adj_5020, n15_adj_5021, 
        n7_c, n9, n11, n5, n74716, n74679, n4, n12, n16, n77439, 
        n77440, n77328, n76864, n77441, n75791, n77528, n77529, 
        n77486, n77115, n77116, n75615, n76471, n36, n38, n75799, 
        n76896;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2872), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter_c[7]), 
            .I3(GND_net), .O(n69121));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter_c[11]), .I1(pwm_counter_c[18]), .I2(pwm_counter_c[15]), 
            .I3(pwm_counter_c[13]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n69121), .I1(\pwm_counter[16] ), .I2(pwm_counter_c[10]), 
            .I3(pwm_counter_c[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(\pwm_counter[20] ), .I1(pwm_counter_c[22]), .I2(pwm_counter_c[14]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(\pwm_counter[19] ), .I3(pwm_counter_c[12]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter_c[17]), .I1(pwm_counter_c[21]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter_c[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(n45));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_counter_2040_add_4_25_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[23]), 
            .I3(n59447), .O(n64468)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2040_add_4_24_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[22]), 
            .I3(n59446), .O(n64508)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_24 (.CI(n59446), .I0(GND_net), .I1(pwm_counter_c[22]), 
            .CO(n59447));
    SB_LUT4 pwm_counter_2040_add_4_23_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[21]), 
            .I3(n59445), .O(n64540)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_23 (.CI(n59445), .I0(GND_net), .I1(pwm_counter_c[21]), 
            .CO(n59446));
    SB_LUT4 pwm_counter_2040_add_4_22_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[20] ), 
            .I3(n59444), .O(n64580)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_22 (.CI(n59444), .I0(GND_net), .I1(\pwm_counter[20] ), 
            .CO(n59445));
    SB_LUT4 pwm_counter_2040_add_4_21_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n59443), .O(n64620)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_21 (.CI(n59443), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n59444));
    SB_LUT4 pwm_counter_2040_add_4_20_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[18]), 
            .I3(n59442), .O(n64660)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_20 (.CI(n59442), .I0(GND_net), .I1(pwm_counter_c[18]), 
            .CO(n59443));
    SB_LUT4 pwm_counter_2040_add_4_19_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[17]), 
            .I3(n59441), .O(n64698)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_19 (.CI(n59441), .I0(GND_net), .I1(pwm_counter_c[17]), 
            .CO(n59442));
    SB_LUT4 pwm_counter_2040_add_4_18_lut (.I0(n45), .I1(GND_net), .I2(\pwm_counter[16] ), 
            .I3(n59440), .O(n64736)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_18 (.CI(n59440), .I0(GND_net), .I1(\pwm_counter[16] ), 
            .CO(n59441));
    SB_LUT4 pwm_counter_2040_add_4_17_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[15]), 
            .I3(n59439), .O(n64766)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_17 (.CI(n59439), .I0(GND_net), .I1(pwm_counter_c[15]), 
            .CO(n59440));
    SB_LUT4 pwm_counter_2040_add_4_16_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[14]), 
            .I3(n59438), .O(n64806)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_16 (.CI(n59438), .I0(GND_net), .I1(pwm_counter_c[14]), 
            .CO(n59439));
    SB_LUT4 pwm_counter_2040_add_4_15_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[13]), 
            .I3(n59437), .O(n64838)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_15 (.CI(n59437), .I0(GND_net), .I1(pwm_counter_c[13]), 
            .CO(n59438));
    SB_LUT4 pwm_counter_2040_add_4_14_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[12]), 
            .I3(n59436), .O(n64876)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_14 (.CI(n59436), .I0(GND_net), .I1(pwm_counter_c[12]), 
            .CO(n59437));
    SB_LUT4 pwm_counter_2040_add_4_13_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[11]), 
            .I3(n59435), .O(n64910)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_13 (.CI(n59435), .I0(GND_net), .I1(pwm_counter_c[11]), 
            .CO(n59436));
    SB_LUT4 pwm_counter_2040_add_4_12_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[10]), 
            .I3(n59434), .O(n64942)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_12 (.CI(n59434), .I0(GND_net), .I1(pwm_counter_c[10]), 
            .CO(n59435));
    SB_LUT4 pwm_counter_2040_add_4_11_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[9]), 
            .I3(n59433), .O(n64982)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_11 (.CI(n59433), .I0(GND_net), .I1(pwm_counter_c[9]), 
            .CO(n59434));
    SB_LUT4 pwm_counter_2040_add_4_10_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n59432), .O(n65032)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_10 (.CI(n59432), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n59433));
    SB_LUT4 pwm_counter_2040_add_4_9_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[7]), 
            .I3(n59431), .O(n65076)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_9 (.CI(n59431), .I0(GND_net), .I1(pwm_counter_c[7]), 
            .CO(n59432));
    SB_LUT4 pwm_counter_2040_add_4_8_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n59430), .O(n65136)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_8 (.CI(n59430), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n59431));
    SB_LUT4 pwm_counter_2040_add_4_7_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[5]), 
            .I3(n59429), .O(n65258)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_7 (.CI(n59429), .I0(GND_net), .I1(pwm_counter_c[5]), 
            .CO(n59430));
    SB_LUT4 pwm_counter_2040_add_4_6_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[4]), 
            .I3(n59428), .O(n65426)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_6 (.CI(n59428), .I0(GND_net), .I1(pwm_counter_c[4]), 
            .CO(n59429));
    SB_LUT4 pwm_counter_2040_add_4_5_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[3]), 
            .I3(n59427), .O(n65556)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_5 (.CI(n59427), .I0(GND_net), .I1(pwm_counter_c[3]), 
            .CO(n59428));
    SB_LUT4 pwm_counter_2040_add_4_4_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[2]), 
            .I3(n59426), .O(n65558)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_4 (.CI(n59426), .I0(GND_net), .I1(pwm_counter_c[2]), 
            .CO(n59427));
    SB_LUT4 pwm_counter_2040_add_4_3_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[1]), 
            .I3(n59425), .O(n65560)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_3 (.CI(n59425), .I0(GND_net), .I1(pwm_counter_c[1]), 
            .CO(n59426));
    SB_LUT4 pwm_counter_2040_add_4_2_lut (.I0(n45), .I1(GND_net), .I2(pwm_counter_c[0]), 
            .I3(VCC_net), .O(n65550)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter_c[0]), 
            .CO(n59425));
    SB_DFFR pwm_counter_2040__i0 (.Q(pwm_counter_c[0]), .C(clk32MHz), .D(n65550), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i23 (.Q(pwm_counter_c[23]), .C(clk32MHz), 
            .D(n64468), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i22 (.Q(pwm_counter_c[22]), .C(clk32MHz), 
            .D(n64508), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i21 (.Q(pwm_counter_c[21]), .C(clk32MHz), 
            .D(n64540), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i20 (.Q(\pwm_counter[20] ), .C(clk32MHz), 
            .D(n64580), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n64620), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i18 (.Q(pwm_counter_c[18]), .C(clk32MHz), 
            .D(n64660), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i17 (.Q(pwm_counter_c[17]), .C(clk32MHz), 
            .D(n64698), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i16 (.Q(\pwm_counter[16] ), .C(clk32MHz), 
            .D(n64736), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i15 (.Q(pwm_counter_c[15]), .C(clk32MHz), 
            .D(n64766), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i14 (.Q(pwm_counter_c[14]), .C(clk32MHz), 
            .D(n64806), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i13 (.Q(pwm_counter_c[13]), .C(clk32MHz), 
            .D(n64838), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i12 (.Q(pwm_counter_c[12]), .C(clk32MHz), 
            .D(n64876), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i11 (.Q(pwm_counter_c[11]), .C(clk32MHz), 
            .D(n64910), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i10 (.Q(pwm_counter_c[10]), .C(clk32MHz), 
            .D(n64942), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i9 (.Q(pwm_counter_c[9]), .C(clk32MHz), .D(n64982), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n65032), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i7 (.Q(pwm_counter_c[7]), .C(clk32MHz), .D(n65076), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n65136), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i5 (.Q(pwm_counter_c[5]), .C(clk32MHz), .D(n65258), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i4 (.Q(pwm_counter_c[4]), .C(clk32MHz), .D(n65426), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i3 (.Q(pwm_counter_c[3]), .C(clk32MHz), .D(n65556), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i2 (.Q(pwm_counter_c[2]), .C(clk32MHz), .D(n65558), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i1 (.Q(pwm_counter_c[1]), .C(clk32MHz), .D(n65560), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(\pwm_setpoint[2] ), .I1(\pwm_setpoint[3] ), 
            .I2(pwm_counter_c[3]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59831_2_lut_4_lut (.I0(\pwm_setpoint[8] ), .I1(pwm_counter[8]), 
            .I2(pwm_counter_c[4]), .I3(\pwm_setpoint[4] ), .O(n75666));
    defparam i59831_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(\pwm_setpoint[4] ), .I1(\pwm_setpoint[8] ), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i58857_2_lut_4_lut (.I0(\pwm_setpoint[6] ), .I1(pwm_counter[6]), 
            .I2(pwm_counter_c[5]), .I3(\pwm_setpoint[5] ), .O(n74692));
    defparam i58857_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(\pwm_setpoint[5] ), .I1(\pwm_setpoint[6] ), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i23332_3_lut_4_lut (.I0(\PWMLimit[6] ), .I1(\data_in_frame[10][6] ), 
            .I2(Kp_23__N_612), .I3(Kp_23__N_1748), .O(n30764));
    defparam i23332_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter_c[22]), .I1(\pwm_setpoint[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5019));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter_c[21]), .I1(\pwm_setpoint[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter_c[12]), .I1(\pwm_setpoint[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter_c[10]), .I1(\pwm_setpoint[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter_c[11]), .I1(\pwm_setpoint[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter_c[9]), .I1(\pwm_setpoint[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5020));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter_c[7]), .I1(\pwm_setpoint[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5021));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i7_2_lut (.I0(pwm_counter_c[3]), .I1(\pwm_setpoint[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n7_c));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter_c[4]), .I1(\pwm_setpoint[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter_c[5]), .I1(\pwm_setpoint[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i5_2_lut (.I0(pwm_counter_c[2]), .I1(\pwm_setpoint[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i58881_4_lut (.I0(n11), .I1(n9), .I2(n7_c), .I3(n5), .O(n74716));
    defparam i58881_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i58844_4_lut (.I0(n17), .I1(n15_adj_5021), .I2(n13), .I3(n74716), 
            .O(n74679));
    defparam i58844_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter_c[0]), .I1(\pwm_setpoint[1] ), 
            .I2(pwm_counter_c[1]), .I3(\pwm_setpoint[0] ), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(n10), .I1(\pwm_setpoint[7] ), .I2(n15_adj_5021), 
            .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(n8), .I1(\pwm_setpoint[9] ), .I2(n19_adj_5020), 
            .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61604_4_lut (.I0(n16), .I1(n6), .I2(n19_adj_5020), .I3(n75666), 
            .O(n77439));   // verilog/pwm.v(21[8:24])
    defparam i61604_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61605_3_lut (.I0(n77439), .I1(\pwm_setpoint[10] ), .I2(n21), 
            .I3(GND_net), .O(n77440));   // verilog/pwm.v(21[8:24])
    defparam i61605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61493_3_lut (.I0(n77440), .I1(\pwm_setpoint[11] ), .I2(n23), 
            .I3(GND_net), .O(n77328));   // verilog/pwm.v(21[8:24])
    defparam i61493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61029_4_lut (.I0(n23), .I1(n21), .I2(n19_adj_5020), .I3(n74679), 
            .O(n76864));
    defparam i61029_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61606_4_lut (.I0(n12), .I1(n4), .I2(n15_adj_5021), .I3(n74692), 
            .O(n77441));   // verilog/pwm.v(21[8:24])
    defparam i61606_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59956_3_lut (.I0(n77328), .I1(\pwm_setpoint[12] ), .I2(n25), 
            .I3(GND_net), .O(n75791));   // verilog/pwm.v(21[8:24])
    defparam i59956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61693_4_lut (.I0(n75791), .I1(n77441), .I2(n25), .I3(n76864), 
            .O(n77528));   // verilog/pwm.v(21[8:24])
    defparam i61693_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61694_3_lut (.I0(n77528), .I1(\pwm_setpoint[13] ), .I2(pwm_counter_c[13]), 
            .I3(GND_net), .O(n77529));   // verilog/pwm.v(21[8:24])
    defparam i61694_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61651_3_lut (.I0(n77529), .I1(\pwm_setpoint[14] ), .I2(pwm_counter_c[14]), 
            .I3(GND_net), .O(n77486));   // verilog/pwm.v(21[8:24])
    defparam i61651_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59962_3_lut (.I0(n77486), .I1(\pwm_setpoint[15] ), .I2(pwm_counter_c[15]), 
            .I3(GND_net), .O(n32));   // verilog/pwm.v(21[8:24])
    defparam i59962_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61280_3_lut (.I0(n34), .I1(\pwm_setpoint[20] ), .I2(n41), 
            .I3(GND_net), .O(n77115));   // verilog/pwm.v(21[8:24])
    defparam i61280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61281_3_lut (.I0(n77115), .I1(\pwm_setpoint[21] ), .I2(n43), 
            .I3(GND_net), .O(n77116));   // verilog/pwm.v(21[8:24])
    defparam i61281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60636_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n75615), 
            .O(n76471));
    defparam i60636_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 duty_23__I_0_i38_3_lut (.I0(n36), .I1(\pwm_setpoint[19] ), .I2(n39), 
            .I3(GND_net), .O(n38));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59964_3_lut (.I0(n77116), .I1(\pwm_setpoint[22] ), .I2(n45_adj_5019), 
            .I3(GND_net), .O(n75799));   // verilog/pwm.v(21[8:24])
    defparam i59964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61061_4_lut (.I0(n75799), .I1(n38), .I2(n45_adj_5019), .I3(n76471), 
            .O(n76896));   // verilog/pwm.v(21[8:24])
    defparam i61061_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61062_3_lut (.I0(n76896), .I1(pwm_counter_c[23]), .I2(\pwm_setpoint[23] ), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i61062_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[10][6] ), .I1(\data_in_frame[12][7] ), 
            .I2(\data_in_frame[12][0] ), .I3(\data_in_frame[11][7] ), .O(n70983));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[10][6] ), .I1(\data_in_frame[12][7] ), 
            .I2(\data_in_frame[10][5] ), .I3(GND_net), .O(n71189));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 duty_23__I_0_i36_3_lut_3_lut (.I0(pwm_counter_c[18]), .I1(\pwm_setpoint[18] ), 
            .I2(\pwm_setpoint[17] ), .I3(GND_net), .O(n36));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59780_3_lut_4_lut (.I0(pwm_counter_c[18]), .I1(\pwm_setpoint[18] ), 
            .I2(\pwm_setpoint[17] ), .I3(pwm_counter_c[17]), .O(n75615));   // verilog/pwm.v(21[8:24])
    defparam i59780_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i2_3_lut_adj_987 (.I0(n66769), .I1(\data_in_frame[15][3] ), 
            .I2(n66751), .I3(GND_net), .O(n68353));
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_988 (.I0(n7), .I1(n69038), .I2(\data_in_frame[10][7] ), 
            .I3(\data_in_frame[11][0] ), .O(n66791));
    defparam i1_4_lut_adj_988.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut (.I0(n26329), .I1(n66791), .I2(\data_in_frame[10][6] ), 
            .I3(GND_net), .O(n68099));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (enable_slow_N_4213, clk16MHz, GND_net, data, baudrate, 
            n28271, data_ready, n29943, ID, \state_7__N_3918[0] , 
            n30719, n30718, n30717, n30716, n30715, n30714, n30713, 
            n30704, n30703, n30702, n30701, n30700, n30699, n30698, 
            n30696, n68385, \state_7__N_4110[0] , \state[0] , scl_enable, 
            scl, sda_enable, sda_out, n11, n29968, n29967, n29965, 
            n29964, n29963, n29959, n29958, n6705, n30749, n8, 
            VCC_net, n44499, \state_7__N_4126[3] , n10, n4, n4_adj_6, 
            n25888, n25930, n44644) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output enable_slow_N_4213;
    input clk16MHz;
    input GND_net;
    output [7:0]data;
    output [31:0]baudrate;
    output n28271;
    output data_ready;
    input n29943;
    output [7:0]ID;
    input \state_7__N_3918[0] ;
    input n30719;
    input n30718;
    input n30717;
    input n30716;
    input n30715;
    input n30714;
    input n30713;
    input n30704;
    input n30703;
    input n30702;
    input n30701;
    input n30700;
    input n30699;
    input n30698;
    input n30696;
    output n68385;
    output \state_7__N_4110[0] ;
    output \state[0] ;
    output scl_enable;
    output scl;
    output sda_enable;
    output sda_out;
    output n11;
    input n29968;
    input n29967;
    input n29965;
    input n29964;
    input n29963;
    input n29959;
    input n29958;
    output n6705;
    input n30749;
    input n8;
    input VCC_net;
    output n44499;
    input \state_7__N_4126[3] ;
    output n10;
    output n4;
    output n4_adj_6;
    output n25888;
    output n25930;
    output n44644;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire ready_prev;
    wire [0:0]n5925;
    
    wire enable;
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire n38052, n44510, n30104, n120, n129, n52816, n30680, n52805, 
        n30681, n25750;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n28, n52852, n135;
    wire [2:0]n1;
    wire [15:0]delay_counter_15__N_3956;
    
    wire n28089;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n52782, n65212, rw, n29944, n28161, n29430, n60798, n4_c, 
        n47, n4_adj_5008, n28756, n74636, n10_c, n8_c, n65062, 
        n30712, n30711, n30710, n30709, n30708, n30707, n30706, 
        n30705, n30695, n30694, n30693, n30692, n30691, n30690, 
        n30689, n30688, n30687, n30686, n30685, n30684, n30683, 
        n30682;
    wire [7:0]state_7__N_3885;
    
    wire n68601;
    wire [15:0]n5391;
    
    wire n58410, n58409, n58408;
    wire [7:0]state_adj_5018;   // verilog/i2c_controller.v(33[12:17])
    
    wire n74670, n58407, n58406, n6936, n58405, n52770, n6935, 
        n58404, n6934, n58403, n6933, n58402, n6932, n58401, n58400, 
        n6930, n58399, n58398, n58397, n58396, n15, n45126, n53, 
        n60213, n10_adj_5011;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n65606, n71484, n17, n7, n28_adj_5013, n26, n27, n25;
    
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5925[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38052));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30436_2_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n44510));
    defparam i30436_2_lut.LUT_INIT = 16'hdddd;
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n30104));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i38758_4_lut (.I0(n120), .I1(n129), .I2(data[7]), .I3(baudrate[31]), 
            .O(n52816));   // verilog/eeprom.v(23[12:16])
    defparam i38758_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i38759_3_lut (.I0(n52816), .I1(baudrate[31]), .I2(state[2]), 
            .I3(GND_net), .O(n30680));   // verilog/eeprom.v(27[11:16])
    defparam i38759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38747_4_lut (.I0(n120), .I1(n129), .I2(data[6]), .I3(baudrate[30]), 
            .O(n52805));   // verilog/eeprom.v(23[12:16])
    defparam i38747_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i38748_3_lut (.I0(n52805), .I1(baudrate[30]), .I2(state[2]), 
            .I3(GND_net), .O(n30681));   // verilog/eeprom.v(27[11:16])
    defparam i38748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1515_Mux_0_i3_3_lut_4_lut (.I0(state[0]), .I1(enable_slow_N_4213), 
            .I2(n25750), .I3(state[1]), .O(n5925[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1515_Mux_0_i3_3_lut_4_lut.LUT_INIT = 16'h04aa;
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(byte_counter[1]), .I2(n28), 
            .I3(GND_net), .O(n52852));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_3_lut_adj_973 (.I0(state[2]), .I1(byte_counter[0]), .I2(n52852), 
            .I3(GND_net), .O(n28271));
    defparam i2_3_lut_adj_973.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(n44510), .O(n30104));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'ha8e8;
    SB_LUT4 i1_2_lut_adj_974 (.I0(byte_counter[0]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n135));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h2222;
    SB_LUT4 i43965_2_lut_3_lut_4_lut (.I0(enable_slow_N_4213), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n1[1]));   // verilog/eeprom.v(68[25:39])
    defparam i43965_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n28089), .D(delay_counter_15__N_3956[13]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n65212));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n29944));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29943));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n28161), .D(n1[1]), .R(n29430));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n28161), .D(n1[2]), .R(n29430));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n28161), .D(n60798), .R(n29430));   // verilog/eeprom.v(68[25:39])
    SB_LUT4 i1_2_lut_adj_975 (.I0(\state_7__N_3918[0] ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'heeee;
    SB_LUT4 i61823_3_lut (.I0(n47), .I1(n44510), .I2(state[0]), .I3(GND_net), 
            .O(n4_adj_5008));
    defparam i61823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(state[1]), .I1(state[2]), .I2(n4_adj_5008), 
            .I3(n4_c), .O(n28756));
    defparam i2_4_lut.LUT_INIT = 16'hecfd;
    SB_LUT4 i59109_3_lut (.I0(n28756), .I1(state[2]), .I2(\state_7__N_3918[0] ), 
            .I3(GND_net), .O(n74636));   // verilog/eeprom.v(27[11:16])
    defparam i59109_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i28_4_lut (.I0(n74636), .I1(n47), .I2(state[1]), .I3(n28756), 
            .O(n10_c));   // verilog/eeprom.v(27[11:16])
    defparam i28_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i27_4_lut (.I0(n10_c), .I1(n8_c), .I2(state[0]), .I3(state[2]), 
            .O(n65062));   // verilog/eeprom.v(27[11:16])
    defparam i27_4_lut.LUT_INIT = 16'hfaca;
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n65062));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30719));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30718));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30717));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30716));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30715));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30714));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30713));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30712));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30711));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30710));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30709));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30708));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30707));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30706));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30705));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30704));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30703));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30702));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30701));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n30700));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n30699));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n30698));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n30696));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30695));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30694));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30693));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30692));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30691));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30690));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30689));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30688));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30687));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30686));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30685));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30684));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30683));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30682));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30681));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30680));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n68601), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1198_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5391[9]), 
            .I3(n58410), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1198_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5391[9]), 
            .I3(n58409), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_16 (.CI(n58409), .I0(delay_counter[14]), .I1(n5391[9]), 
            .CO(n58410));
    SB_LUT4 add_1198_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5391[9]), 
            .I3(n58408), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_15 (.CI(n58408), .I0(delay_counter[13]), .I1(n5391[9]), 
            .CO(n58409));
    SB_LUT4 i58958_2_lut_3_lut (.I0(state_adj_5018[1]), .I1(state_adj_5018[2]), 
            .I2(state[1]), .I3(GND_net), .O(n74670));
    defparam i58958_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 add_1198_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5391[9]), 
            .I3(n58407), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_14 (.CI(n58407), .I0(delay_counter[12]), .I1(n5391[9]), 
            .CO(n58408));
    SB_LUT4 add_1198_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5391[9]), 
            .I3(n58406), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_13 (.CI(n58406), .I0(delay_counter[11]), .I1(n5391[9]), 
            .CO(n58407));
    SB_LUT4 add_1198_12_lut (.I0(n52770), .I1(delay_counter[10]), .I2(n5391[9]), 
            .I3(n58405), .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_12 (.CI(n58405), .I0(delay_counter[10]), .I1(n5391[9]), 
            .CO(n58406));
    SB_LUT4 add_1198_11_lut (.I0(n52770), .I1(delay_counter[9]), .I2(n5391[9]), 
            .I3(n58404), .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_11 (.CI(n58404), .I0(delay_counter[9]), .I1(n5391[9]), 
            .CO(n58405));
    SB_LUT4 add_1198_10_lut (.I0(n52770), .I1(delay_counter[8]), .I2(n5391[9]), 
            .I3(n58403), .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_10 (.CI(n58403), .I0(delay_counter[8]), .I1(n5391[9]), 
            .CO(n58404));
    SB_LUT4 add_1198_9_lut (.I0(n52770), .I1(delay_counter[7]), .I2(n5391[9]), 
            .I3(n58402), .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_9 (.CI(n58402), .I0(delay_counter[7]), .I1(n5391[9]), 
            .CO(n58403));
    SB_LUT4 add_1198_8_lut (.I0(n52770), .I1(delay_counter[6]), .I2(n5391[9]), 
            .I3(n58401), .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_8 (.CI(n58401), .I0(delay_counter[6]), .I1(n5391[9]), 
            .CO(n58402));
    SB_LUT4 add_1198_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5391[9]), 
            .I3(n58400), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_7 (.CI(n58400), .I0(delay_counter[5]), .I1(n5391[9]), 
            .CO(n58401));
    SB_LUT4 add_1198_6_lut (.I0(n52770), .I1(delay_counter[4]), .I2(n5391[9]), 
            .I3(n58399), .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_6 (.CI(n58399), .I0(delay_counter[4]), .I1(n5391[9]), 
            .CO(n58400));
    SB_LUT4 add_1198_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5391[9]), 
            .I3(n58398), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_5 (.CI(n58398), .I0(delay_counter[3]), .I1(n5391[9]), 
            .CO(n58399));
    SB_LUT4 add_1198_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5391[9]), 
            .I3(n58397), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_4 (.CI(n58397), .I0(delay_counter[2]), .I1(n5391[9]), 
            .CO(n58398));
    SB_LUT4 add_1198_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5391[9]), 
            .I3(n58396), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_3 (.CI(n58396), .I0(delay_counter[1]), .I1(n5391[9]), 
            .CO(n58397));
    SB_LUT4 add_1198_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5391[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5391[9]), 
            .CO(n58396));
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n28089), .D(delay_counter_15__N_3956[15]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n28089), .D(delay_counter_15__N_3956[14]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n28089), .D(delay_counter_15__N_3956[12]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n28089), .D(delay_counter_15__N_3956[11]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n28089), .D(n6936), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n28089), 
            .D(n6935), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n28089), 
            .D(n6934), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n28089), 
            .D(n6933), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n28089), 
            .D(n6932), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n28089), 
            .D(delay_counter_15__N_3956[5]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n28089), 
            .D(n6930), .S(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n28089), 
            .D(delay_counter_15__N_3956[3]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n28089), 
            .D(delay_counter_15__N_3956[2]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n28089), 
            .D(delay_counter_15__N_3956[1]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n28089), 
            .D(delay_counter_15__N_3956[0]), .R(n52782));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i12_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(n38052), .I3(data_ready), 
            .O(n29944));   // verilog/eeprom.v(27[11:16])
    defparam i12_4_lut_4_lut.LUT_INIT = 16'hfa08;
    SB_LUT4 i2_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(state[2]), 
            .I3(\state_7__N_3918[0] ), .O(n28161));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0908;
    SB_LUT4 i3_4_lut (.I0(ready_prev), .I1(n45126), .I2(state[0]), .I3(state[1]), 
            .O(n28));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i15218_3_lut_4_lut (.I0(n28161), .I1(state[2]), .I2(state[0]), 
            .I3(state[1]), .O(n29430));   // verilog/eeprom.v(68[25:39])
    defparam i15218_3_lut_4_lut.LUT_INIT = 16'h8aaa;
    SB_LUT4 i2_3_lut_adj_976 (.I0(state[2]), .I1(byte_counter[0]), .I2(n53), 
            .I3(GND_net), .O(n68385));
    defparam i2_3_lut_adj_976.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(rw), .I2(n60213), .I3(state[2]), 
            .O(n10_adj_5011));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut.LUT_INIT = 16'h888a;
    SB_LUT4 i1_4_lut_adj_977 (.I0(n10_adj_5011), .I1(rw), .I2(state[0]), 
            .I3(state[2]), .O(n65212));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut_adj_977.LUT_INIT = 16'heeae;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4213), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n60798));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i1_4_lut_adj_978 (.I0(n45126), .I1(saved_addr[0]), .I2(rw), 
            .I3(\state_7__N_4110[0] ), .O(n65606));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_978.LUT_INIT = 16'hd8cc;
    SB_LUT4 i1_2_lut_3_lut_adj_979 (.I0(state[1]), .I1(enable_slow_N_4213), 
            .I2(ready_prev), .I3(GND_net), .O(n8_c));   // verilog/eeprom.v(27[11:16])
    defparam i1_2_lut_3_lut_adj_979.LUT_INIT = 16'ha2a2;
    SB_LUT4 i18_2_lut (.I0(state[2]), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n52770));
    defparam i18_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i61940_2_lut (.I0(n25750), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5391[9]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i61940_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i55658_3_lut (.I0(\state[0] ), .I1(n25750), .I2(state_adj_5018[3]), 
            .I3(GND_net), .O(n71484));
    defparam i55658_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n74670), .I1(n8_c), .I2(state[0]), .I3(n71484), 
            .O(n17));
    defparam i24_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i2_4_lut_adj_980 (.I0(n17), .I1(state[2]), .I2(\state_7__N_3918[0] ), 
            .I3(state[1]), .O(n68601));
    defparam i2_4_lut_adj_980.LUT_INIT = 16'heefe;
    SB_LUT4 i38764_4_lut (.I0(state[1]), .I1(n15), .I2(state[2]), .I3(state[0]), 
            .O(state_7__N_3885[1]));   // verilog/eeprom.v(27[11:16])
    defparam i38764_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 i2_3_lut_4_lut (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(n28), .I3(byte_counter[2]), .O(n120));   // verilog/eeprom.v(30[11:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_981 (.I0(byte_counter[0]), .I1(byte_counter[1]), 
            .I2(byte_counter[2]), .I3(GND_net), .O(n15));   // verilog/eeprom.v(30[11:23])
    defparam i1_2_lut_3_lut_adj_981.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(\state[0] ), .I1(state_adj_5018[3]), 
            .I2(n7), .I3(n25750), .O(n47));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_983 (.I0(\state[0] ), .I1(state_adj_5018[3]), 
            .I2(state_adj_5018[2]), .I3(state_adj_5018[1]), .O(n45126));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(state[0]), 
            .I3(state[1]), .O(n52782));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h0052;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(state[2]), .I1(n15), .I2(state[0]), 
            .I3(state[1]), .O(n28089));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0552;
    SB_LUT4 i2_3_lut_4_lut_adj_984 (.I0(byte_counter[1]), .I1(n28), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n129));
    defparam i2_3_lut_4_lut_adj_984.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_985 (.I0(byte_counter[1]), .I1(n28), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n53));
    defparam i1_2_lut_3_lut_adj_985.LUT_INIT = 16'hfbfb;
    SB_LUT4 i43972_3_lut_4_lut (.I0(n44510), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n1[2]));   // verilog/eeprom.v(68[25:39])
    defparam i43972_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i2_2_lut (.I0(state_adj_5018[1]), .I1(state_adj_5018[2]), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(55[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(delay_counter[10]), .I1(delay_counter[15]), .I2(delay_counter[8]), 
            .I3(delay_counter[14]), .O(n28_adj_5013));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[3]), .I2(delay_counter[7]), 
            .I3(delay_counter[1]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[2]), .I1(delay_counter[12]), .I2(delay_counter[6]), 
            .I3(delay_counter[5]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28_adj_5013), 
            .O(n25750));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_986 (.I0(state[0]), .I1(enable_slow_N_4213), .I2(n25750), 
            .I3(GND_net), .O(n60213));
    defparam i2_3_lut_adj_986.LUT_INIT = 16'hfbfb;
    SB_LUT4 i16500_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[0]), .I3(baudrate[0]), 
            .O(n30712));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16500_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16493_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[7]), .I3(baudrate[7]), 
            .O(n30705));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16493_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16494_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[6]), .I3(baudrate[6]), 
            .O(n30706));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16494_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16495_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[5]), .I3(baudrate[5]), 
            .O(n30707));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16495_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16496_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[4]), .I3(baudrate[4]), 
            .O(n30708));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16496_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16497_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[3]), .I3(baudrate[3]), 
            .O(n30709));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16497_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16498_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[2]), .I3(baudrate[2]), 
            .O(n30710));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16498_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16499_3_lut_4_lut (.I0(n53), .I1(n135), .I2(data[1]), .I3(baudrate[1]), 
            .O(n30711));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16499_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16483_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30695));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16483_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16476_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30688));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16476_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16477_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30689));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16477_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16478_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30690));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16478_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16479_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30691));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16479_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16480_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30692));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16480_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16481_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30693));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16481_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16482_3_lut_4_lut (.I0(n52852), .I1(n135), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30694));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16482_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16473_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[2]), 
            .I3(baudrate[26]), .O(n30685));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16473_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16475_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[0]), 
            .I3(baudrate[24]), .O(n30687));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16475_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16470_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[5]), 
            .I3(baudrate[29]), .O(n30682));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16470_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16471_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[4]), 
            .I3(baudrate[28]), .O(n30683));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16471_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16472_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[3]), 
            .I3(baudrate[27]), .O(n30684));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16472_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16474_3_lut_4_lut (.I0(state[2]), .I1(n129), .I2(data[1]), 
            .I3(baudrate[25]), .O(n30686));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16474_3_lut_4_lut.LUT_INIT = 16'hfb40;
    i2c_controller i2c (.scl_enable(scl_enable), .scl(scl), .GND_net(GND_net), 
            .sda_enable(sda_enable), .sda_out(sda_out), .clk16MHz(clk16MHz), 
            .\state_7__N_4110[0] (\state_7__N_4110[0] ), .\state[3] (state_adj_5018[3]), 
            .\state[1] (state_adj_5018[1]), .\state[0] (\state[0] ), .\state[2] (state_adj_5018[2]), 
            .\saved_addr[0] (saved_addr[0]), .n7(n7), .enable_slow_N_4213(enable_slow_N_4213), 
            .n11(n11), .n29968(n29968), .data({data}), .n29967(n29967), 
            .n29965(n29965), .n29964(n29964), .n29963(n29963), .n29959(n29959), 
            .n29958(n29958), .n65606(n65606), .n6705(n6705), .n30749(n30749), 
            .n8(n8), .VCC_net(VCC_net), .n44499(n44499), .\state_7__N_4126[3] (\state_7__N_4126[3] ), 
            .enable(enable), .n10(n10), .n4(n4), .n4_adj_5(n4_adj_6), 
            .n25888(n25888), .n25930(n25930), .n44644(n44644)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (scl_enable, scl, GND_net, sda_enable, sda_out, 
            clk16MHz, \state_7__N_4110[0] , \state[3] , \state[1] , 
            \state[0] , \state[2] , \saved_addr[0] , n7, enable_slow_N_4213, 
            n11, n29968, data, n29967, n29965, n29964, n29963, 
            n29959, n29958, n65606, n6705, n30749, n8, VCC_net, 
            n44499, \state_7__N_4126[3] , enable, n10, n4, n4_adj_5, 
            n25888, n25930, n44644) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output scl_enable;
    output scl;
    input GND_net;
    output sda_enable;
    output sda_out;
    input clk16MHz;
    output \state_7__N_4110[0] ;
    output \state[3] ;
    output \state[1] ;
    output \state[0] ;
    output \state[2] ;
    output \saved_addr[0] ;
    input n7;
    output enable_slow_N_4213;
    output n11;
    input n29968;
    output [7:0]data;
    input n29967;
    input n29965;
    input n29964;
    input n29963;
    input n29959;
    input n29958;
    input n65606;
    output n6705;
    input n30749;
    input n8;
    input VCC_net;
    output n44499;
    input \state_7__N_4126[3] ;
    input enable;
    output n10;
    output n4;
    output n4_adj_5;
    output n25888;
    output n25930;
    output n44644;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire sda_out_adj_4998, i2c_clk_N_4199, scl_enable_N_4200, enable_slow_N_4212, 
        n28149, n28, n77673, n11_c, n66988, n28141;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    wire [1:0]n6774;
    
    wire n65310, n28143;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n29408;
    wire [7:0]n119;
    
    wire n28224, n29177, n5, n45056, n44799, n45054, n69207, n68997, 
        n15, n11_adj_5000, n58417, n58416, n58415, n58414, n58413, 
        n58412, n58411, n68244, n68423, n59593, n59592, n59591, 
        n59590, n59589, n11_adj_5001, n11_adj_5002, n4_c, n6698, 
        n44594, n9, n12, n4_adj_5003, n74671, n7042, n9_adj_5006, 
        n10_adj_5007;
    
    SB_LUT4 i30459_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i30459_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2555_2_lut (.I0(sda_out_adj_4998), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2555_2_lut.LUT_INIT = 16'h8888;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n28149), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i61838_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n77673));
    defparam i61838_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n11_c), .I1(n77673), .I2(n28), .I3(n66988), 
            .O(n28141));
    defparam i1_4_lut_adj_963.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1830_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6774[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1830_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i31160_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n66988));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i31160_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(\state[0] ), .I1(n7), .I2(\state[3] ), .I3(n11_c), 
            .O(n65310));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_964 (.I0(n11_c), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n66988), .O(n28143));
    defparam i1_4_lut_adj_964.LUT_INIT = 16'h0a22;
    SB_LUT4 i61988_2_lut (.I0(enable_slow_N_4213), .I1(\state_7__N_4110[0] ), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));   // verilog/i2c_controller.v(44[32:47])
    defparam i61988_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i51329_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(scl_enable_N_4200));
    defparam i51329_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29968));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29967));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29965));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29964));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29963));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29959));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29958));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n65606));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n28224), .D(n119[1]), 
            .S(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n28224), .D(n119[2]), 
            .S(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n28224), .D(n119[3]), 
            .R(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n28224), .D(n119[4]), 
            .R(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n28224), .D(n119[5]), 
            .R(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n28224), .D(n119[6]), 
            .R(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n28224), .D(n119[7]), 
            .R(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6705), .D(n5), 
            .S(n45056));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6705), .D(n44799), 
            .S(n45054));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6705), .D(n69207), 
            .S(n68997));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29408));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30749));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i30425_3_lut_4_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n44499));   // verilog/i2c_controller.v(151[5:14])
    defparam i30425_3_lut_4_lut_4_lut.LUT_INIT = 16'hfcfd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5000));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n58417), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n58416), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n58416), .I0(counter[6]), .I1(VCC_net), 
            .CO(n58417));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n58415), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n58415), .I0(counter[5]), .I1(VCC_net), 
            .CO(n58416));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n58414), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n58414), .I0(counter[4]), .I1(VCC_net), 
            .CO(n58415));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n58413), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n58413), .I0(counter[3]), .I1(VCC_net), 
            .CO(n58414));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n58412), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n58412), .I0(counter[2]), .I1(VCC_net), 
            .CO(n58413));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n58411), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n58411), .I0(counter[1]), .I1(VCC_net), 
            .CO(n58412));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n58411));
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n28143), 
            .D(n68244), .S(n65310));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4998), .C(i2c_clk), .E(n28141), 
            .D(n68423), .S(n65310));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n28224), .D(n119[0]), 
            .S(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_2057_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n59593), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2057_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n59592), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_6 (.CI(n59592), .I0(GND_net), .I1(counter2[4]), 
            .CO(n59593));
    SB_LUT4 counter2_2057_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n59591), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_5 (.CI(n59591), .I0(GND_net), .I1(counter2[3]), 
            .CO(n59592));
    SB_LUT4 counter2_2057_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n59590), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_4 (.CI(n59590), .I0(GND_net), .I1(counter2[2]), 
            .CO(n59591));
    SB_LUT4 counter2_2057_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n59589), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_3 (.CI(n59589), .I0(GND_net), .I1(counter2[1]), 
            .CO(n59590));
    SB_LUT4 counter2_2057_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n59589));
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5001));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_965 (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5002), 
            .I2(n11_c), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h2a2f;
    SB_LUT4 i62374_3_lut (.I0(n6705), .I1(n15), .I2(n11), .I3(GND_net), 
            .O(n45054));
    defparam i62374_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i62323_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5002), 
            .I2(GND_net), .I3(GND_net), .O(n44799));
    defparam i62323_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i62375_4_lut (.I0(n6705), .I1(\state[0] ), .I2(n11_adj_5001), 
            .I3(n7), .O(n45056));
    defparam i62375_4_lut.LUT_INIT = 16'h0a8a;
    SB_LUT4 i61891_4_lut (.I0(\state[3] ), .I1(n6698), .I2(n44594), .I3(n44499), 
            .O(n6705));
    defparam i61891_4_lut.LUT_INIT = 16'h5f13;
    SB_LUT4 i1_4_lut_adj_966 (.I0(n11_adj_5000), .I1(n11_adj_5002), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4126[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_966.LUT_INIT = 16'h5575;
    SB_LUT4 equal_276_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_276_i9_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6698));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\state[3] ), .I1(n6698), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_5003));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i58959_4_lut (.I0(n7), .I1(n4_adj_5003), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n74671));
    defparam i58959_4_lut.LUT_INIT = 16'hfcdd;
    SB_LUT4 i14_4_lut (.I0(n74671), .I1(n9), .I2(n7042), .I3(\state_7__N_4126[3] ), 
            .O(n28224));
    defparam i14_4_lut.LUT_INIT = 16'h35f5;
    SB_LUT4 i14965_2_lut_4_lut (.I0(n28224), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n29177));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14965_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_967 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n25888));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_967.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5006));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_968 (.I0(n15), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n25930));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_968.LUT_INIT = 16'hbbbb;
    SB_LUT4 i30570_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n44644));
    defparam i30570_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_adj_5002));   // verilog/i2c_controller.v(44[32:47])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i61985_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i61985_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n7042));   // verilog/i2c_controller.v(44[32:47])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6774[1]), 
            .I3(\state[1] ), .O(n68423));   // verilog/i2c_controller.v(44[32:47])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_adj_969 (.I0(enable), .I1(enable_slow_N_4213), 
            .I2(\state_7__N_4110[0] ), .I3(GND_net), .O(n28149));
    defparam i1_2_lut_3_lut_adj_969.LUT_INIT = 16'hbaba;
    SB_LUT4 i2_3_lut_4_lut_adj_970 (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n68244));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_970.LUT_INIT = 16'h1110;
    SB_LUT4 i62370_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(n6705), 
            .I3(\state[1] ), .O(n68997));   // verilog/i2c_controller.v(151[5:14])
    defparam i62370_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 equal_1562_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11_c));   // verilog/i2c_controller.v(151[5:14])
    defparam equal_1562_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i30520_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(GND_net), .O(n44594));
    defparam i30520_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut_adj_971 (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_c), 
            .I3(n9_adj_5006), .O(n69207));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_971.LUT_INIT = 16'hf0f4;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_5007));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_5007), .I2(counter2[0]), 
            .I3(GND_net), .O(n29408));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_972 (.I0(i2c_clk), .I1(n29408), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4199));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (PWMLimit, GND_net, \Kp[6] , \Kp[4] , \Ki[9] , 
            n349, \Ki[10] , IntegralLimit, \Kp[1] , \Kp[0] , \Ki[11] , 
            \Ki[12] , \Kp[7] , \Ki[13] , \Ki[1] , n350, \Kp[8] , 
            \Ki[0] , \Kp[2] , \Kp[9] , \Kp[10] , \Ki[2] , \Kp[3] , 
            \Ki[3] , \Kp[11] , \Kp[5] , \Ki[4] , \Kp[12] , \Kp[13] , 
            \Kp[14] , \Kp[15] , n284, n258, n356, n357, \Ki[5] , 
            \Ki[6] , \Ki[7] , \Ki[8] , n337, n313, \Ki[14] , \Ki[15] , 
            n339, n340, n358, duty, n45105, n342, n343, n344, 
            n322, n348, n359, n336, control_update, clk16MHz, reset, 
            n345, n346, n347, VCC_net, setpoint, motor_state, \PID_CONTROLLER.integral , 
            n239, n247, n467, n6, n37336, n58049, n37146, n475, 
            n30514, n30513, n30512, n30511, n30510, n30509, n30508, 
            n30507, n30506, n30505, n30503, n30501, n30500, n30499, 
            n30498, n30497, n30496, n30495, n30494, n30493, n30488, 
            n30487, n30479, deadband, n29773, n460, n65754, n22, 
            n351, n38, \control_mode[5] , \control_mode[0] , \control_mode[1] , 
            \control_mode[6] , \control_mode[7] , n110, n9, n16, n34707, 
            n20, n25, n33, n37, n41, n22_adj_1, n486, n35808, 
            n24, n36173, n291, n25794, n352, n299, n38_adj_2, 
            n8, n25_adj_3, n10, n39, n20419, n20420, n56, n40, 
            n353, n354, n20466, n355, n21, n37_adj_4, n57846, 
            n20493, n20465) /* synthesis syn_module_defined=1 */ ;
    input [23:0]PWMLimit;
    input GND_net;
    input \Kp[6] ;
    input \Kp[4] ;
    input \Ki[9] ;
    input n349;
    input \Ki[10] ;
    input [23:0]IntegralLimit;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Kp[7] ;
    input \Ki[13] ;
    input \Ki[1] ;
    output n350;
    input \Kp[8] ;
    input \Ki[0] ;
    input \Kp[2] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Ki[2] ;
    input \Kp[3] ;
    input \Ki[3] ;
    input \Kp[11] ;
    input \Kp[5] ;
    input \Ki[4] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    output n284;
    output n258;
    output n356;
    output n357;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    output n337;
    output n313;
    input \Ki[14] ;
    input \Ki[15] ;
    output n339;
    output n340;
    output n358;
    output [23:0]duty;
    output n45105;
    output n342;
    output n343;
    output n344;
    output n322;
    output n348;
    output n359;
    output n336;
    output control_update;
    input clk16MHz;
    input reset;
    output n345;
    output n346;
    input n347;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output [23:0]\PID_CONTROLLER.integral ;
    output n239;
    output n247;
    output n467;
    input n6;
    input n37336;
    input n58049;
    input n37146;
    output n475;
    input n30514;
    input n30513;
    input n30512;
    input n30511;
    input n30510;
    input n30509;
    input n30508;
    input n30507;
    input n30506;
    input n30505;
    input n30503;
    input n30501;
    input n30500;
    input n30499;
    input n30498;
    input n30497;
    input n30496;
    input n30495;
    input n30494;
    input n30493;
    input n30488;
    input n30487;
    input n30479;
    input [23:0]deadband;
    input n29773;
    output n460;
    output n65754;
    input n22;
    output n351;
    input n38;
    input \control_mode[5] ;
    input \control_mode[0] ;
    input \control_mode[1] ;
    input \control_mode[6] ;
    input \control_mode[7] ;
    input n110;
    input n9;
    output n16;
    input n34707;
    output n20;
    input n25;
    input n33;
    input n37;
    input n41;
    input n22_adj_1;
    output n486;
    input n35808;
    output n24;
    input n36173;
    output n291;
    input n25794;
    output n352;
    output n299;
    output n38_adj_2;
    output n8;
    input n25_adj_3;
    input n10;
    input n39;
    input n20419;
    input n20420;
    input n56;
    input n40;
    output n353;
    output n354;
    output n20466;
    output n355;
    input n21;
    input n37_adj_4;
    output n57846;
    input n20493;
    output n20465;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    wire [23:0]n207;
    
    wire n454, n323, n688, n761;
    wire [23:0]n1_adj_4996;
    wire [23:0]n285;
    
    wire n58319, n58522;
    wire [11:0]n19061;
    
    wire n58523;
    wire [12:0]n18698;
    
    wire n250, n58521, n110_c, n41_c, n58320, n834, n907, n527, 
        n980, n101, n600, n32, n58318, n183, n58317, n673, n746, 
        n58316, n174, n256, n247_c, n819, n329, n402, n320, 
        n892, n475_c, n548, n965, n621, n694, n767, n1038, n840, 
        n1111;
    wire [23:0]n233;
    wire [23:0]n310;
    
    wire n80, n11, n153, n226, n393, n299_c, n466, n86, n17_adj_4435, 
        n159, n372, n445, n518, n591, n232, n305_adj_4436, n539, 
        n58315, n378, n451, n524, n597, n664, n670, n743, n737, 
        n816, n810, n883, n956, n1029, n1102, n58214;
    wire [43:0]n360;
    wire [47:0]n46;
    
    wire n58215, n889, n962, n77, n8_adj_4438, n150, n1035, n1108, 
        n223_adj_4439, n296, n369, n442, n515, n588, n125, n661, 
        n56_c, n198, n734, n807, n880, n953, n1026, n1099, n271, 
        n57894, n70879, n74, n5_adj_4442, n344_adj_4443, n147;
    wire [2:0]n20468;
    
    wire n4_adj_4444;
    wire [4:0]n20370;
    
    wire n417, n347_c, n6_adj_4445, n66283, n220, n293_adj_4446, 
        n366, n439, n70875, n512, n585, n658, n731, n62, n804, 
        n877, n950, n57908, n58123, n1023, n490, n1096, n70865, 
        n79606, n70869, n8_adj_4447, n6_adj_4448, n68674, n177, 
        n58520, n58314, n35, n104;
    wire [23:0]n455;
    
    wire n78630, counter_31__N_3714, n116, n47, n612, n41_adj_4450, 
        n189, n183_adj_4452, n256_adj_4453, n262, n58176, n329_adj_4454, 
        n335, n58213, n402_adj_4455, n58212, n408, n58177, n475_adj_4456, 
        n58211, n481, n554, n548_adj_4457, n621_adj_4458, n627, 
        n700, n694_adj_4459, n11880, n74615, n4734, n78777, n767_adj_4460, 
        n58210, n840_adj_4461, n58175, n107, n180, n253, n326, 
        n399, n472, n545, n618, n691;
    wire [23:0]n535;
    
    wire n78780, n764, n837, n58174, n58209, n58208, n58207, n685, 
        n78930, n58173, n78906, n78894, n78888, n58206, n58205, 
        n78882, n78876, n78870, n58172, n58204, n78858, n58203, 
        n877_adj_4464, n448, n58202, n521, n594, n667, n740, n950_adj_4465, 
        n813, n886, n959, n758, n1032, n1105, n910, n831, n1023_adj_4466, 
        n58201, n58200, n74604, n78717, n78720, n78846, n74603, 
        n78711, n78714, n78816, n904, n75342, n74602, n78705, 
        n75364, n78708, n58199, n75267, n58198;
    wire [0:0]n12496;
    wire [21:0]n13003;
    
    wire n59846, n59845, n59844, n59843, n59842, n59841, n59840, 
        n75291, n59839, n59838, n59837, n59836, n59835, n59834, 
        n74601, n78699, n59833, n78702, n59832, n59831, n59830, 
        n59829, n78696, n78690, n59828, n59827, n59826, n78684, 
        n59825;
    wire [20:0]n13968;
    
    wire n59824, n59823, n59822, n59821, n78678, n78672, n59820, 
        n59819, n59818, n59817, n59816, n78666, n59815, n59814, 
        n59813, n59812, n78660, n59811, n59810, n59809, n59808, 
        n59807, n59806, n59805, n59804;
    wire [19:0]n14846;
    
    wire n59803, n59802, n59801, n59800, n59799, n59798, n59797, 
        n59796, n59795, n59794, n59793, n59792, n59791, n59790;
    wire [0:0]n11920;
    wire [21:0]n12379;
    
    wire n58903, n59789, n59788, n59787, n59786, n59785, n59784, 
        n58902, n58901;
    wire [10:0]n19372;
    wire [9:0]n19635;
    
    wire n59783, n59782, n59781, n59780, n59779, n59778, n59777, 
        n58900, n59776, n58899, n58898, n59775, n59774;
    wire [18:0]n15642;
    
    wire n59773, n58897, n58896, n1096_adj_4475, n58895, n59772, 
        n59771, n59770, n59769, n58894, n59768, n396, n469_adj_4476, 
        n59767, n542, n615, n688_adj_4477, n761_adj_4478, n834_adj_4479, 
        n59766, n907_adj_4480, n59765, n59764, n58893, n59763, n980_adj_4481, 
        n125_adj_4482, n59762, n59761, n198_adj_4483, n271_adj_4484, 
        n59760, n344_adj_4485, n59759, n417_adj_4486, n58892;
    wire [3:0]n20462;
    wire [4:0]n20416;
    
    wire n375, n59758, n204, n302_adj_4488, n59757;
    wire [1:0]n20499;
    wire [2:0]n20490;
    
    wire n804_adj_4490, n58891, n131, n62_adj_4491, n229, n59756, 
        n156, n59755, n14_adj_4492, n83;
    wire [17:0]n16360;
    
    wire n59754, n59753, n59752, n59751, n1108_adj_4493, n59750, 
        n1035_adj_4494, n59749, n962_adj_4495, n59748, n490_adj_4496, 
        n889_adj_4497, n59747, n70829, n70833, n816_adj_4498, n59746, 
        n731_adj_4499, n58890, n743_adj_4500, n59745, n70831, n670_adj_4501, 
        n59744, n57998, n70839, n4_adj_4502, n597_adj_4503, n59743, 
        n8_adj_4504, n524_adj_4505, n59742, n658_adj_4506, n58889, 
        n6_adj_4507, n69074, n451_adj_4508, n59741, n378_adj_4509, 
        n59740, n305_adj_4510, n59739, n585_adj_4512, n58888, n232_adj_4513, 
        n59738, n512_adj_4514, n58887, n159_adj_4515, n59737, n17_adj_4516, 
        n86_adj_4517, n439_adj_4519, n58886;
    wire [8:0]n19854;
    
    wire n770, n59736, n697, n59735, n366_adj_4521, n58885, n624, 
        n59734, n101_adj_4522, n32_adj_4523, n551, n59733, n478, 
        n59732, n293_adj_4524, n58884, n174_adj_4525, n58197, n405, 
        n59731, n247_adj_4527, n220_adj_4528, n58883, n320_adj_4529, 
        n393_adj_4530, n466_adj_4531, n332_adj_4532, n59730, n539_adj_4533, 
        n259, n59729, n612_adj_4534, n186, n59728, n685_adj_4535, 
        n44, n113, n147_adj_4537, n58882, n758_adj_4538;
    wire [16:0]n17004;
    
    wire n59727, n59726, n74600, n78693, n59725, n831_adj_4539, 
        n904_adj_4540, n1111_adj_4541, n59724, n977, n1050, n1038_adj_4542, 
        n59723, n98, n965_adj_4543, n59722, n29, n171, n892_adj_4544, 
        n59721, n819_adj_4545, n59720, n244_adj_4546, n317_adj_4548, 
        n390_adj_4549, n463, n746_adj_4550, n59719, n673_adj_4551, 
        n59718, n536, n609, n600_adj_4552, n59717, n682, n755, 
        n527_adj_4553, n59716, n828, n454_adj_4555, n59715, n381, 
        n59714, n901, n74599, n78687, n974, n308_adj_4557, n59713, 
        n235_adj_4559, n59712, n1047, n162, n59711, n74598, n78681, 
        n1120, n122, n20_adj_4561, n89;
    wire [15:0]n17578;
    
    wire n59710, n53, n59709, n195, n1114, n59708, n268, n5_adj_4563, 
        n74_adj_4564, n1041, n59707, n341, n968, n59706, n895, 
        n59705, n414, n822, n59704, n487, n560, n749, n59703, 
        n676, n59702, n74597, n78675, n603, n59701, n530, n59700, 
        n457, n59699, n384_adj_4568, n59698, n311_adj_4569, n59697, 
        n238_adj_4570, n59696, n165, n59695, n23_adj_4574, n92;
    wire [9:0]n19776;
    wire [8:0]n19972;
    
    wire n770_adj_4575, n58881;
    wire [7:0]n20033;
    
    wire n700_adj_4576, n59694, n697_adj_4577, n58880, n627_adj_4578, 
        n59693, n95, n554_adj_4579, n59692, n26, n168, n481_adj_4580, 
        n59691, n408_adj_4582, n59690, n241_adj_4583, n335_adj_4584, 
        n59689, n262_adj_4585, n59688, n189_adj_4586, n59687, n47_adj_4587, 
        n116_adj_4588;
    wire [14:0]n18086;
    
    wire n59686, n1117, n59685, n1044, n59684, n314_adj_4590, n971, 
        n59683, n898, n59682, n825, n59681, n752, n59680, n679, 
        n59679, n606, n59678, n533, n59677, n460_c, n59676, n387_adj_4591, 
        n59675, n314_adj_4592, n59674, n241_adj_4593, n59673, n168_adj_4594, 
        n59672, n26_adj_4595, n95_adj_4596;
    wire [13:0]n18532;
    
    wire n1120_adj_4597, n59671, n1047_adj_4598, n59670, n974_adj_4599, 
        n59669, n901_adj_4600, n59668, n74596, n78669;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n387_adj_4601, n460_adj_4602, n828_adj_4604, n59667, n755_adj_4607, 
        n59666, n682_adj_4608, n59665, n74595, n78663, n624_adj_4609, 
        n58879, n609_adj_4610, n59664, n536_adj_4611, n59663, n463_adj_4612, 
        n59662, n390_adj_4613, n59661, n317_adj_4614, n59660, n244_adj_4615, 
        n59659, n171_adj_4616, n59658, n29_adj_4617, n98_adj_4618;
    wire [6:0]n20176;
    
    wire n630, n59657, n551_adj_4619, n58878, n557, n59656, n484, 
        n59655, n478_adj_4620, n58877, n411, n59654, n405_adj_4621, 
        n58876, n338, n59653, n265, n59652, n332_adj_4622, n58875, 
        n259_adj_4623, n58874, n192, n59651, n186_adj_4624, n58873, 
        n50, n119, n44_adj_4625, n113_adj_4626;
    wire [12:0]n18920;
    
    wire n1050_adj_4627, n59650, n977_adj_4628, n59649, n59648, n59647, 
        n59646, n59645, n59644, n59643, n59642, n59641, n533_adj_4630, 
        n606_adj_4631, n679_adj_4632, n752_adj_4633, n825_adj_4634, 
        n898_adj_4635, n59640, n971_adj_4636, n1044_adj_4637, n1117_adj_4638, 
        n59639, n59638;
    wire [11:0]n19254;
    
    wire n59637, n59636, n59635, n59634, n59633, n45170;
    wire [23:0]n1_adj_4997;
    
    wire n615_adj_4645, n59632;
    wire [20:0]n13441;
    
    wire n58850, n542_adj_4646, n59631, n58849, n58848, n58847, 
        n58846, n910_adj_4647, n58438, n58845, n58844, n469_adj_4648, 
        n59630, n1099_adj_4649, n58843, n837_adj_4650, n58437, n1026_adj_4651, 
        n58842, n764_adj_4652, n58436, n953_adj_4653, n58841, n691_adj_4654, 
        n58435, n880_adj_4655, n58840, n78654, n618_adj_4656, n58434, 
        n807_adj_4657, n58839, n734_adj_4658, n58838, n661_adj_4659, 
        n58837, n545_adj_4660, n58433, n588_adj_4661, n58836, n472_adj_4662, 
        n58432, n515_adj_4663, n58835, n399_adj_4664, n58431, n442_adj_4665, 
        n58834, n326_adj_4666, n58430, n369_adj_4667, n58833, n296_adj_4668, 
        n58832, n223_adj_4669, n58831, n150_adj_4670, n58830, n396_adj_4671, 
        n59629, n8_adj_4672, n77_adj_4673, n253_adj_4674, n58429;
    wire [19:0]n14365;
    
    wire n58829, n58828, n180_adj_4675, n58428, n323_adj_4676, n59628, 
        n58827, n38_c, n107_adj_4677, n58826, n58825, n58824, n1102_adj_4680, 
        n58823, n1029_adj_4681, n58822, n956_adj_4683, n58821, n883_adj_4684, 
        n58820, n250_adj_4685, n59627, n810_adj_4686, n58819, n737_adj_4687, 
        n58818, n177_adj_4688, n59626, n664_adj_4689, n58817, n591_adj_4690, 
        n58816, n518_adj_4691, n58815, n445_adj_4692, n58814, n372_adj_4693, 
        n58813, n299_adj_4694, n58812, n35_adj_4695, n104_adj_4696, 
        n226_adj_4697, n58811, n153_adj_4698, n58810, n11_adj_4699, 
        n80_adj_4700;
    wire [5:0]n20287;
    
    wire n560_adj_4701, n59625, n487_adj_4702, n59624, n414_adj_4703, 
        n59623, n41_adj_4705, n39_c, n45, n43, n37_c, n29_adj_4709, 
        n31, n74663, n78927, n21_adj_4711, n23_adj_4712, n25_adj_4713, 
        n17_adj_4714, n19_adj_4715, n9_adj_4716;
    wire [18:0]n15204;
    
    wire n58788, n58787, n35_adj_4719, n33_c, n11_adj_4721, n15_adj_4722, 
        n27, n13_adj_4723, n58786, n58785, n58784, n41_adj_4727, 
        n39_adj_4728, n45_adj_4729, n43_adj_4730, n37_adj_4731, n1105_adj_4732, 
        n58783, n29_adj_4733, n1032_adj_4734, n58782, n959_adj_4735, 
        n58781, n31_adj_4736, n23_adj_4737, n25_adj_4738, n35_adj_4739, 
        n11_adj_4740, n886_adj_4741, n58780, n13_adj_4742, n813_adj_4743, 
        n58779, n740_adj_4744, n58778, n27_adj_4745, n58196, n341_adj_4746, 
        n59622, n15_adj_4747, n33_adj_4748, n9_adj_4749, n17_adj_4750, 
        n19_adj_4751, n21_adj_4752, n105, n25796, n667_adj_4754, n58777, 
        n594_adj_4755, n58776, n521_adj_4756, n58775, n448_adj_4757, 
        n58774, n75495, n75457, n12_adj_4758, n10_adj_4759, n30, 
        n375_adj_4760, n58773, n302_adj_4761, n58772, n75511, n76409, 
        n76399, n77387, n76794, n77503, n16_adj_4762, n6_adj_4763, 
        n77109, n229_adj_4764, n58771, n156_adj_4765, n58770, n77110, 
        n8_adj_4766, n24_adj_4767, n75421, n75410, n76900, n75809, 
        n4_adj_4768, n14_adj_4769, n83_adj_4770, n92_adj_4772, n23_adj_4773, 
        n268_adj_4775, n59621, n165_adj_4776, n195_adj_4777, n59620, 
        n238_adj_4778, n77107, n311_adj_4779, n77108, n53_adj_4780, 
        n122_adj_4781, n384_adj_4782, n75444, n457_adj_4783, n75440, 
        n77447, n75811, n77607, n530_adj_4785, n603_adj_4786, n77608, 
        n676_adj_4787;
    wire [10:0]n19538;
    
    wire n59619, n749_adj_4788, n822_adj_4791, n895_adj_4793, n968_adj_4794, 
        n77557, n59618, n59617, n1041_adj_4795, n59616, n75427, 
        n59615, n59614, n77409, n75817, n59613, n77411, n59612, 
        n59611, n59610, n1114_adj_4798, n119_adj_4799, n59609, n50_adj_4800, 
        n59608, n59607, n192_adj_4802, n265_adj_4803, n6_adj_4804, 
        n59606;
    wire [7:0]n20130;
    
    wire n58749, n58748, n59605, n59604, n58747, n338_adj_4806, 
        n58746, n411_adj_4807, n484_adj_4808, n59603, n557_adj_4809, 
        n58745, n630_adj_4810, n59602, n58744, n59601, n58743, n59600, 
        n59599, n58742, n59598, n59597, n59596;
    wire [17:0]n15963;
    
    wire n58741, n59595, n59594, n58740, n89_adj_4818, n20_adj_4819, 
        n58739, n58738, n162_adj_4821, n43_adj_4822, n235_adj_4823, 
        n58737, n39_adj_4824, n58736, n58195, n58735, n58194, n58382, 
        n58734, n58171, n58381, n308_adj_4827, n4_adj_4828, n6_adj_4829, 
        n8_adj_4831, n381_adj_4832, n75597, n77443, n58733, n77444, 
        n77324, n58732, n58380, n58731, n58730, n58729, n58379, 
        n58193, n58728, n58378, n58727, n58726, n58725, n58377, 
        n58724, n58376, n27_adj_4835, n58375, n58374, n29_adj_4836, 
        n31_adj_4837, n35_adj_4838, n23_adj_4839, n75572, n75558, 
        n28, n30_adj_4842, n58373, n58372, n58371, n58370, n58369, 
        n58368;
    wire [16:0]n16646;
    
    wire n58704, n58703, n58367, n58702, n58366, n58192, n58701, 
        n58700, n58365, n58699, n58364, n58698, n58191, n58170, 
        n58169, n58697, n58363, n58168, n58696, n26_adj_4843, n34, 
        n58695, n58362, n24_adj_4845, n75556, n77445, n58694, n77446, 
        n58693, n58190, n58692, n58361, n77322, n58360, n58691, 
        n58690, n77177, n58189, n75566, n77343, n58689, n75807, 
        n58688, n47_adj_4849, n58359, n77487;
    wire [23:0]n48;
    
    wire n58358, n77488, n58357, n58188, n37_adj_4851, n35_adj_4852, 
        n58356, n13_adj_4853, n15_adj_4854, n19_adj_4855, n17_adj_4856, 
        n7_adj_4857, n58355, n58354, n11_adj_4859, n5_adj_4860, n75140, 
        n58353, n58187, n8_adj_4861;
    wire [6:0]n20254;
    
    wire n58669, n58668, n58667, n58666, n6_adj_4862, n58665, n58352, 
        n58664, n58663, n16_adj_4863, n4_adj_4865;
    wire [15:0]n17257;
    
    wire n58662, n58661, n58660, n58351, n58186, n58350, n77034, 
        n58659, n58658, n58657, n58349, n58656, n58185, n58348, 
        n77035, n75136, n58347, n58655, n58654, n58653, n58652, 
        n58346, n58651, n75134, n77331, n58650, n58649, n58648, 
        n58184, n58647, n58345, n75859, n58344, n77568, n77569, 
        n58183, n58343, n58342, n58341, n58340, n58339, n58338, 
        n58337, n74481, n58182, n58336, n58335, n58334, n58181, 
        n41_adj_4868, n39_adj_4869, n29_adj_4870, n58333, n31_adj_4871, 
        n58332, n33_adj_4872;
    wire [14:0]n17800;
    
    wire n58629, n58628, n27_adj_4873, n75126, n30_adj_4874, n28_adj_4875, 
        n58627, n38_adj_4876, n58626, n58625, n58624, n77030, n77031, 
        n75120, n58623, n58622, n75118, n77457, n58621, n75861, 
        n77597, n58620, n77598, n77548, n58619, n58618, n58180, 
        n58617, n58179, n58178, n58616, n58331, n7054, n35_adj_4877, 
        n7_adj_4878, n58615, n58330, n9_adj_4879, n31_adj_4880, n58329, 
        n23_adj_4881, n58328, n25_adj_4882, n33_adj_4883, n29_adj_4884, 
        n27_adj_4885, n17_adj_4886, n19_adj_4887, n21_adj_4888, n11_adj_4889, 
        n13_adj_4890, n15_adj_4891, n75158, n76155, n76678, n76676, 
        n75162, n75051, n12_adj_4892, n4_adj_4893, n77036, n77037, 
        n10_adj_4894, n30_adj_4896, n75154, n75152, n76908, n75857, 
        n8_adj_4897, n6_adj_4898, n58327;
    wire [5:0]n20348;
    
    wire n58598, n16_adj_4899, n58597, n75200, n77455, n77456, n77304, 
        n58326, n58596, n58325, n58595, n58594, n77103, n58324, 
        n58593;
    wire [13:0]n18279;
    
    wire n58592, n58323, n77421, n75855, n77423, n58591, n37_adj_4903, 
        n58590, n58236, n35_adj_4904, n58322, n41_adj_4905, n58235, 
        n58589, n29_adj_4906, n58588, n31_adj_4907, n58321, n58587, 
        n58586, n58234, n58585, n58584, n33_adj_4908, n4_adj_4909, 
        n58583, n58582, n76906, n23_adj_4911, n58581, n58580, n59529, 
        n59528, n58579, n58233, n58232, n58231, n58230, n59527, 
        n27_adj_4912, n17_adj_4913, n19_adj_4914, n58229, n75075, 
        n58228, n21_adj_4915, n58227, n58563, n58562, n59526, n58561, 
        n58226, n59525, n13_adj_4916, n58560, n75251, n15_adj_4917, 
        n59524, n58559, n59523, n76201, n76706, n59522, n58558, 
        n59521, n58557, n58556, n58555, n58225, n59520, n76704, 
        n75237, n59519, n58554, n58553, n59518, n58224, n58552, 
        n77060, n59517, n75225, n58551, n58223, n18_adj_4921, n16_adj_4922, 
        n58222, n58221, n58220, n58219, n74594, n78657, n58218, 
        n58536, n36, n75235, n58535, n58534, n58533, n77061, n58532, 
        n75227, n58217, n58531, n58530, n58216, n58529, n58528, 
        n77453, n75843, n58527, n42, n58526, n75148, n58525, n79219, 
        n58524, n44_adj_4924, n76910, n14_adj_4925, n12_adj_4926, 
        n22_adj_4927, n77451, n77452, n77312, n77127, n77595, n75841, 
        n77643, n77644, n76911, n77642, n44588, n74632, n78903, 
        n7052, n25756, n67040, n75081, n12_adj_4928, n10_adj_4929, 
        n30_adj_4930, n75112, n76075, n76071, n77301, n76628, n77475, 
        n6_adj_4931, n77026, n77027, n16_adj_4932, n8_adj_4933, n24_adj_4934, 
        n75095, n75057, n76914, n75869, n4_adj_4935, n76626, n76627, 
        n75077, n77265, n75871, n77532, n77533, n77478, n75065, 
        n77221, n75877, n77424, n74593, n78651, n4_adj_4936, n68521, 
        n25798, n6_adj_4937, n75406, n75338, n6_adj_4938, n74631, 
        n78891, n74630, n78885, n74629, n78879, n74628, n78873, 
        n74627, n78867, n74626, n78855, n25754, n74592, n78627, 
        n74624, n74625, n78843, n71340, n23_adj_4940, n22_adj_4941, 
        n26_adj_4942, n41_adj_4943, n39_adj_4944, n45_adj_4945, n43_adj_4946, 
        n23_adj_4947, n25_adj_4948, n29_adj_4949, n31_adj_4950, n35_adj_4951, 
        n33_adj_4952, n11_adj_4953, n13_adj_4954, n15_adj_4955, n27_adj_4956, 
        n9_adj_4957, n17_adj_4958, n19_adj_4959, n75316, n75305, n12_adj_4961, 
        n10_adj_4962, n30_adj_4963, n76269, n76259, n77355, n76726, 
        n77493, n16_adj_4965, n77095, n77096, n8_adj_4966, n24_adj_4967, 
        n75271, n76904, n75829, n4_adj_4968, n77093, n77094, n75297, 
        n77481, n75831, n77593, n77594, n77553, n75275, n77417, 
        n75837, n77419, n4_adj_4969, n41_adj_4970, n39_adj_4971, n45_adj_4972, 
        n43_adj_4973, n37_adj_4974, n29_adj_4975, n31_adj_4976, n23_adj_4977, 
        n25_adj_4978, n35_adj_4979, n11_adj_4980, n13_adj_4981, n15_adj_4982, 
        n27_adj_4983, n33_adj_4984, n9_adj_4985, n17_adj_4986, n19_adj_4987, 
        n21_adj_4988, n75388, n75376, n12_adj_4989, n10_adj_4990, 
        n30_adj_4991, n76333, n76323, n77371, n76760, n77499, n16_adj_4992, 
        n77101, n77102, n8_adj_4993, n24_adj_4994, n75346, n76902, 
        n75819, n4_adj_4995, n77099, n77100, n75370, n77449, n75821, 
        n77591, n77592, n77555, n75350, n77413, n75827, n77415, 
        n78813;
    
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[6]), 
            .I3(n58319), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_5 (.CI(n58522), .I0(n19061[2]), .I1(n323), .CO(n58523));
    SB_LUT4 add_6481_4_lut (.I0(GND_net), .I1(n19061[1]), .I2(n250), .I3(n58521), 
            .O(n18698[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_4 (.CI(n58521), .I0(n19061[1]), .I1(n250), .CO(n58522));
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n58319), .I0(GND_net), .I1(n1_adj_4996[6]), 
            .CO(n58320));
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[5]), 
            .I3(n58318), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n58318), .I0(GND_net), .I1(n1_adj_4996[5]), 
            .CO(n58319));
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[4]), 
            .I3(n58317), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n58317), .I0(GND_net), .I1(n1_adj_4996[4]), 
            .CO(n58318));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[3]), 
            .I3(n58316), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n58316), .I0(GND_net), .I1(n1_adj_4996[3]), 
            .CO(n58317));
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n247_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n356));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n11));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n299_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4435));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4436));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[2]), 
            .I3(n58315), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n313));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n339));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_25_3 (.CI(n58214), .I0(n360[1]), .I1(n46[1]), .CO(n58215));
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n340));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n357));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n357), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4438));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31029_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45105));   // verilog/motorControl.v(42[14] 73[8])
    defparam i31029_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n342));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n343));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n348));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut (.I0(n207[23]), .I1(\Kp[2] ), .I2(n57894), .I3(n207[22]), 
            .O(n70879));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n358));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n358), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4442));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4443));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_944 (.I0(n207[22]), .I1(n20468[1]), .I2(n4_adj_4444), 
            .I3(\Kp[3] ), .O(n20370[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_944.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_945 (.I0(n20468[1]), .I1(n6_adj_4445), .I2(n347_c), 
            .I3(n66283), .O(n20370[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4446));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i43863_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n57894));   // verilog/motorControl.v(61[20:26])
    defparam i43863_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(n70875), .I1(n207[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4444));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i43924_4_lut (.I0(n20468[1]), .I1(\Kp[3] ), .I2(n4_adj_4444), 
            .I3(n207[22]), .O(n6_adj_4445));   // verilog/motorControl.v(61[20:26])
    defparam i43924_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i40_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n70875));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i55580_3_lut (.I0(n207[23]), .I1(n70875), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n66283));   // verilog/motorControl.v(61[20:26])
    defparam i55580_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44055_3_lut (.I0(n207[23]), .I1(n57908), .I2(n58123), .I3(GND_net), 
            .O(n20468[1]));   // verilog/motorControl.v(61[20:26])
    defparam i44055_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_946 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n58123), 
            .I3(n207[22]), .O(n70865));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_545_2_lut (.I0(n20468[1]), .I1(n66283), .I2(GND_net), 
            .I3(GND_net), .O(n79606));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_545_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n57908), .I1(n70865), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n70869));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h9666;
    SB_LUT4 i43932_4_lut (.I0(n79606), .I1(\Kp[4] ), .I2(n6_adj_4445), 
            .I3(n207[22]), .O(n8_adj_4447));   // verilog/motorControl.v(61[20:26])
    defparam i43932_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n336));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43885_4_lut (.I0(n20468[1]), .I1(\Kp[3] ), .I2(n70875), .I3(n207[23]), 
            .O(n6_adj_4448));   // verilog/motorControl.v(61[20:26])
    defparam i43885_4_lut.LUT_INIT = 16'he800;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n58315), .I0(GND_net), .I1(n1_adj_4996[2]), 
            .CO(n58316));
    SB_LUT4 i1_4_lut_adj_948 (.I0(n6_adj_4448), .I1(n8_adj_4447), .I2(n70869), 
            .I3(n66283), .O(n68674));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 add_6481_3_lut (.I0(GND_net), .I1(n19061[0]), .I2(n177), .I3(n58520), 
            .O(n18698[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_3 (.CI(n58520), .I0(n19061[0]), .I1(n177), .CO(n58521));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[1]), 
            .I3(n58314), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n18698[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n46[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n78630), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_CARRY add_6481_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n58520));
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4450));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4452));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4453));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n58314), .I0(GND_net), .I1(n1_adj_4996[1]), 
            .CO(n58315));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n46[0]), .CO(n58214));
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n58176), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4996[0]), 
            .CO(n58314));
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n58213), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4455));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n58212), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_24 (.CI(n58212), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n58213));
    SB_CARRY sub_15_add_2_11 (.CI(n58176), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n58177));
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4456));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n58211), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4457));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4458));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4459));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_23 (.CI(n58211), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n58212));
    SB_LUT4 n11880_bdd_4_lut_62918 (.I0(n11880), .I1(n74615), .I2(setpoint[13]), 
            .I3(n4734), .O(n78777));
    defparam n11880_bdd_4_lut_62918.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4460));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n58210), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4461));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n58175), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78777_bdd_4_lut (.I0(n78777), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4734), .O(n78780));
    defparam n78777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_10 (.CI(n58175), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n58176));
    SB_CARRY add_16_22 (.CI(n58210), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n58211));
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n58174), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n58174), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n58175));
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n58209), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n58209), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n58210));
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n58208), .O(n239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_20 (.CI(n58208), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n58209));
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n58207), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n78930), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n58173), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_19 (.CI(n58207), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n58208));
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n78906), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n78894), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n78888), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n58206), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_18 (.CI(n58206), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n58207));
    SB_CARRY sub_15_add_2_8 (.CI(n58173), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n58174));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n58205), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n78882), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n78876), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_16_17 (.CI(n58205), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n58206));
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n78870), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n58172), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n58204), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n78858), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_16_16 (.CI(n58204), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n58205));
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n58203), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_15 (.CI(n58203), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n58204));
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4464));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_7 (.CI(n58172), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n58173));
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n58202), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_14 (.CI(n58202), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n58203));
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4465));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4466));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n58201), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_13 (.CI(n58201), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n58202));
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n58200), .O(n247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11880_bdd_4_lut_62889 (.I0(n11880), .I1(n74604), .I2(setpoint[12]), 
            .I3(n4734), .O(n78717));
    defparam n11880_bdd_4_lut_62889.LUT_INIT = 16'he4aa;
    SB_LUT4 n78717_bdd_4_lut (.I0(n78717), .I1(n535[12]), .I2(n467), .I3(n4734), 
            .O(n78720));
    defparam n78717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n78846), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n11880_bdd_4_lut_62840 (.I0(n11880), .I1(n74603), .I2(setpoint[11]), 
            .I3(n4734), .O(n78711));
    defparam n11880_bdd_4_lut_62840.LUT_INIT = 16'he4aa;
    SB_CARRY add_16_12 (.CI(n58200), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n58201));
    SB_LUT4 n78711_bdd_4_lut (.I0(n78711), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4734), .O(n78714));
    defparam n78711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n78816), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59507_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n75342));
    defparam i59507_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n11880_bdd_4_lut_62835 (.I0(n11880), .I1(n74602), .I2(setpoint[10]), 
            .I3(n4734), .O(n78705));
    defparam n11880_bdd_4_lut_62835.LUT_INIT = 16'he4aa;
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n78780), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n78720), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n78714), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i59529_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n75364));
    defparam i59529_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n78705_bdd_4_lut (.I0(n78705), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4734), .O(n78708));
    defparam n78705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n58199), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n58199), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n58200));
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n78708), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i59432_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n75267));
    defparam i59432_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n58198), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n336), .I1(n13003[21]), .I2(GND_net), 
            .I3(n59846), .O(n12496[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n13003[20]), .I2(GND_net), 
            .I3(n59845), .O(n46[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_23 (.CI(n59845), .I0(n13003[20]), .I1(GND_net), 
            .CO(n59846));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n13003[19]), .I2(GND_net), 
            .I3(n59844), .O(n46[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_22 (.CI(n59844), .I0(n13003[19]), .I1(GND_net), 
            .CO(n59845));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n13003[18]), .I2(GND_net), 
            .I3(n59843), .O(n46[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_21 (.CI(n59843), .I0(n13003[18]), .I1(GND_net), 
            .CO(n59844));
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n13003[17]), .I2(GND_net), 
            .I3(n59842), .O(n46[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n59842), .I0(n13003[17]), .I1(GND_net), 
            .CO(n59843));
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n13003[16]), .I2(GND_net), 
            .I3(n59841), .O(n46[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_19 (.CI(n59841), .I0(n13003[16]), .I1(GND_net), 
            .CO(n59842));
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n13003[15]), .I2(GND_net), 
            .I3(n59840), .O(n46[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_18 (.CI(n59840), .I0(n13003[15]), .I1(GND_net), 
            .CO(n59841));
    SB_LUT4 i59456_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n75291));
    defparam i59456_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n13003[14]), .I2(GND_net), 
            .I3(n59839), .O(n46[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_17 (.CI(n59839), .I0(n13003[14]), .I1(GND_net), 
            .CO(n59840));
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n13003[13]), .I2(n1096), 
            .I3(n59838), .O(n46[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_16 (.CI(n59838), .I0(n13003[13]), .I1(n1096), 
            .CO(n59839));
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n13003[12]), .I2(n1023), 
            .I3(n59837), .O(n46[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_15 (.CI(n59837), .I0(n13003[12]), .I1(n1023), 
            .CO(n59838));
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n13003[11]), .I2(n950), 
            .I3(n59836), .O(n46[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_14 (.CI(n59836), .I0(n13003[11]), .I1(n950), 
            .CO(n59837));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n13003[10]), .I2(n877), 
            .I3(n59835), .O(n46[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_13 (.CI(n59835), .I0(n13003[10]), .I1(n877), 
            .CO(n59836));
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n13003[9]), .I2(n804), 
            .I3(n59834), .O(n46[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_12 (.CI(n59834), .I0(n13003[9]), .I1(n804), 
            .CO(n59835));
    SB_LUT4 n11880_bdd_4_lut_62830 (.I0(n11880), .I1(n74601), .I2(setpoint[9]), 
            .I3(n4734), .O(n78699));
    defparam n11880_bdd_4_lut_62830.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n13003[8]), .I2(n731), 
            .I3(n59833), .O(n46[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n78702), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY mult_24_add_1225_11 (.CI(n59833), .I0(n13003[8]), .I1(n731), 
            .CO(n59834));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n13003[7]), .I2(n658), 
            .I3(n59832), .O(n46[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n59832), .I0(n13003[7]), .I1(n658), 
            .CO(n59833));
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n13003[6]), .I2(n585), 
            .I3(n59831), .O(n46[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_9 (.CI(n59831), .I0(n13003[6]), .I1(n585), 
            .CO(n59832));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n13003[5]), .I2(n512), 
            .I3(n59830), .O(n46[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n59830), .I0(n13003[5]), .I1(n512), 
            .CO(n59831));
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n13003[4]), .I2(n439), 
            .I3(n59829), .O(n46[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_7 (.CI(n59829), .I0(n13003[4]), .I1(n439), 
            .CO(n59830));
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n78696), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 n78699_bdd_4_lut (.I0(n78699), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4734), .O(n78702));
    defparam n78699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n78690), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n13003[3]), .I2(n366), 
            .I3(n59828), .O(n46[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_6 (.CI(n59828), .I0(n13003[3]), .I1(n366), 
            .CO(n59829));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n13003[2]), .I2(n293_adj_4446), 
            .I3(n59827), .O(n46[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_5 (.CI(n59827), .I0(n13003[2]), .I1(n293_adj_4446), 
            .CO(n59828));
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n13003[1]), .I2(n220), 
            .I3(n59826), .O(n46[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n78684), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY mult_24_add_1225_4 (.CI(n59826), .I0(n13003[1]), .I1(n220), 
            .CO(n59827));
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n13003[0]), .I2(n147), 
            .I3(n59825), .O(n46[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_3 (.CI(n59825), .I0(n13003[0]), .I1(n147), 
            .CO(n59826));
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4442), .I2(n74), 
            .I3(GND_net), .O(n46[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5_adj_4442), .I1(n74), 
            .CO(n59825));
    SB_LUT4 add_6189_23_lut (.I0(GND_net), .I1(n13968[20]), .I2(GND_net), 
            .I3(n59824), .O(n13003[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6189_22_lut (.I0(GND_net), .I1(n13968[19]), .I2(GND_net), 
            .I3(n59823), .O(n13003[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_22 (.CI(n59823), .I0(n13968[19]), .I1(GND_net), 
            .CO(n59824));
    SB_LUT4 add_6189_21_lut (.I0(GND_net), .I1(n13968[18]), .I2(GND_net), 
            .I3(n59822), .O(n13003[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_21 (.CI(n59822), .I0(n13968[18]), .I1(GND_net), 
            .CO(n59823));
    SB_LUT4 add_6189_20_lut (.I0(GND_net), .I1(n13968[17]), .I2(GND_net), 
            .I3(n59821), .O(n13003[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n78678), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_6189_20 (.CI(n59821), .I0(n13968[17]), .I1(GND_net), 
            .CO(n59822));
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n78672), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6189_19_lut (.I0(GND_net), .I1(n13968[16]), .I2(GND_net), 
            .I3(n59820), .O(n13003[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_19 (.CI(n59820), .I0(n13968[16]), .I1(GND_net), 
            .CO(n59821));
    SB_LUT4 add_6189_18_lut (.I0(GND_net), .I1(n13968[15]), .I2(GND_net), 
            .I3(n59819), .O(n13003[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_18 (.CI(n59819), .I0(n13968[15]), .I1(GND_net), 
            .CO(n59820));
    SB_LUT4 add_6189_17_lut (.I0(GND_net), .I1(n13968[14]), .I2(GND_net), 
            .I3(n59818), .O(n13003[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_17 (.CI(n59818), .I0(n13968[14]), .I1(GND_net), 
            .CO(n59819));
    SB_LUT4 add_6189_16_lut (.I0(GND_net), .I1(n13968[13]), .I2(n1099), 
            .I3(n59817), .O(n13003[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_16 (.CI(n59817), .I0(n13968[13]), .I1(n1099), .CO(n59818));
    SB_LUT4 add_6189_15_lut (.I0(GND_net), .I1(n13968[12]), .I2(n1026), 
            .I3(n59816), .O(n13003[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_15 (.CI(n59816), .I0(n13968[12]), .I1(n1026), .CO(n59817));
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n78666), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6189_14_lut (.I0(GND_net), .I1(n13968[11]), .I2(n953), 
            .I3(n59815), .O(n13003[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_14 (.CI(n59815), .I0(n13968[11]), .I1(n953), .CO(n59816));
    SB_LUT4 add_6189_13_lut (.I0(GND_net), .I1(n13968[10]), .I2(n880), 
            .I3(n59814), .O(n13003[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_13 (.CI(n59814), .I0(n13968[10]), .I1(n880), .CO(n59815));
    SB_LUT4 add_6189_12_lut (.I0(GND_net), .I1(n13968[9]), .I2(n807), 
            .I3(n59813), .O(n13003[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_12 (.CI(n59813), .I0(n13968[9]), .I1(n807), .CO(n59814));
    SB_LUT4 add_6189_11_lut (.I0(GND_net), .I1(n13968[8]), .I2(n734), 
            .I3(n59812), .O(n13003[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n78660), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_6189_11 (.CI(n59812), .I0(n13968[8]), .I1(n734), .CO(n59813));
    SB_LUT4 add_6189_10_lut (.I0(GND_net), .I1(n13968[7]), .I2(n661), 
            .I3(n59811), .O(n13003[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_10 (.CI(n59811), .I0(n13968[7]), .I1(n661), .CO(n59812));
    SB_LUT4 add_6189_9_lut (.I0(GND_net), .I1(n13968[6]), .I2(n588), .I3(n59810), 
            .O(n13003[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_9 (.CI(n59810), .I0(n13968[6]), .I1(n588), .CO(n59811));
    SB_LUT4 add_6189_8_lut (.I0(GND_net), .I1(n13968[5]), .I2(n515), .I3(n59809), 
            .O(n13003[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_8 (.CI(n59809), .I0(n13968[5]), .I1(n515), .CO(n59810));
    SB_LUT4 add_6189_7_lut (.I0(GND_net), .I1(n13968[4]), .I2(n442), .I3(n59808), 
            .O(n13003[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_7 (.CI(n59808), .I0(n13968[4]), .I1(n442), .CO(n59809));
    SB_LUT4 add_6189_6_lut (.I0(GND_net), .I1(n13968[3]), .I2(n369), .I3(n59807), 
            .O(n13003[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_6 (.CI(n59807), .I0(n13968[3]), .I1(n369), .CO(n59808));
    SB_LUT4 add_6189_5_lut (.I0(GND_net), .I1(n13968[2]), .I2(n296), .I3(n59806), 
            .O(n13003[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_5 (.CI(n59806), .I0(n13968[2]), .I1(n296), .CO(n59807));
    SB_LUT4 add_6189_4_lut (.I0(GND_net), .I1(n13968[1]), .I2(n223_adj_4439), 
            .I3(n59805), .O(n13003[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_4 (.CI(n59805), .I0(n13968[1]), .I1(n223_adj_4439), 
            .CO(n59806));
    SB_LUT4 add_6189_3_lut (.I0(GND_net), .I1(n13968[0]), .I2(n150), .I3(n59804), 
            .O(n13003[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_3 (.CI(n59804), .I0(n13968[0]), .I1(n150), .CO(n59805));
    SB_LUT4 add_6189_2_lut (.I0(GND_net), .I1(n8_adj_4438), .I2(n77), 
            .I3(GND_net), .O(n13003[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6189_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6189_2 (.CI(GND_net), .I0(n8_adj_4438), .I1(n77), .CO(n59804));
    SB_LUT4 add_6232_22_lut (.I0(GND_net), .I1(n14846[19]), .I2(GND_net), 
            .I3(n59803), .O(n13968[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6232_21_lut (.I0(GND_net), .I1(n14846[18]), .I2(GND_net), 
            .I3(n59802), .O(n13968[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_21 (.CI(n59802), .I0(n14846[18]), .I1(GND_net), 
            .CO(n59803));
    SB_LUT4 add_6232_20_lut (.I0(GND_net), .I1(n14846[17]), .I2(GND_net), 
            .I3(n59801), .O(n13968[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_20 (.CI(n59801), .I0(n14846[17]), .I1(GND_net), 
            .CO(n59802));
    SB_LUT4 add_6232_19_lut (.I0(GND_net), .I1(n14846[16]), .I2(GND_net), 
            .I3(n59800), .O(n13968[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_19 (.CI(n59800), .I0(n14846[16]), .I1(GND_net), 
            .CO(n59801));
    SB_LUT4 add_6232_18_lut (.I0(GND_net), .I1(n14846[15]), .I2(GND_net), 
            .I3(n59799), .O(n13968[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_18 (.CI(n59799), .I0(n14846[15]), .I1(GND_net), 
            .CO(n59800));
    SB_LUT4 add_6232_17_lut (.I0(GND_net), .I1(n14846[14]), .I2(GND_net), 
            .I3(n59798), .O(n13968[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_17 (.CI(n59798), .I0(n14846[14]), .I1(GND_net), 
            .CO(n59799));
    SB_LUT4 add_6232_16_lut (.I0(GND_net), .I1(n14846[13]), .I2(n1102), 
            .I3(n59797), .O(n13968[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_16 (.CI(n59797), .I0(n14846[13]), .I1(n1102), .CO(n59798));
    SB_LUT4 add_6232_15_lut (.I0(GND_net), .I1(n14846[12]), .I2(n1029), 
            .I3(n59796), .O(n13968[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_15 (.CI(n59796), .I0(n14846[12]), .I1(n1029), .CO(n59797));
    SB_LUT4 add_6232_14_lut (.I0(GND_net), .I1(n14846[11]), .I2(n956), 
            .I3(n59795), .O(n13968[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_14 (.CI(n59795), .I0(n14846[11]), .I1(n956), .CO(n59796));
    SB_LUT4 add_6232_13_lut (.I0(GND_net), .I1(n14846[10]), .I2(n883), 
            .I3(n59794), .O(n13968[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_13 (.CI(n59794), .I0(n14846[10]), .I1(n883), .CO(n59795));
    SB_LUT4 add_6232_12_lut (.I0(GND_net), .I1(n14846[9]), .I2(n810), 
            .I3(n59793), .O(n13968[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_12 (.CI(n59793), .I0(n14846[9]), .I1(n810), .CO(n59794));
    SB_LUT4 add_6232_11_lut (.I0(GND_net), .I1(n14846[8]), .I2(n737), 
            .I3(n59792), .O(n13968[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_11 (.CI(n59792), .I0(n14846[8]), .I1(n737), .CO(n59793));
    SB_LUT4 add_6232_10_lut (.I0(GND_net), .I1(n14846[7]), .I2(n664), 
            .I3(n59791), .O(n13968[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_10 (.CI(n59791), .I0(n14846[7]), .I1(n664), .CO(n59792));
    SB_LUT4 add_6232_9_lut (.I0(GND_net), .I1(n14846[6]), .I2(n591), .I3(n59790), 
            .O(n13968[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_9 (.CI(n59790), .I0(n14846[6]), .I1(n591), .CO(n59791));
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n12379[21]), .I2(GND_net), 
            .I3(n58903), .O(n11920[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6232_8_lut (.I0(GND_net), .I1(n14846[5]), .I2(n518), .I3(n59789), 
            .O(n13968[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_8 (.CI(n59789), .I0(n14846[5]), .I1(n518), .CO(n59790));
    SB_LUT4 add_6232_7_lut (.I0(GND_net), .I1(n14846[4]), .I2(n445), .I3(n59788), 
            .O(n13968[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_7 (.CI(n59788), .I0(n14846[4]), .I1(n445), .CO(n59789));
    SB_LUT4 add_6232_6_lut (.I0(GND_net), .I1(n14846[3]), .I2(n372), .I3(n59787), 
            .O(n13968[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_6 (.CI(n59787), .I0(n14846[3]), .I1(n372), .CO(n59788));
    SB_LUT4 add_6232_5_lut (.I0(GND_net), .I1(n14846[2]), .I2(n299_c), 
            .I3(n59786), .O(n13968[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_5 (.CI(n59786), .I0(n14846[2]), .I1(n299_c), .CO(n59787));
    SB_LUT4 add_6232_4_lut (.I0(GND_net), .I1(n14846[1]), .I2(n226), .I3(n59785), 
            .O(n13968[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_4 (.CI(n59785), .I0(n14846[1]), .I1(n226), .CO(n59786));
    SB_LUT4 add_6232_3_lut (.I0(GND_net), .I1(n14846[0]), .I2(n153), .I3(n59784), 
            .O(n13968[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n12379[20]), .I2(GND_net), 
            .I3(n58902), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n58902), .I0(n12379[20]), .I1(GND_net), 
            .CO(n58903));
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n12379[19]), .I2(GND_net), 
            .I3(n58901), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_22 (.CI(n58901), .I0(n12379[19]), .I1(GND_net), 
            .CO(n58902));
    SB_CARRY add_6232_3 (.CI(n59784), .I0(n14846[0]), .I1(n153), .CO(n59785));
    SB_LUT4 add_6232_2_lut (.I0(GND_net), .I1(n11), .I2(n80), .I3(GND_net), 
            .O(n13968[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6232_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6232_2 (.CI(GND_net), .I0(n11), .I1(n80), .CO(n59784));
    SB_LUT4 add_6529_12_lut (.I0(GND_net), .I1(n19635[9]), .I2(n840), 
            .I3(n59783), .O(n19372[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6529_11_lut (.I0(GND_net), .I1(n19635[8]), .I2(n767), 
            .I3(n59782), .O(n19372[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_11 (.CI(n59782), .I0(n19635[8]), .I1(n767), .CO(n59783));
    SB_LUT4 add_6529_10_lut (.I0(GND_net), .I1(n19635[7]), .I2(n694), 
            .I3(n59781), .O(n19372[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_10 (.CI(n59781), .I0(n19635[7]), .I1(n694), .CO(n59782));
    SB_LUT4 add_6529_9_lut (.I0(GND_net), .I1(n19635[6]), .I2(n621), .I3(n59780), 
            .O(n19372[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_9 (.CI(n59780), .I0(n19635[6]), .I1(n621), .CO(n59781));
    SB_LUT4 add_6529_8_lut (.I0(GND_net), .I1(n19635[5]), .I2(n548), .I3(n59779), 
            .O(n19372[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_8 (.CI(n59779), .I0(n19635[5]), .I1(n548), .CO(n59780));
    SB_LUT4 add_6529_7_lut (.I0(GND_net), .I1(n19635[4]), .I2(n475_c), 
            .I3(n59778), .O(n19372[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_7 (.CI(n59778), .I0(n19635[4]), .I1(n475_c), .CO(n59779));
    SB_LUT4 add_6529_6_lut (.I0(GND_net), .I1(n19635[3]), .I2(n402), .I3(n59777), 
            .O(n19372[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_6 (.CI(n59777), .I0(n19635[3]), .I1(n402), .CO(n59778));
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n12379[18]), .I2(GND_net), 
            .I3(n58900), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6529_5_lut (.I0(GND_net), .I1(n19635[2]), .I2(n329), .I3(n59776), 
            .O(n19372[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n58900), .I0(n12379[18]), .I1(GND_net), 
            .CO(n58901));
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n12379[17]), .I2(GND_net), 
            .I3(n58899), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_20 (.CI(n58899), .I0(n12379[17]), .I1(GND_net), 
            .CO(n58900));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n12379[16]), .I2(GND_net), 
            .I3(n58898), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n58898), .I0(n12379[16]), .I1(GND_net), 
            .CO(n58899));
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6529_5 (.CI(n59776), .I0(n19635[2]), .I1(n329), .CO(n59777));
    SB_LUT4 add_6529_4_lut (.I0(GND_net), .I1(n19635[1]), .I2(n256), .I3(n59775), 
            .O(n19372[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_4 (.CI(n59775), .I0(n19635[1]), .I1(n256), .CO(n59776));
    SB_LUT4 add_6529_3_lut (.I0(GND_net), .I1(n19635[0]), .I2(n183), .I3(n59774), 
            .O(n19372[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_3 (.CI(n59774), .I0(n19635[0]), .I1(n183), .CO(n59775));
    SB_LUT4 add_6529_2_lut (.I0(GND_net), .I1(n41_c), .I2(n110_c), .I3(GND_net), 
            .O(n19372[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6529_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6529_2 (.CI(GND_net), .I0(n41_c), .I1(n110_c), .CO(n59774));
    SB_LUT4 add_6272_21_lut (.I0(GND_net), .I1(n15642[18]), .I2(GND_net), 
            .I3(n59773), .O(n14846[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n12379[15]), .I2(GND_net), 
            .I3(n58897), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_18 (.CI(n58897), .I0(n12379[15]), .I1(GND_net), 
            .CO(n58898));
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n12379[14]), .I2(GND_net), 
            .I3(n58896), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_17 (.CI(n58896), .I0(n12379[14]), .I1(GND_net), 
            .CO(n58897));
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n12379[13]), .I2(n1096_adj_4475), 
            .I3(n58895), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6272_20_lut (.I0(GND_net), .I1(n15642[17]), .I2(GND_net), 
            .I3(n59772), .O(n14846[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_20 (.CI(n59772), .I0(n15642[17]), .I1(GND_net), 
            .CO(n59773));
    SB_LUT4 add_6272_19_lut (.I0(GND_net), .I1(n15642[16]), .I2(GND_net), 
            .I3(n59771), .O(n14846[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_19 (.CI(n59771), .I0(n15642[16]), .I1(GND_net), 
            .CO(n59772));
    SB_LUT4 add_6272_18_lut (.I0(GND_net), .I1(n15642[15]), .I2(GND_net), 
            .I3(n59770), .O(n14846[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_18 (.CI(n59770), .I0(n15642[15]), .I1(GND_net), 
            .CO(n59771));
    SB_LUT4 add_6272_17_lut (.I0(GND_net), .I1(n15642[14]), .I2(GND_net), 
            .I3(n59769), .O(n14846[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n58895), .I0(n12379[13]), .I1(n1096_adj_4475), 
            .CO(n58896));
    SB_CARRY add_6272_17 (.CI(n59769), .I0(n15642[14]), .I1(GND_net), 
            .CO(n59770));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n12379[12]), .I2(n1023_adj_4466), 
            .I3(n58894), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6272_16_lut (.I0(GND_net), .I1(n15642[13]), .I2(n1105), 
            .I3(n59768), .O(n14846[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4476));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_16 (.CI(n59768), .I0(n15642[13]), .I1(n1105), .CO(n59769));
    SB_LUT4 add_6272_15_lut (.I0(GND_net), .I1(n15642[12]), .I2(n1032), 
            .I3(n59767), .O(n14846[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4477));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4478));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4479));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_15 (.CI(n59767), .I0(n15642[12]), .I1(n1032), .CO(n59768));
    SB_LUT4 add_6272_14_lut (.I0(GND_net), .I1(n15642[11]), .I2(n959), 
            .I3(n59766), .O(n14846[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4480));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_14 (.CI(n59766), .I0(n15642[11]), .I1(n959), .CO(n59767));
    SB_LUT4 add_6272_13_lut (.I0(GND_net), .I1(n15642[10]), .I2(n886), 
            .I3(n59765), .O(n14846[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_13 (.CI(n59765), .I0(n15642[10]), .I1(n886), .CO(n59766));
    SB_LUT4 add_6272_12_lut (.I0(GND_net), .I1(n15642[9]), .I2(n813), 
            .I3(n59764), .O(n14846[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_12 (.CI(n59764), .I0(n15642[9]), .I1(n813), .CO(n59765));
    SB_CARRY mult_23_add_1221_15 (.CI(n58894), .I0(n12379[12]), .I1(n1023_adj_4466), 
            .CO(n58895));
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n12379[11]), .I2(n950_adj_4465), 
            .I3(n58893), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6272_11_lut (.I0(GND_net), .I1(n15642[8]), .I2(n740), 
            .I3(n59763), .O(n14846[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_11 (.CI(n59763), .I0(n15642[8]), .I1(n740), .CO(n59764));
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4482));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_10_lut (.I0(GND_net), .I1(n15642[7]), .I2(n667), 
            .I3(n59762), .O(n14846[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_10 (.CI(n59762), .I0(n15642[7]), .I1(n667), .CO(n59763));
    SB_LUT4 add_6272_9_lut (.I0(GND_net), .I1(n15642[6]), .I2(n594), .I3(n59761), 
            .O(n14846[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4483));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4484));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_9 (.CI(n59761), .I0(n15642[6]), .I1(n594), .CO(n59762));
    SB_LUT4 add_6272_8_lut (.I0(GND_net), .I1(n15642[5]), .I2(n521), .I3(n59760), 
            .O(n14846[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4485));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_8 (.CI(n59760), .I0(n15642[5]), .I1(n521), .CO(n59761));
    SB_CARRY mult_23_add_1221_14 (.CI(n58893), .I0(n12379[11]), .I1(n950_adj_4465), 
            .CO(n58894));
    SB_LUT4 add_6272_7_lut (.I0(GND_net), .I1(n15642[4]), .I2(n448), .I3(n59759), 
            .O(n14846[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4486));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n12379[10]), .I2(n877_adj_4464), 
            .I3(n58892), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_13 (.CI(n58892), .I0(n12379[10]), .I1(n877_adj_4464), 
            .CO(n58893));
    SB_LUT4 i1_4_lut_adj_949 (.I0(n20462[2]), .I1(n6), .I2(n37336), .I3(\Ki[4] ), 
            .O(n20416[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h9666;
    SB_CARRY add_6272_7 (.CI(n59759), .I0(n15642[4]), .I1(n448), .CO(n59760));
    SB_LUT4 add_6272_6_lut (.I0(GND_net), .I1(n15642[3]), .I2(n375), .I3(n59758), 
            .O(n14846[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_6 (.CI(n59758), .I0(n15642[3]), .I1(n375), .CO(n59759));
    SB_LUT4 mult_24_i138_2_lut (.I0(\Ki[2] ), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_5_lut (.I0(GND_net), .I1(n15642[2]), .I2(n302_adj_4488), 
            .I3(n59757), .O(n14846[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_5 (.CI(n59757), .I0(n15642[2]), .I1(n302_adj_4488), 
            .CO(n59758));
    SB_LUT4 i1_4_lut_adj_950 (.I0(n20499[0]), .I1(n58049), .I2(\Ki[2] ), 
            .I3(n339), .O(n20490[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h9666;
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n12379[9]), .I2(n804_adj_4490), 
            .I3(n58891), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i89_2_lut (.I0(\Ki[1] ), .I1(n340), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i42_2_lut (.I0(\Ki[0] ), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4491));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_4_lut (.I0(GND_net), .I1(n15642[1]), .I2(n229), .I3(n59756), 
            .O(n14846[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_4 (.CI(n59756), .I0(n15642[1]), .I1(n229), .CO(n59757));
    SB_LUT4 add_6272_3_lut (.I0(GND_net), .I1(n15642[0]), .I2(n156), .I3(n59755), 
            .O(n14846[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_3 (.CI(n59755), .I0(n15642[0]), .I1(n156), .CO(n59756));
    SB_LUT4 add_6272_2_lut (.I0(GND_net), .I1(n14_adj_4492), .I2(n83), 
            .I3(GND_net), .O(n14846[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_2 (.CI(GND_net), .I0(n14_adj_4492), .I1(n83), .CO(n59755));
    SB_LUT4 add_6310_20_lut (.I0(GND_net), .I1(n16360[17]), .I2(GND_net), 
            .I3(n59754), .O(n15642[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6310_19_lut (.I0(GND_net), .I1(n16360[16]), .I2(GND_net), 
            .I3(n59753), .O(n15642[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_19 (.CI(n59753), .I0(n16360[16]), .I1(GND_net), 
            .CO(n59754));
    SB_LUT4 add_6310_18_lut (.I0(GND_net), .I1(n16360[15]), .I2(GND_net), 
            .I3(n59752), .O(n15642[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_18 (.CI(n59752), .I0(n16360[15]), .I1(GND_net), 
            .CO(n59753));
    SB_CARRY mult_23_add_1221_12 (.CI(n58891), .I0(n12379[9]), .I1(n804_adj_4490), 
            .CO(n58892));
    SB_LUT4 add_6310_17_lut (.I0(GND_net), .I1(n16360[14]), .I2(GND_net), 
            .I3(n59751), .O(n15642[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_17 (.CI(n59751), .I0(n16360[14]), .I1(GND_net), 
            .CO(n59752));
    SB_LUT4 add_6310_16_lut (.I0(GND_net), .I1(n16360[13]), .I2(n1108_adj_4493), 
            .I3(n59750), .O(n15642[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_16 (.CI(n59750), .I0(n16360[13]), .I1(n1108_adj_4493), 
            .CO(n59751));
    SB_LUT4 add_6310_15_lut (.I0(GND_net), .I1(n16360[12]), .I2(n1035_adj_4494), 
            .I3(n59749), .O(n15642[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_15 (.CI(n59749), .I0(n16360[12]), .I1(n1035_adj_4494), 
            .CO(n59750));
    SB_LUT4 add_6310_14_lut (.I0(GND_net), .I1(n16360[11]), .I2(n962_adj_4495), 
            .I3(n59748), .O(n15642[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4496));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6310_14 (.CI(n59748), .I0(n16360[11]), .I1(n962_adj_4495), 
            .CO(n59749));
    SB_LUT4 add_6310_13_lut (.I0(GND_net), .I1(n16360[10]), .I2(n889_adj_4497), 
            .I3(n59747), .O(n15642[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_951 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n337), .I3(n336), 
            .O(n70829));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h93a0;
    SB_CARRY add_6310_13 (.CI(n59747), .I0(n16360[10]), .I1(n889_adj_4497), 
            .CO(n59748));
    SB_LUT4 i1_4_lut_adj_952 (.I0(n37336), .I1(\Ki[4] ), .I2(\Ki[5] ), 
            .I3(n340), .O(n70833));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_6310_12_lut (.I0(GND_net), .I1(n16360[9]), .I2(n816_adj_4498), 
            .I3(n59746), .O(n15642[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n12379[8]), .I2(n731_adj_4499), 
            .I3(n58890), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_11 (.CI(n58890), .I0(n12379[8]), .I1(n731_adj_4499), 
            .CO(n58891));
    SB_CARRY add_6310_12 (.CI(n59746), .I0(n16360[9]), .I1(n816_adj_4498), 
            .CO(n59747));
    SB_LUT4 add_6310_11_lut (.I0(GND_net), .I1(n16360[8]), .I2(n743_adj_4500), 
            .I3(n59745), .O(n15642[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_953 (.I0(\Ki[3] ), .I1(n37146), .I2(n339), .I3(\Ki[2] ), 
            .O(n70831));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h6ca0;
    SB_CARRY add_6310_11 (.CI(n59745), .I0(n16360[8]), .I1(n743_adj_4500), 
            .CO(n59746));
    SB_LUT4 add_6310_10_lut (.I0(GND_net), .I1(n16360[7]), .I2(n670_adj_4501), 
            .I3(n59744), .O(n15642[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_954 (.I0(n70831), .I1(n57998), .I2(n70833), .I3(n70829), 
            .O(n70839));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_CARRY add_6310_10 (.CI(n59744), .I0(n16360[7]), .I1(n670_adj_4501), 
            .CO(n59745));
    SB_LUT4 i44005_4_lut (.I0(n20499[0]), .I1(\Ki[2] ), .I2(n58049), .I3(n339), 
            .O(n4_adj_4502));   // verilog/motorControl.v(61[29:40])
    defparam i44005_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_6310_9_lut (.I0(GND_net), .I1(n16360[6]), .I2(n597_adj_4503), 
            .I3(n59743), .O(n15642[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i43837_4_lut (.I0(n20462[2]), .I1(n37336), .I2(n6), .I3(\Ki[4] ), 
            .O(n8_adj_4504));   // verilog/motorControl.v(61[29:40])
    defparam i43837_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY add_6310_9 (.CI(n59743), .I0(n16360[6]), .I1(n597_adj_4503), 
            .CO(n59744));
    SB_LUT4 add_6310_8_lut (.I0(GND_net), .I1(n16360[5]), .I2(n524_adj_4505), 
            .I3(n59742), .O(n15642[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_8 (.CI(n59742), .I0(n16360[5]), .I1(n524_adj_4505), 
            .CO(n59743));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n12379[7]), .I2(n658_adj_4506), 
            .I3(n58889), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_10 (.CI(n58889), .I0(n12379[7]), .I1(n658_adj_4506), 
            .CO(n58890));
    SB_LUT4 i1_4_lut_adj_955 (.I0(n6_adj_4507), .I1(n8_adj_4504), .I2(n4_adj_4502), 
            .I3(n70839), .O(n69074));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 add_6310_7_lut (.I0(GND_net), .I1(n16360[4]), .I2(n451_adj_4508), 
            .I3(n59741), .O(n15642[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_7 (.CI(n59741), .I0(n16360[4]), .I1(n451_adj_4508), 
            .CO(n59742));
    SB_LUT4 add_6310_6_lut (.I0(GND_net), .I1(n16360[3]), .I2(n378_adj_4509), 
            .I3(n59740), .O(n15642[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_6 (.CI(n59740), .I0(n16360[3]), .I1(n378_adj_4509), 
            .CO(n59741));
    SB_LUT4 add_6310_5_lut (.I0(GND_net), .I1(n16360[2]), .I2(n305_adj_4510), 
            .I3(n59739), .O(n15642[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n12379[6]), .I2(n585_adj_4512), 
            .I3(n58888), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_5 (.CI(n59739), .I0(n16360[2]), .I1(n305_adj_4510), 
            .CO(n59740));
    SB_CARRY mult_23_add_1221_9 (.CI(n58888), .I0(n12379[6]), .I1(n585_adj_4512), 
            .CO(n58889));
    SB_LUT4 add_6310_4_lut (.I0(GND_net), .I1(n16360[1]), .I2(n232_adj_4513), 
            .I3(n59738), .O(n15642[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_4 (.CI(n59738), .I0(n16360[1]), .I1(n232_adj_4513), 
            .CO(n59739));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n12379[5]), .I2(n512_adj_4514), 
            .I3(n58887), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_8 (.CI(n58887), .I0(n12379[5]), .I1(n512_adj_4514), 
            .CO(n58888));
    SB_LUT4 add_6310_3_lut (.I0(GND_net), .I1(n16360[0]), .I2(n159_adj_4515), 
            .I3(n59737), .O(n15642[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6310_3 (.CI(n59737), .I0(n16360[0]), .I1(n159_adj_4515), 
            .CO(n59738));
    SB_LUT4 add_6310_2_lut (.I0(GND_net), .I1(n17_adj_4516), .I2(n86_adj_4517), 
            .I3(GND_net), .O(n15642[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6310_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6310_2 (.CI(GND_net), .I0(n17_adj_4516), .I1(n86_adj_4517), 
            .CO(n59737));
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n12379[4]), .I2(n439_adj_4519), 
            .I3(n58886), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_7 (.CI(n58886), .I0(n12379[4]), .I1(n439_adj_4519), 
            .CO(n58887));
    SB_LUT4 add_6550_11_lut (.I0(GND_net), .I1(n19854[8]), .I2(n770), 
            .I3(n59736), .O(n19635[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_10_lut (.I0(GND_net), .I1(n19854[7]), .I2(n697), 
            .I3(n59735), .O(n19635[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_10 (.CI(n59735), .I0(n19854[7]), .I1(n697), .CO(n59736));
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n12379[3]), .I2(n366_adj_4521), 
            .I3(n58885), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n58885), .I0(n12379[3]), .I1(n366_adj_4521), 
            .CO(n58886));
    SB_LUT4 add_6550_9_lut (.I0(GND_net), .I1(n19854[6]), .I2(n624), .I3(n59734), 
            .O(n19635[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4522));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4523));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6550_9 (.CI(n59734), .I0(n19854[6]), .I1(n624), .CO(n59735));
    SB_LUT4 add_6550_8_lut (.I0(GND_net), .I1(n19854[5]), .I2(n551), .I3(n59733), 
            .O(n19635[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_8 (.CI(n59733), .I0(n19854[5]), .I1(n551), .CO(n59734));
    SB_LUT4 add_6550_7_lut (.I0(GND_net), .I1(n19854[4]), .I2(n478), .I3(n59732), 
            .O(n19635[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_7 (.CI(n59732), .I0(n19854[4]), .I1(n478), .CO(n59733));
    SB_CARRY add_16_10 (.CI(n58198), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n58199));
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n12379[2]), .I2(n293_adj_4524), 
            .I3(n58884), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4525));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_5 (.CI(n58884), .I0(n12379[2]), .I1(n293_adj_4524), 
            .CO(n58885));
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n58197), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_6_lut (.I0(GND_net), .I1(n19854[3]), .I2(n405), .I3(n59731), 
            .O(n19635[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_6 (.CI(n59731), .I0(n19854[3]), .I1(n405), .CO(n59732));
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4527));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n12379[1]), .I2(n220_adj_4528), 
            .I3(n58883), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4529));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4530));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4531));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6550_5_lut (.I0(GND_net), .I1(n19854[2]), .I2(n332_adj_4532), 
            .I3(n59730), .O(n19635[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4533));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6550_5 (.CI(n59730), .I0(n19854[2]), .I1(n332_adj_4532), 
            .CO(n59731));
    SB_LUT4 add_6550_4_lut (.I0(GND_net), .I1(n19854[1]), .I2(n259), .I3(n59729), 
            .O(n19635[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_4 (.CI(n58883), .I0(n12379[1]), .I1(n220_adj_4528), 
            .CO(n58884));
    SB_CARRY add_6550_4 (.CI(n59729), .I0(n19854[1]), .I1(n259), .CO(n59730));
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4534));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6550_3_lut (.I0(GND_net), .I1(n19854[0]), .I2(n186), .I3(n59728), 
            .O(n19635[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4535));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6550_3 (.CI(n59728), .I0(n19854[0]), .I1(n186), .CO(n59729));
    SB_LUT4 add_6550_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19635[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n12379[0]), .I2(n147_adj_4537), 
            .I3(n58882), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4538));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6550_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n59728));
    SB_LUT4 add_6346_19_lut (.I0(GND_net), .I1(n17004[16]), .I2(GND_net), 
            .I3(n59727), .O(n16360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6346_18_lut (.I0(GND_net), .I1(n17004[15]), .I2(GND_net), 
            .I3(n59726), .O(n16360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11880_bdd_4_lut_62825 (.I0(n11880), .I1(n74600), .I2(setpoint[8]), 
            .I3(n4734), .O(n78693));
    defparam n11880_bdd_4_lut_62825.LUT_INIT = 16'he4aa;
    SB_CARRY add_6346_18 (.CI(n59726), .I0(n17004[15]), .I1(GND_net), 
            .CO(n59727));
    SB_LUT4 add_6346_17_lut (.I0(GND_net), .I1(n17004[14]), .I2(GND_net), 
            .I3(n59725), .O(n16360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_17 (.CI(n59725), .I0(n17004[14]), .I1(GND_net), 
            .CO(n59726));
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4540));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6346_16_lut (.I0(GND_net), .I1(n17004[13]), .I2(n1111_adj_4541), 
            .I3(n59724), .O(n16360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_16 (.CI(n59724), .I0(n17004[13]), .I1(n1111_adj_4541), 
            .CO(n59725));
    SB_LUT4 add_6346_15_lut (.I0(GND_net), .I1(n17004[12]), .I2(n1038_adj_4542), 
            .I3(n59723), .O(n16360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_15 (.CI(n59723), .I0(n17004[12]), .I1(n1038_adj_4542), 
            .CO(n59724));
    SB_LUT4 add_6346_14_lut (.I0(GND_net), .I1(n17004[11]), .I2(n965_adj_4543), 
            .I3(n59722), .O(n16360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_14 (.CI(n59722), .I0(n17004[11]), .I1(n965_adj_4543), 
            .CO(n59723));
    SB_LUT4 add_6346_13_lut (.I0(GND_net), .I1(n17004[10]), .I2(n892_adj_4544), 
            .I3(n59721), .O(n16360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_13 (.CI(n59721), .I0(n17004[10]), .I1(n892_adj_4544), 
            .CO(n59722));
    SB_LUT4 add_6346_12_lut (.I0(GND_net), .I1(n17004[9]), .I2(n819_adj_4545), 
            .I3(n59720), .O(n16360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4546));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78693_bdd_4_lut (.I0(n78693), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4734), .O(n78696));
    defparam n78693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4548));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4549));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_12 (.CI(n59720), .I0(n17004[9]), .I1(n819_adj_4545), 
            .CO(n59721));
    SB_LUT4 add_6346_11_lut (.I0(GND_net), .I1(n17004[8]), .I2(n746_adj_4550), 
            .I3(n59719), .O(n16360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_11 (.CI(n59719), .I0(n17004[8]), .I1(n746_adj_4550), 
            .CO(n59720));
    SB_LUT4 add_6346_10_lut (.I0(GND_net), .I1(n17004[7]), .I2(n673_adj_4551), 
            .I3(n59718), .O(n16360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_10 (.CI(n59718), .I0(n17004[7]), .I1(n673_adj_4551), 
            .CO(n59719));
    SB_LUT4 add_6346_9_lut (.I0(GND_net), .I1(n17004[6]), .I2(n600_adj_4552), 
            .I3(n59717), .O(n16360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_9 (.CI(n59717), .I0(n17004[6]), .I1(n600_adj_4552), 
            .CO(n59718));
    SB_LUT4 add_6346_8_lut (.I0(GND_net), .I1(n17004[5]), .I2(n527_adj_4553), 
            .I3(n59716), .O(n16360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_8 (.CI(n59716), .I0(n17004[5]), .I1(n527_adj_4553), 
            .CO(n59717));
    SB_LUT4 add_6346_7_lut (.I0(GND_net), .I1(n17004[4]), .I2(n454_adj_4555), 
            .I3(n59715), .O(n16360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_7 (.CI(n59715), .I0(n17004[4]), .I1(n454_adj_4555), 
            .CO(n59716));
    SB_LUT4 add_6346_6_lut (.I0(GND_net), .I1(n17004[3]), .I2(n381), .I3(n59714), 
            .O(n16360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62820 (.I0(n11880), .I1(n74599), .I2(setpoint[7]), 
            .I3(n4734), .O(n78687));
    defparam n11880_bdd_4_lut_62820.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_6 (.CI(n59714), .I0(n17004[3]), .I1(n381), .CO(n59715));
    SB_LUT4 add_6346_5_lut (.I0(GND_net), .I1(n17004[2]), .I2(n308_adj_4557), 
            .I3(n59713), .O(n16360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n78687_bdd_4_lut (.I0(n78687), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4734), .O(n78690));
    defparam n78687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_6346_5 (.CI(n59713), .I0(n17004[2]), .I1(n308_adj_4557), 
            .CO(n59714));
    SB_LUT4 add_6346_4_lut (.I0(GND_net), .I1(n17004[1]), .I2(n235_adj_4559), 
            .I3(n59712), .O(n16360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6346_4 (.CI(n59712), .I0(n17004[1]), .I1(n235_adj_4559), 
            .CO(n59713));
    SB_LUT4 add_6346_3_lut (.I0(GND_net), .I1(n17004[0]), .I2(n162), .I3(n59711), 
            .O(n16360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11880_bdd_4_lut_62815 (.I0(n11880), .I1(n74598), .I2(setpoint[6]), 
            .I3(n4734), .O(n78681));
    defparam n11880_bdd_4_lut_62815.LUT_INIT = 16'he4aa;
    SB_LUT4 n78681_bdd_4_lut (.I0(n78681), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4734), .O(n78684));
    defparam n78681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6346_3 (.CI(n59711), .I0(n17004[0]), .I1(n162), .CO(n59712));
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6346_2_lut (.I0(GND_net), .I1(n20_adj_4561), .I2(n89), 
            .I3(GND_net), .O(n16360[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6346_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6346_2 (.CI(GND_net), .I0(n20_adj_4561), .I1(n89), .CO(n59711));
    SB_LUT4 add_6380_18_lut (.I0(GND_net), .I1(n17578[15]), .I2(GND_net), 
            .I3(n59710), .O(n17004[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6380_17_lut (.I0(GND_net), .I1(n17578[14]), .I2(GND_net), 
            .I3(n59709), .O(n17004[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_17 (.CI(n59709), .I0(n17578[14]), .I1(GND_net), 
            .CO(n59710));
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6380_16_lut (.I0(GND_net), .I1(n17578[13]), .I2(n1114), 
            .I3(n59708), .O(n17004[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_16 (.CI(n59708), .I0(n17578[13]), .I1(n1114), .CO(n59709));
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4475));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_3 (.CI(n58882), .I0(n12379[0]), .I1(n147_adj_4537), 
            .CO(n58883));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_4563), .I2(n74_adj_4564), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6380_15_lut (.I0(GND_net), .I1(n17578[12]), .I2(n1041), 
            .I3(n59707), .O(n17004[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_15 (.CI(n59707), .I0(n17578[12]), .I1(n1041), .CO(n59708));
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6380_14_lut (.I0(GND_net), .I1(n17578[11]), .I2(n968), 
            .I3(n59706), .O(n17004[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_14 (.CI(n59706), .I0(n17578[11]), .I1(n968), .CO(n59707));
    SB_LUT4 add_6380_13_lut (.I0(GND_net), .I1(n17578[10]), .I2(n895), 
            .I3(n59705), .O(n17004[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6380_13 (.CI(n59705), .I0(n17578[10]), .I1(n895), .CO(n59706));
    SB_LUT4 add_6380_12_lut (.I0(GND_net), .I1(n17578[9]), .I2(n822), 
            .I3(n59704), .O(n17004[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6380_12 (.CI(n59704), .I0(n17578[9]), .I1(n822), .CO(n59705));
    SB_LUT4 add_6380_11_lut (.I0(GND_net), .I1(n17578[8]), .I2(n749), 
            .I3(n59703), .O(n17004[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6380_11 (.CI(n59703), .I0(n17578[8]), .I1(n749), .CO(n59704));
    SB_LUT4 add_6380_10_lut (.I0(GND_net), .I1(n17578[7]), .I2(n676), 
            .I3(n59702), .O(n17004[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11880_bdd_4_lut_62810 (.I0(n11880), .I1(n74597), .I2(setpoint[5]), 
            .I3(n4734), .O(n78675));
    defparam n11880_bdd_4_lut_62810.LUT_INIT = 16'he4aa;
    SB_CARRY add_6380_10 (.CI(n59702), .I0(n17578[7]), .I1(n676), .CO(n59703));
    SB_LUT4 add_6380_9_lut (.I0(GND_net), .I1(n17578[6]), .I2(n603), .I3(n59701), 
            .O(n17004[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_9 (.CI(n59701), .I0(n17578[6]), .I1(n603), .CO(n59702));
    SB_LUT4 add_6380_8_lut (.I0(GND_net), .I1(n17578[5]), .I2(n530), .I3(n59700), 
            .O(n17004[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_8 (.CI(n59700), .I0(n17578[5]), .I1(n530), .CO(n59701));
    SB_LUT4 add_6380_7_lut (.I0(GND_net), .I1(n17578[4]), .I2(n457), .I3(n59699), 
            .O(n17004[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_7 (.CI(n59699), .I0(n17578[4]), .I1(n457), .CO(n59700));
    SB_LUT4 add_6380_6_lut (.I0(GND_net), .I1(n17578[3]), .I2(n384_adj_4568), 
            .I3(n59698), .O(n17004[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_6 (.CI(n59698), .I0(n17578[3]), .I1(n384_adj_4568), 
            .CO(n59699));
    SB_LUT4 add_6380_5_lut (.I0(GND_net), .I1(n17578[2]), .I2(n311_adj_4569), 
            .I3(n59697), .O(n17004[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_5 (.CI(n59697), .I0(n17578[2]), .I1(n311_adj_4569), 
            .CO(n59698));
    SB_LUT4 add_6380_4_lut (.I0(GND_net), .I1(n17578[1]), .I2(n238_adj_4570), 
            .I3(n59696), .O(n17004[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_4 (.CI(n59696), .I0(n17578[1]), .I1(n238_adj_4570), 
            .CO(n59697));
    SB_LUT4 add_6380_3_lut (.I0(GND_net), .I1(n17578[0]), .I2(n165), .I3(n59695), 
            .O(n17004[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6380_3 (.CI(n59695), .I0(n17578[0]), .I1(n165), .CO(n59696));
    SB_LUT4 add_6380_2_lut (.I0(GND_net), .I1(n23_adj_4574), .I2(n92), 
            .I3(GND_net), .O(n17004[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6380_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5_adj_4563), .I1(n74_adj_4564), 
            .CO(n58882));
    SB_LUT4 add_6562_11_lut (.I0(GND_net), .I1(n19972[8]), .I2(n770_adj_4575), 
            .I3(n58881), .O(n19776[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6380_2 (.CI(GND_net), .I0(n23_adj_4574), .I1(n92), .CO(n59695));
    SB_LUT4 add_6569_10_lut (.I0(GND_net), .I1(n20033[7]), .I2(n700_adj_4576), 
            .I3(n59694), .O(n19854[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_10_lut (.I0(GND_net), .I1(n19972[7]), .I2(n697_adj_4577), 
            .I3(n58880), .O(n19776[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6569_9_lut (.I0(GND_net), .I1(n20033[6]), .I2(n627_adj_4578), 
            .I3(n59693), .O(n19854[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_9 (.CI(n59693), .I0(n20033[6]), .I1(n627_adj_4578), 
            .CO(n59694));
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6569_8_lut (.I0(GND_net), .I1(n20033[5]), .I2(n554_adj_4579), 
            .I3(n59692), .O(n19854[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_8 (.CI(n59692), .I0(n20033[5]), .I1(n554_adj_4579), 
            .CO(n59693));
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6569_7_lut (.I0(GND_net), .I1(n20033[4]), .I2(n481_adj_4580), 
            .I3(n59691), .O(n19854[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6569_7 (.CI(n59691), .I0(n20033[4]), .I1(n481_adj_4580), 
            .CO(n59692));
    SB_LUT4 add_6569_6_lut (.I0(GND_net), .I1(n20033[3]), .I2(n408_adj_4582), 
            .I3(n59690), .O(n19854[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_6 (.CI(n59690), .I0(n20033[3]), .I1(n408_adj_4582), 
            .CO(n59691));
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4583));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6569_5_lut (.I0(GND_net), .I1(n20033[2]), .I2(n335_adj_4584), 
            .I3(n59689), .O(n19854[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_5 (.CI(n59689), .I0(n20033[2]), .I1(n335_adj_4584), 
            .CO(n59690));
    SB_LUT4 add_6569_4_lut (.I0(GND_net), .I1(n20033[1]), .I2(n262_adj_4585), 
            .I3(n59688), .O(n19854[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_4 (.CI(n59688), .I0(n20033[1]), .I1(n262_adj_4585), 
            .CO(n59689));
    SB_LUT4 add_6569_3_lut (.I0(GND_net), .I1(n20033[0]), .I2(n189_adj_4586), 
            .I3(n59687), .O(n19854[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_3 (.CI(n59687), .I0(n20033[0]), .I1(n189_adj_4586), 
            .CO(n59688));
    SB_LUT4 add_6569_2_lut (.I0(GND_net), .I1(n47_adj_4587), .I2(n116_adj_4588), 
            .I3(GND_net), .O(n19854[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6569_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6569_2 (.CI(GND_net), .I0(n47_adj_4587), .I1(n116_adj_4588), 
            .CO(n59687));
    SB_LUT4 add_6412_17_lut (.I0(GND_net), .I1(n18086[14]), .I2(GND_net), 
            .I3(n59686), .O(n17578[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6412_16_lut (.I0(GND_net), .I1(n18086[13]), .I2(n1117), 
            .I3(n59685), .O(n17578[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n78675_bdd_4_lut (.I0(n78675), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4734), .O(n78678));
    defparam n78675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_6412_16 (.CI(n59685), .I0(n18086[13]), .I1(n1117), .CO(n59686));
    SB_LUT4 add_6412_15_lut (.I0(GND_net), .I1(n18086[12]), .I2(n1044), 
            .I3(n59684), .O(n17578[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_15 (.CI(n59684), .I0(n18086[12]), .I1(n1044), .CO(n59685));
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4590));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6412_14_lut (.I0(GND_net), .I1(n18086[11]), .I2(n971), 
            .I3(n59683), .O(n17578[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_14 (.CI(n59683), .I0(n18086[11]), .I1(n971), .CO(n59684));
    SB_LUT4 add_6412_13_lut (.I0(GND_net), .I1(n18086[10]), .I2(n898), 
            .I3(n59682), .O(n17578[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_13 (.CI(n59682), .I0(n18086[10]), .I1(n898), .CO(n59683));
    SB_LUT4 add_6412_12_lut (.I0(GND_net), .I1(n18086[9]), .I2(n825), 
            .I3(n59681), .O(n17578[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_12 (.CI(n59681), .I0(n18086[9]), .I1(n825), .CO(n59682));
    SB_LUT4 add_6412_11_lut (.I0(GND_net), .I1(n18086[8]), .I2(n752), 
            .I3(n59680), .O(n17578[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_10 (.CI(n58880), .I0(n19972[7]), .I1(n697_adj_4577), 
            .CO(n58881));
    SB_CARRY add_6412_11 (.CI(n59680), .I0(n18086[8]), .I1(n752), .CO(n59681));
    SB_LUT4 add_6412_10_lut (.I0(GND_net), .I1(n18086[7]), .I2(n679), 
            .I3(n59679), .O(n17578[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_10 (.CI(n59679), .I0(n18086[7]), .I1(n679), .CO(n59680));
    SB_LUT4 add_6412_9_lut (.I0(GND_net), .I1(n18086[6]), .I2(n606), .I3(n59678), 
            .O(n17578[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_9 (.CI(n59678), .I0(n18086[6]), .I1(n606), .CO(n59679));
    SB_LUT4 add_6412_8_lut (.I0(GND_net), .I1(n18086[5]), .I2(n533), .I3(n59677), 
            .O(n17578[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_8 (.CI(n59677), .I0(n18086[5]), .I1(n533), .CO(n59678));
    SB_LUT4 add_6412_7_lut (.I0(GND_net), .I1(n18086[4]), .I2(n460_c), 
            .I3(n59676), .O(n17578[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_7 (.CI(n59676), .I0(n18086[4]), .I1(n460_c), .CO(n59677));
    SB_LUT4 add_6412_6_lut (.I0(GND_net), .I1(n18086[3]), .I2(n387_adj_4591), 
            .I3(n59675), .O(n17578[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_6 (.CI(n59675), .I0(n18086[3]), .I1(n387_adj_4591), 
            .CO(n59676));
    SB_LUT4 add_6412_5_lut (.I0(GND_net), .I1(n18086[2]), .I2(n314_adj_4592), 
            .I3(n59674), .O(n17578[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_5 (.CI(n59674), .I0(n18086[2]), .I1(n314_adj_4592), 
            .CO(n59675));
    SB_LUT4 add_6412_4_lut (.I0(GND_net), .I1(n18086[1]), .I2(n241_adj_4593), 
            .I3(n59673), .O(n17578[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_4 (.CI(n59673), .I0(n18086[1]), .I1(n241_adj_4593), 
            .CO(n59674));
    SB_LUT4 add_6412_3_lut (.I0(GND_net), .I1(n18086[0]), .I2(n168_adj_4594), 
            .I3(n59672), .O(n17578[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_3 (.CI(n59672), .I0(n18086[0]), .I1(n168_adj_4594), 
            .CO(n59673));
    SB_LUT4 add_6412_2_lut (.I0(GND_net), .I1(n26_adj_4595), .I2(n95_adj_4596), 
            .I3(GND_net), .O(n17578[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6412_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6412_2 (.CI(GND_net), .I0(n26_adj_4595), .I1(n95_adj_4596), 
            .CO(n59672));
    SB_LUT4 add_6442_16_lut (.I0(GND_net), .I1(n18532[13]), .I2(n1120_adj_4597), 
            .I3(n59671), .O(n18086[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_15_lut (.I0(GND_net), .I1(n18532[12]), .I2(n1047_adj_4598), 
            .I3(n59670), .O(n18086[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_15 (.CI(n59670), .I0(n18532[12]), .I1(n1047_adj_4598), 
            .CO(n59671));
    SB_LUT4 add_6442_14_lut (.I0(GND_net), .I1(n18532[11]), .I2(n974_adj_4599), 
            .I3(n59669), .O(n18086[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_14 (.CI(n59669), .I0(n18532[11]), .I1(n974_adj_4599), 
            .CO(n59670));
    SB_LUT4 add_6442_13_lut (.I0(GND_net), .I1(n18532[10]), .I2(n901_adj_4600), 
            .I3(n59668), .O(n18086[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_13 (.CI(n59668), .I0(n18532[10]), .I1(n901_adj_4600), 
            .CO(n59669));
    SB_LUT4 n11880_bdd_4_lut_62805 (.I0(n11880), .I1(n74596), .I2(setpoint[4]), 
            .I3(n4734), .O(n78669));
    defparam n11880_bdd_4_lut_62805.LUT_INIT = 16'he4aa;
    SB_DFFSR counter_2045_2046__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4601));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4602));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78669_bdd_4_lut (.I0(n78669), .I1(n535[4]), .I2(n475), .I3(n4734), 
            .O(n78672));
    defparam n78669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_6442_12_lut (.I0(GND_net), .I1(n18532[9]), .I2(n828_adj_4604), 
            .I3(n59667), .O(n18086[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_12 (.CI(n59667), .I0(n18532[9]), .I1(n828_adj_4604), 
            .CO(n59668));
    SB_DFFSR counter_2045_2046__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 add_6442_11_lut (.I0(GND_net), .I1(n18532[8]), .I2(n755_adj_4607), 
            .I3(n59666), .O(n18086[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_11 (.CI(n59666), .I0(n18532[8]), .I1(n755_adj_4607), 
            .CO(n59667));
    SB_LUT4 add_6442_10_lut (.I0(GND_net), .I1(n18532[7]), .I2(n682_adj_4608), 
            .I3(n59665), .O(n18086[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_10 (.CI(n59665), .I0(n18532[7]), .I1(n682_adj_4608), 
            .CO(n59666));
    SB_LUT4 n11880_bdd_4_lut_62800 (.I0(n11880), .I1(n74595), .I2(setpoint[3]), 
            .I3(n4734), .O(n78663));
    defparam n11880_bdd_4_lut_62800.LUT_INIT = 16'he4aa;
    SB_LUT4 add_6562_9_lut (.I0(GND_net), .I1(n19972[6]), .I2(n624_adj_4609), 
            .I3(n58879), .O(n19776[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6442_9_lut (.I0(GND_net), .I1(n18532[6]), .I2(n609_adj_4610), 
            .I3(n59664), .O(n18086[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_9 (.CI(n59664), .I0(n18532[6]), .I1(n609_adj_4610), 
            .CO(n59665));
    SB_LUT4 add_6442_8_lut (.I0(GND_net), .I1(n18532[5]), .I2(n536_adj_4611), 
            .I3(n59663), .O(n18086[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_8 (.CI(n59663), .I0(n18532[5]), .I1(n536_adj_4611), 
            .CO(n59664));
    SB_LUT4 add_6442_7_lut (.I0(GND_net), .I1(n18532[4]), .I2(n463_adj_4612), 
            .I3(n59662), .O(n18086[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_7 (.CI(n59662), .I0(n18532[4]), .I1(n463_adj_4612), 
            .CO(n59663));
    SB_LUT4 add_6442_6_lut (.I0(GND_net), .I1(n18532[3]), .I2(n390_adj_4613), 
            .I3(n59661), .O(n18086[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_6 (.CI(n59661), .I0(n18532[3]), .I1(n390_adj_4613), 
            .CO(n59662));
    SB_LUT4 add_6442_5_lut (.I0(GND_net), .I1(n18532[2]), .I2(n317_adj_4614), 
            .I3(n59660), .O(n18086[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_9 (.CI(n58879), .I0(n19972[6]), .I1(n624_adj_4609), 
            .CO(n58880));
    SB_CARRY add_6442_5 (.CI(n59660), .I0(n18532[2]), .I1(n317_adj_4614), 
            .CO(n59661));
    SB_LUT4 add_6442_4_lut (.I0(GND_net), .I1(n18532[1]), .I2(n244_adj_4615), 
            .I3(n59659), .O(n18086[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n78663_bdd_4_lut (.I0(n78663), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4734), .O(n78666));
    defparam n78663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_6442_4 (.CI(n59659), .I0(n18532[1]), .I1(n244_adj_4615), 
            .CO(n59660));
    SB_LUT4 add_6442_3_lut (.I0(GND_net), .I1(n18532[0]), .I2(n171_adj_4616), 
            .I3(n59658), .O(n18086[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_3 (.CI(n59658), .I0(n18532[0]), .I1(n171_adj_4616), 
            .CO(n59659));
    SB_LUT4 add_6442_2_lut (.I0(GND_net), .I1(n29_adj_4617), .I2(n98_adj_4618), 
            .I3(GND_net), .O(n18086[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6442_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6442_2 (.CI(GND_net), .I0(n29_adj_4617), .I1(n98_adj_4618), 
            .CO(n59658));
    SB_LUT4 add_6586_9_lut (.I0(GND_net), .I1(n20176[6]), .I2(n630), .I3(n59657), 
            .O(n20033[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_8_lut (.I0(GND_net), .I1(n19972[5]), .I2(n551_adj_4619), 
            .I3(n58878), .O(n19776[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_8 (.CI(n58878), .I0(n19972[5]), .I1(n551_adj_4619), 
            .CO(n58879));
    SB_LUT4 add_6586_8_lut (.I0(GND_net), .I1(n20176[5]), .I2(n557), .I3(n59656), 
            .O(n20033[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_8 (.CI(n59656), .I0(n20176[5]), .I1(n557), .CO(n59657));
    SB_LUT4 add_6586_7_lut (.I0(GND_net), .I1(n20176[4]), .I2(n484), .I3(n59655), 
            .O(n20033[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_7 (.CI(n59655), .I0(n20176[4]), .I1(n484), .CO(n59656));
    SB_LUT4 add_6562_7_lut (.I0(GND_net), .I1(n19972[4]), .I2(n478_adj_4620), 
            .I3(n58877), .O(n19776[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_7 (.CI(n58877), .I0(n19972[4]), .I1(n478_adj_4620), 
            .CO(n58878));
    SB_LUT4 add_6586_6_lut (.I0(GND_net), .I1(n20176[3]), .I2(n411), .I3(n59654), 
            .O(n20033[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_6_lut (.I0(GND_net), .I1(n19972[3]), .I2(n405_adj_4621), 
            .I3(n58876), .O(n19776[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_6 (.CI(n59654), .I0(n20176[3]), .I1(n411), .CO(n59655));
    SB_CARRY add_6562_6 (.CI(n58876), .I0(n19972[3]), .I1(n405_adj_4621), 
            .CO(n58877));
    SB_LUT4 add_6586_5_lut (.I0(GND_net), .I1(n20176[2]), .I2(n338), .I3(n59653), 
            .O(n20033[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_5 (.CI(n59653), .I0(n20176[2]), .I1(n338), .CO(n59654));
    SB_LUT4 add_6586_4_lut (.I0(GND_net), .I1(n20176[1]), .I2(n265), .I3(n59652), 
            .O(n20033[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6562_5_lut (.I0(GND_net), .I1(n19972[2]), .I2(n332_adj_4622), 
            .I3(n58875), .O(n19776[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_5 (.CI(n58875), .I0(n19972[2]), .I1(n332_adj_4622), 
            .CO(n58876));
    SB_LUT4 add_6562_4_lut (.I0(GND_net), .I1(n19972[1]), .I2(n259_adj_4623), 
            .I3(n58874), .O(n19776[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_4 (.CI(n58874), .I0(n19972[1]), .I1(n259_adj_4623), 
            .CO(n58875));
    SB_CARRY add_6586_4 (.CI(n59652), .I0(n20176[1]), .I1(n265), .CO(n59653));
    SB_LUT4 add_6586_3_lut (.I0(GND_net), .I1(n20176[0]), .I2(n192), .I3(n59651), 
            .O(n20033[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6586_3 (.CI(n59651), .I0(n20176[0]), .I1(n192), .CO(n59652));
    SB_LUT4 add_6562_3_lut (.I0(GND_net), .I1(n19972[0]), .I2(n186_adj_4624), 
            .I3(n58873), .O(n19776[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6586_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20033[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6586_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_3 (.CI(n58873), .I0(n19972[0]), .I1(n186_adj_4624), 
            .CO(n58874));
    SB_CARRY add_6586_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n59651));
    SB_LUT4 add_6562_2_lut (.I0(GND_net), .I1(n44_adj_4625), .I2(n113_adj_4626), 
            .I3(GND_net), .O(n19776[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6562_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6470_15_lut (.I0(GND_net), .I1(n18920[12]), .I2(n1050_adj_4627), 
            .I3(n59650), .O(n18532[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6470_14_lut (.I0(GND_net), .I1(n18920[11]), .I2(n977_adj_4628), 
            .I3(n59649), .O(n18532[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6562_2 (.CI(GND_net), .I0(n44_adj_4625), .I1(n113_adj_4626), 
            .CO(n58873));
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4628));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6470_14 (.CI(n59649), .I0(n18920[11]), .I1(n977_adj_4628), 
            .CO(n59650));
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n345));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6470_13_lut (.I0(GND_net), .I1(n18920[10]), .I2(n904), 
            .I3(n59648), .O(n18532[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4626));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4625));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_13 (.CI(n59648), .I0(n18920[10]), .I1(n904), .CO(n59649));
    SB_LUT4 add_6470_12_lut (.I0(GND_net), .I1(n18920[9]), .I2(n831), 
            .I3(n59647), .O(n18532[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_12 (.CI(n59647), .I0(n18920[9]), .I1(n831), .CO(n59648));
    SB_LUT4 add_6470_11_lut (.I0(GND_net), .I1(n18920[8]), .I2(n758), 
            .I3(n59646), .O(n18532[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_11 (.CI(n59646), .I0(n18920[8]), .I1(n758), .CO(n59647));
    SB_LUT4 add_6470_10_lut (.I0(GND_net), .I1(n18920[7]), .I2(n685), 
            .I3(n59645), .O(n18532[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_10 (.CI(n59645), .I0(n18920[7]), .I1(n685), .CO(n59646));
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_9_lut (.I0(GND_net), .I1(n18920[6]), .I2(n612), .I3(n59644), 
            .O(n18532[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30514), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30513), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30512), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30511), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30510), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_6470_9 (.CI(n59644), .I0(n18920[6]), .I1(n612), .CO(n59645));
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30509), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30508), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30507), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30506), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30505), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30503), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30501), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30500), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30499), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30498), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30497), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30496), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30495), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30494), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30493), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30488), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30487), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30479), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6470_8_lut (.I0(GND_net), .I1(n18920[5]), .I2(n539), .I3(n59643), 
            .O(n18532[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_8 (.CI(n59643), .I0(n18920[5]), .I1(n539), .CO(n59644));
    SB_LUT4 add_6470_7_lut (.I0(GND_net), .I1(n18920[4]), .I2(n466), .I3(n59642), 
            .O(n18532[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_7 (.CI(n59642), .I0(n18920[4]), .I1(n466), .CO(n59643));
    SB_LUT4 add_6470_6_lut (.I0(GND_net), .I1(n18920[3]), .I2(n393), .I3(n59641), 
            .O(n18532[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4623));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4631));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4632));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4633));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4622));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4634));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_6 (.CI(n59641), .I0(n18920[3]), .I1(n393), .CO(n59642));
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4635));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_5_lut (.I0(GND_net), .I1(n18920[2]), .I2(n320), .I3(n59640), 
            .O(n18532[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4636));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4637));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_5 (.CI(n59640), .I0(n18920[2]), .I1(n320), .CO(n59641));
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4638));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6470_4_lut (.I0(GND_net), .I1(n18920[1]), .I2(n247_c), 
            .I3(n59639), .O(n18532[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_4 (.CI(n59639), .I0(n18920[1]), .I1(n247_c), .CO(n59640));
    SB_LUT4 add_6470_3_lut (.I0(GND_net), .I1(n18920[0]), .I2(n174), .I3(n59638), 
            .O(n18532[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6470_3 (.CI(n59638), .I0(n18920[0]), .I1(n174), .CO(n59639));
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6470_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18532[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6470_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6470_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n59638));
    SB_LUT4 add_6496_14_lut (.I0(GND_net), .I1(n19254[11]), .I2(n980), 
            .I3(n59637), .O(n18920[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4621));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6496_13_lut (.I0(GND_net), .I1(n19254[10]), .I2(n907), 
            .I3(n59636), .O(n18920[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_13 (.CI(n59636), .I0(n19254[10]), .I1(n907), .CO(n59637));
    SB_LUT4 add_6496_12_lut (.I0(GND_net), .I1(n19254[9]), .I2(n834), 
            .I3(n59635), .O(n18920[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_12 (.CI(n59635), .I0(n19254[9]), .I1(n834), .CO(n59636));
    SB_LUT4 add_6496_11_lut (.I0(GND_net), .I1(n19254[8]), .I2(n761), 
            .I3(n59634), .O(n18920[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_11 (.CI(n59634), .I0(n19254[8]), .I1(n761), .CO(n59635));
    SB_LUT4 add_6496_10_lut (.I0(GND_net), .I1(n19254[7]), .I2(n688), 
            .I3(n59633), .O(n18920[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31093_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45170));   // verilog/motorControl.v(61[20:40])
    defparam i31093_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6496_10 (.CI(n59633), .I0(n19254[7]), .I1(n688), .CO(n59634));
    SB_LUT4 add_6496_9_lut (.I0(GND_net), .I1(n19254[6]), .I2(n615_adj_4645), 
            .I3(n59632), .O(n18920[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_9 (.CI(n59632), .I0(n19254[6]), .I1(n615_adj_4645), 
            .CO(n59633));
    SB_LUT4 add_6139_23_lut (.I0(GND_net), .I1(n13441[20]), .I2(GND_net), 
            .I3(n58850), .O(n12379[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6496_8_lut (.I0(GND_net), .I1(n19254[5]), .I2(n542_adj_4646), 
            .I3(n59631), .O(n18920[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6496_8 (.CI(n59631), .I0(n19254[5]), .I1(n542_adj_4646), 
            .CO(n59632));
    SB_LUT4 add_6139_22_lut (.I0(GND_net), .I1(n13441[19]), .I2(GND_net), 
            .I3(n58849), .O(n12379[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_22 (.CI(n58849), .I0(n13441[19]), .I1(GND_net), 
            .CO(n58850));
    SB_LUT4 add_6139_21_lut (.I0(GND_net), .I1(n13441[18]), .I2(GND_net), 
            .I3(n58848), .O(n12379[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_21 (.CI(n58848), .I0(n13441[18]), .I1(GND_net), 
            .CO(n58849));
    SB_LUT4 add_6139_20_lut (.I0(GND_net), .I1(n13441[17]), .I2(GND_net), 
            .I3(n58847), .O(n12379[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_20 (.CI(n58847), .I0(n13441[17]), .I1(GND_net), 
            .CO(n58848));
    SB_LUT4 add_6139_19_lut (.I0(GND_net), .I1(n13441[16]), .I2(GND_net), 
            .I3(n58846), .O(n12379[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_19 (.CI(n58846), .I0(n13441[16]), .I1(GND_net), 
            .CO(n58847));
    SB_LUT4 add_6506_13_lut (.I0(GND_net), .I1(n19372[10]), .I2(n910_adj_4647), 
            .I3(n58438), .O(n19061[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6139_18_lut (.I0(GND_net), .I1(n13441[15]), .I2(GND_net), 
            .I3(n58845), .O(n12379[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_18 (.CI(n58845), .I0(n13441[15]), .I1(GND_net), 
            .CO(n58846));
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29773), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6139_17_lut (.I0(GND_net), .I1(n13441[14]), .I2(GND_net), 
            .I3(n58844), .O(n12379[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6496_7_lut (.I0(GND_net), .I1(n19254[4]), .I2(n469_adj_4648), 
            .I3(n59630), .O(n18920[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_7 (.CI(n59630), .I0(n19254[4]), .I1(n469_adj_4648), 
            .CO(n59631));
    SB_CARRY add_6139_17 (.CI(n58844), .I0(n13441[14]), .I1(GND_net), 
            .CO(n58845));
    SB_LUT4 add_6139_16_lut (.I0(GND_net), .I1(n13441[13]), .I2(n1099_adj_4649), 
            .I3(n58843), .O(n12379[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_16 (.CI(n58843), .I0(n13441[13]), .I1(n1099_adj_4649), 
            .CO(n58844));
    SB_LUT4 add_6506_12_lut (.I0(GND_net), .I1(n19372[9]), .I2(n837_adj_4650), 
            .I3(n58437), .O(n19061[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_12 (.CI(n58437), .I0(n19372[9]), .I1(n837_adj_4650), 
            .CO(n58438));
    SB_LUT4 add_6139_15_lut (.I0(GND_net), .I1(n13441[12]), .I2(n1026_adj_4651), 
            .I3(n58842), .O(n12379[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_15 (.CI(n58842), .I0(n13441[12]), .I1(n1026_adj_4651), 
            .CO(n58843));
    SB_LUT4 add_6506_11_lut (.I0(GND_net), .I1(n19372[8]), .I2(n764_adj_4652), 
            .I3(n58436), .O(n19061[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_11 (.CI(n58436), .I0(n19372[8]), .I1(n764_adj_4652), 
            .CO(n58437));
    SB_LUT4 add_6139_14_lut (.I0(GND_net), .I1(n13441[11]), .I2(n953_adj_4653), 
            .I3(n58841), .O(n12379[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_14 (.CI(n58841), .I0(n13441[11]), .I1(n953_adj_4653), 
            .CO(n58842));
    SB_LUT4 add_6506_10_lut (.I0(GND_net), .I1(n19372[7]), .I2(n691_adj_4654), 
            .I3(n58435), .O(n19061[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_10 (.CI(n58435), .I0(n19372[7]), .I1(n691_adj_4654), 
            .CO(n58436));
    SB_LUT4 add_6139_13_lut (.I0(GND_net), .I1(n13441[10]), .I2(n880_adj_4655), 
            .I3(n58840), .O(n12379[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_13 (.CI(n58840), .I0(n13441[10]), .I1(n880_adj_4655), 
            .CO(n58841));
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n78654), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_6506_9_lut (.I0(GND_net), .I1(n19372[6]), .I2(n618_adj_4656), 
            .I3(n58434), .O(n19061[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_9 (.CI(n58434), .I0(n19372[6]), .I1(n618_adj_4656), 
            .CO(n58435));
    SB_LUT4 add_6139_12_lut (.I0(GND_net), .I1(n13441[9]), .I2(n807_adj_4657), 
            .I3(n58839), .O(n12379[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_12 (.CI(n58839), .I0(n13441[9]), .I1(n807_adj_4657), 
            .CO(n58840));
    SB_LUT4 add_6139_11_lut (.I0(GND_net), .I1(n13441[8]), .I2(n734_adj_4658), 
            .I3(n58838), .O(n12379[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_11 (.CI(n58838), .I0(n13441[8]), .I1(n734_adj_4658), 
            .CO(n58839));
    SB_LUT4 add_6139_10_lut (.I0(GND_net), .I1(n13441[7]), .I2(n661_adj_4659), 
            .I3(n58837), .O(n12379[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_10 (.CI(n58837), .I0(n13441[7]), .I1(n661_adj_4659), 
            .CO(n58838));
    SB_LUT4 add_6506_8_lut (.I0(GND_net), .I1(n19372[5]), .I2(n545_adj_4660), 
            .I3(n58433), .O(n19061[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_8 (.CI(n58433), .I0(n19372[5]), .I1(n545_adj_4660), 
            .CO(n58434));
    SB_LUT4 add_6139_9_lut (.I0(GND_net), .I1(n13441[6]), .I2(n588_adj_4661), 
            .I3(n58836), .O(n12379[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4620));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6139_9 (.CI(n58836), .I0(n13441[6]), .I1(n588_adj_4661), 
            .CO(n58837));
    SB_LUT4 add_6506_7_lut (.I0(GND_net), .I1(n19372[4]), .I2(n472_adj_4662), 
            .I3(n58432), .O(n19061[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_7 (.CI(n58432), .I0(n19372[4]), .I1(n472_adj_4662), 
            .CO(n58433));
    SB_LUT4 add_6139_8_lut (.I0(GND_net), .I1(n13441[5]), .I2(n515_adj_4663), 
            .I3(n58835), .O(n12379[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_8 (.CI(n58835), .I0(n13441[5]), .I1(n515_adj_4663), 
            .CO(n58836));
    SB_LUT4 add_6506_6_lut (.I0(GND_net), .I1(n19372[3]), .I2(n399_adj_4664), 
            .I3(n58431), .O(n19061[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_6 (.CI(n58431), .I0(n19372[3]), .I1(n399_adj_4664), 
            .CO(n58432));
    SB_LUT4 add_6139_7_lut (.I0(GND_net), .I1(n13441[4]), .I2(n442_adj_4665), 
            .I3(n58834), .O(n12379[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_7 (.CI(n58834), .I0(n13441[4]), .I1(n442_adj_4665), 
            .CO(n58835));
    SB_LUT4 add_6506_5_lut (.I0(GND_net), .I1(n19372[2]), .I2(n326_adj_4666), 
            .I3(n58430), .O(n19061[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_5 (.CI(n58430), .I0(n19372[2]), .I1(n326_adj_4666), 
            .CO(n58431));
    SB_LUT4 add_6139_6_lut (.I0(GND_net), .I1(n13441[3]), .I2(n369_adj_4667), 
            .I3(n58833), .O(n12379[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_6 (.CI(n58833), .I0(n13441[3]), .I1(n369_adj_4667), 
            .CO(n58834));
    SB_LUT4 add_6139_5_lut (.I0(GND_net), .I1(n13441[2]), .I2(n296_adj_4668), 
            .I3(n58832), .O(n12379[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_5 (.CI(n58832), .I0(n13441[2]), .I1(n296_adj_4668), 
            .CO(n58833));
    SB_LUT4 add_6139_4_lut (.I0(GND_net), .I1(n13441[1]), .I2(n223_adj_4669), 
            .I3(n58831), .O(n12379[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6139_4 (.CI(n58831), .I0(n13441[1]), .I1(n223_adj_4669), 
            .CO(n58832));
    SB_LUT4 add_6139_3_lut (.I0(GND_net), .I1(n13441[0]), .I2(n150_adj_4670), 
            .I3(n58830), .O(n12379[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6496_6_lut (.I0(GND_net), .I1(n19254[3]), .I2(n396_adj_4671), 
            .I3(n59629), .O(n18920[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_3 (.CI(n58830), .I0(n13441[0]), .I1(n150_adj_4670), 
            .CO(n58831));
    SB_CARRY add_6496_6 (.CI(n59629), .I0(n19254[3]), .I1(n396_adj_4671), 
            .CO(n59630));
    SB_LUT4 add_6139_2_lut (.I0(GND_net), .I1(n8_adj_4672), .I2(n77_adj_4673), 
            .I3(GND_net), .O(n12379[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6139_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6139_2 (.CI(GND_net), .I0(n8_adj_4672), .I1(n77_adj_4673), 
            .CO(n58830));
    SB_LUT4 add_6506_4_lut (.I0(GND_net), .I1(n19372[1]), .I2(n253_adj_4674), 
            .I3(n58429), .O(n19061[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_4 (.CI(n58429), .I0(n19372[1]), .I1(n253_adj_4674), 
            .CO(n58430));
    SB_LUT4 add_6208_22_lut (.I0(GND_net), .I1(n14365[19]), .I2(GND_net), 
            .I3(n58829), .O(n13441[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_21_lut (.I0(GND_net), .I1(n14365[18]), .I2(GND_net), 
            .I3(n58828), .O(n13441[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_3_lut (.I0(GND_net), .I1(n19372[0]), .I2(n180_adj_4675), 
            .I3(n58428), .O(n19061[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_3 (.CI(n58428), .I0(n19372[0]), .I1(n180_adj_4675), 
            .CO(n58429));
    SB_LUT4 add_6496_5_lut (.I0(GND_net), .I1(n19254[2]), .I2(n323_adj_4676), 
            .I3(n59628), .O(n18920[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_21 (.CI(n58828), .I0(n14365[18]), .I1(GND_net), 
            .CO(n58829));
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6208_20_lut (.I0(GND_net), .I1(n14365[17]), .I2(GND_net), 
            .I3(n58827), .O(n13441[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6506_2_lut (.I0(GND_net), .I1(n38_c), .I2(n107_adj_4677), 
            .I3(GND_net), .O(n19061[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6506_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6506_2 (.CI(GND_net), .I0(n38_c), .I1(n107_adj_4677), 
            .CO(n58428));
    SB_CARRY add_6208_20 (.CI(n58827), .I0(n14365[17]), .I1(GND_net), 
            .CO(n58828));
    SB_LUT4 add_6208_19_lut (.I0(GND_net), .I1(n14365[16]), .I2(GND_net), 
            .I3(n58826), .O(n13441[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_19 (.CI(n58826), .I0(n14365[16]), .I1(GND_net), 
            .CO(n58827));
    SB_LUT4 add_6208_18_lut (.I0(GND_net), .I1(n14365[15]), .I2(GND_net), 
            .I3(n58825), .O(n13441[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_18 (.CI(n58825), .I0(n14365[15]), .I1(GND_net), 
            .CO(n58826));
    SB_LUT4 add_6208_17_lut (.I0(GND_net), .I1(n14365[14]), .I2(GND_net), 
            .I3(n58824), .O(n13441[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_17 (.CI(n58824), .I0(n14365[14]), .I1(GND_net), 
            .CO(n58825));
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6496_5 (.CI(n59628), .I0(n19254[2]), .I1(n323_adj_4676), 
            .CO(n59629));
    SB_LUT4 add_6208_16_lut (.I0(GND_net), .I1(n14365[13]), .I2(n1102_adj_4680), 
            .I3(n58823), .O(n13441[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_16 (.CI(n58823), .I0(n14365[13]), .I1(n1102_adj_4680), 
            .CO(n58824));
    SB_LUT4 add_6208_15_lut (.I0(GND_net), .I1(n14365[12]), .I2(n1029_adj_4681), 
            .I3(n58822), .O(n13441[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4619));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6208_15 (.CI(n58822), .I0(n14365[12]), .I1(n1029_adj_4681), 
            .CO(n58823));
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6208_14_lut (.I0(GND_net), .I1(n14365[11]), .I2(n956_adj_4683), 
            .I3(n58821), .O(n13441[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_14 (.CI(n58821), .I0(n14365[11]), .I1(n956_adj_4683), 
            .CO(n58822));
    SB_LUT4 add_6208_13_lut (.I0(GND_net), .I1(n14365[10]), .I2(n883_adj_4684), 
            .I3(n58820), .O(n13441[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_13 (.CI(n58820), .I0(n14365[10]), .I1(n883_adj_4684), 
            .CO(n58821));
    SB_LUT4 add_6496_4_lut (.I0(GND_net), .I1(n19254[1]), .I2(n250_adj_4685), 
            .I3(n59627), .O(n18920[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_12_lut (.I0(GND_net), .I1(n14365[9]), .I2(n810_adj_4686), 
            .I3(n58819), .O(n13441[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_12 (.CI(n58819), .I0(n14365[9]), .I1(n810_adj_4686), 
            .CO(n58820));
    SB_LUT4 add_6208_11_lut (.I0(GND_net), .I1(n14365[8]), .I2(n737_adj_4687), 
            .I3(n58818), .O(n13441[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_4 (.CI(n59627), .I0(n19254[1]), .I1(n250_adj_4685), 
            .CO(n59628));
    SB_CARRY add_6208_11 (.CI(n58818), .I0(n14365[8]), .I1(n737_adj_4687), 
            .CO(n58819));
    SB_LUT4 add_6496_3_lut (.I0(GND_net), .I1(n19254[0]), .I2(n177_adj_4688), 
            .I3(n59626), .O(n18920[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6208_10_lut (.I0(GND_net), .I1(n14365[7]), .I2(n664_adj_4689), 
            .I3(n58817), .O(n13441[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_10 (.CI(n58817), .I0(n14365[7]), .I1(n664_adj_4689), 
            .CO(n58818));
    SB_LUT4 add_6208_9_lut (.I0(GND_net), .I1(n14365[6]), .I2(n591_adj_4690), 
            .I3(n58816), .O(n13441[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_9 (.CI(n58816), .I0(n14365[6]), .I1(n591_adj_4690), 
            .CO(n58817));
    SB_LUT4 add_6208_8_lut (.I0(GND_net), .I1(n14365[5]), .I2(n518_adj_4691), 
            .I3(n58815), .O(n13441[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_8 (.CI(n58815), .I0(n14365[5]), .I1(n518_adj_4691), 
            .CO(n58816));
    SB_LUT4 add_6208_7_lut (.I0(GND_net), .I1(n14365[4]), .I2(n445_adj_4692), 
            .I3(n58814), .O(n13441[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_7 (.CI(n58814), .I0(n14365[4]), .I1(n445_adj_4692), 
            .CO(n58815));
    SB_LUT4 add_6208_6_lut (.I0(GND_net), .I1(n14365[3]), .I2(n372_adj_4693), 
            .I3(n58813), .O(n13441[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_6 (.CI(n58813), .I0(n14365[3]), .I1(n372_adj_4693), 
            .CO(n58814));
    SB_LUT4 add_6208_5_lut (.I0(GND_net), .I1(n14365[2]), .I2(n299_adj_4694), 
            .I3(n58812), .O(n13441[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_3 (.CI(n59626), .I0(n19254[0]), .I1(n177_adj_4688), 
            .CO(n59627));
    SB_LUT4 add_6496_2_lut (.I0(GND_net), .I1(n35_adj_4695), .I2(n104_adj_4696), 
            .I3(GND_net), .O(n18920[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6496_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6496_2 (.CI(GND_net), .I0(n35_adj_4695), .I1(n104_adj_4696), 
            .CO(n59626));
    SB_CARRY add_6208_5 (.CI(n58812), .I0(n14365[2]), .I1(n299_adj_4694), 
            .CO(n58813));
    SB_LUT4 add_6208_4_lut (.I0(GND_net), .I1(n14365[1]), .I2(n226_adj_4697), 
            .I3(n58811), .O(n13441[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_4 (.CI(n58811), .I0(n14365[1]), .I1(n226_adj_4697), 
            .CO(n58812));
    SB_LUT4 add_6208_3_lut (.I0(GND_net), .I1(n14365[0]), .I2(n153_adj_4698), 
            .I3(n58810), .O(n13441[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_3 (.CI(n58810), .I0(n14365[0]), .I1(n153_adj_4698), 
            .CO(n58811));
    SB_LUT4 add_6208_2_lut (.I0(GND_net), .I1(n11_adj_4699), .I2(n80_adj_4700), 
            .I3(GND_net), .O(n13441[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6208_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6208_2 (.CI(GND_net), .I0(n11_adj_4699), .I1(n80_adj_4700), 
            .CO(n58810));
    SB_LUT4 add_6601_8_lut (.I0(GND_net), .I1(n20287[5]), .I2(n560_adj_4701), 
            .I3(n59625), .O(n20176[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_7_lut (.I0(GND_net), .I1(n20287[4]), .I2(n487_adj_4702), 
            .I3(n59624), .O(n20176[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_7 (.CI(n59624), .I0(n20287[4]), .I1(n487_adj_4702), 
            .CO(n59625));
    SB_LUT4 add_6601_6_lut (.I0(GND_net), .I1(n20287[3]), .I2(n414_adj_4703), 
            .I3(n59623), .O(n20176[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4705));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n460), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_c));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_c));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4709));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n11880_bdd_4_lut (.I0(n11880), .I1(n74663), .I2(setpoint[23]), 
            .I3(n4734), .O(n78927));
    defparam n11880_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4711));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4712));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n467), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4713));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4714));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4715));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6601_6 (.CI(n59623), .I0(n20287[3]), .I1(n414_adj_4703), 
            .CO(n59624));
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n475), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4716));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6250_21_lut (.I0(GND_net), .I1(n15204[18]), .I2(GND_net), 
            .I3(n58788), .O(n14365[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_20_lut (.I0(GND_net), .I1(n15204[17]), .I2(GND_net), 
            .I3(n58787), .O(n14365[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_20 (.CI(n58787), .I0(n15204[17]), .I1(GND_net), 
            .CO(n58788));
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4719));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_c));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4721));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4722));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4723));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6250_19_lut (.I0(GND_net), .I1(n15204[16]), .I2(GND_net), 
            .I3(n58786), .O(n14365[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_19 (.CI(n58786), .I0(n15204[16]), .I1(GND_net), 
            .CO(n58787));
    SB_LUT4 add_6250_18_lut (.I0(GND_net), .I1(n15204[15]), .I2(GND_net), 
            .I3(n58785), .O(n14365[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_18 (.CI(n58785), .I0(n15204[15]), .I1(GND_net), 
            .CO(n58786));
    SB_LUT4 add_6250_17_lut (.I0(GND_net), .I1(n15204[14]), .I2(GND_net), 
            .I3(n58784), .O(n14365[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6250_17 (.CI(n58784), .I0(n15204[14]), .I1(GND_net), 
            .CO(n58785));
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n78927_bdd_4_lut (.I0(n78927), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4734), .O(n78930));
    defparam n78927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4727));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4728));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4729));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4730));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4731));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6250_16_lut (.I0(GND_net), .I1(n15204[13]), .I2(n1105_adj_4732), 
            .I3(n58783), .O(n14365[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4733));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6250_16 (.CI(n58783), .I0(n15204[13]), .I1(n1105_adj_4732), 
            .CO(n58784));
    SB_LUT4 add_6250_15_lut (.I0(GND_net), .I1(n15204[12]), .I2(n1032_adj_4734), 
            .I3(n58782), .O(n14365[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_15 (.CI(n58782), .I0(n15204[12]), .I1(n1032_adj_4734), 
            .CO(n58783));
    SB_LUT4 add_6250_14_lut (.I0(GND_net), .I1(n15204[11]), .I2(n959_adj_4735), 
            .I3(n58781), .O(n14365[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_14 (.CI(n58781), .I0(n15204[11]), .I1(n959_adj_4735), 
            .CO(n58782));
    SB_CARRY add_16_9 (.CI(n58197), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n58198));
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4736));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4737));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4738));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4739));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4740));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6250_13_lut (.I0(GND_net), .I1(n15204[10]), .I2(n886_adj_4741), 
            .I3(n58780), .O(n14365[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4742));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6250_13 (.CI(n58780), .I0(n15204[10]), .I1(n886_adj_4741), 
            .CO(n58781));
    SB_LUT4 add_6250_12_lut (.I0(GND_net), .I1(n15204[9]), .I2(n813_adj_4743), 
            .I3(n58779), .O(n14365[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_12 (.CI(n58779), .I0(n15204[9]), .I1(n813_adj_4743), 
            .CO(n58780));
    SB_LUT4 add_6250_11_lut (.I0(GND_net), .I1(n15204[8]), .I2(n740_adj_4744), 
            .I3(n58778), .O(n14365[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4745));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n58196), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_11 (.CI(n58778), .I0(n15204[8]), .I1(n740_adj_4744), 
            .CO(n58779));
    SB_LUT4 add_6601_5_lut (.I0(GND_net), .I1(n20287[2]), .I2(n341_adj_4746), 
            .I3(n59622), .O(n20176[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4747));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4748));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4749));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4750));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4751));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4752));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n105), .I1(control_update), .I2(n65754), .I3(n22), 
            .O(n25796));
    defparam i3_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 add_6250_10_lut (.I0(GND_net), .I1(n15204[7]), .I2(n667_adj_4754), 
            .I3(n58777), .O(n14365[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_10 (.CI(n58777), .I0(n15204[7]), .I1(n667_adj_4754), 
            .CO(n58778));
    SB_LUT4 add_6250_9_lut (.I0(GND_net), .I1(n15204[6]), .I2(n594_adj_4755), 
            .I3(n58776), .O(n14365[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_9 (.CI(n58776), .I0(n15204[6]), .I1(n594_adj_4755), 
            .CO(n58777));
    SB_LUT4 add_6250_8_lut (.I0(GND_net), .I1(n15204[5]), .I2(n521_adj_4756), 
            .I3(n58775), .O(n14365[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_8 (.CI(n58775), .I0(n15204[5]), .I1(n521_adj_4756), 
            .CO(n58776));
    SB_LUT4 add_6250_7_lut (.I0(GND_net), .I1(n15204[4]), .I2(n448_adj_4757), 
            .I3(n58774), .O(n14365[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59660_4_lut (.I0(n21_adj_4752), .I1(n19_adj_4751), .I2(n17_adj_4750), 
            .I3(n9_adj_4749), .O(n75495));
    defparam i59660_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59622_4_lut (.I0(n27_adj_4745), .I1(n15_adj_4747), .I2(n13_adj_4742), 
            .I3(n11_adj_4740), .O(n75457));
    defparam i59622_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4748), 
            .I3(GND_net), .O(n12_adj_4758));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4742), 
            .I3(GND_net), .O(n10_adj_4759));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4758), .I1(n535[17]), .I2(n35_adj_4739), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6250_7 (.CI(n58774), .I0(n15204[4]), .I1(n448_adj_4757), 
            .CO(n58775));
    SB_LUT4 add_6250_6_lut (.I0(GND_net), .I1(n15204[3]), .I2(n375_adj_4760), 
            .I3(n58773), .O(n14365[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_6 (.CI(n58773), .I0(n15204[3]), .I1(n375_adj_4760), 
            .CO(n58774));
    SB_LUT4 add_6250_5_lut (.I0(GND_net), .I1(n15204[2]), .I2(n302_adj_4761), 
            .I3(n58772), .O(n14365[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60574_4_lut (.I0(n13_adj_4742), .I1(n11_adj_4740), .I2(n9_adj_4749), 
            .I3(n75511), .O(n76409));
    defparam i60574_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60564_4_lut (.I0(n19_adj_4751), .I1(n17_adj_4750), .I2(n15_adj_4747), 
            .I3(n76409), .O(n76399));
    defparam i60564_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61552_4_lut (.I0(n25_adj_4738), .I1(n23_adj_4737), .I2(n21_adj_4752), 
            .I3(n76399), .O(n77387));
    defparam i61552_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i60959_4_lut (.I0(n31_adj_4736), .I1(n29_adj_4733), .I2(n27_adj_4745), 
            .I3(n77387), .O(n76794));
    defparam i60959_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61668_4_lut (.I0(n37_adj_4731), .I1(n35_adj_4739), .I2(n33_adj_4748), 
            .I3(n76794), .O(n77503));
    defparam i61668_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4730), 
            .I3(GND_net), .O(n16_adj_4762));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61274_3_lut (.I0(n6_adj_4763), .I1(n535[10]), .I2(n21_adj_4752), 
            .I3(GND_net), .O(n77109));   // verilog/motorControl.v(47[25:43])
    defparam i61274_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6250_5 (.CI(n58772), .I0(n15204[2]), .I1(n302_adj_4761), 
            .CO(n58773));
    SB_LUT4 add_6250_4_lut (.I0(GND_net), .I1(n15204[1]), .I2(n229_adj_4764), 
            .I3(n58771), .O(n14365[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_4 (.CI(n58771), .I0(n15204[1]), .I1(n229_adj_4764), 
            .CO(n58772));
    SB_LUT4 add_6250_3_lut (.I0(GND_net), .I1(n15204[0]), .I2(n156_adj_4765), 
            .I3(n58770), .O(n14365[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61275_3_lut (.I0(n77109), .I1(n535[11]), .I2(n23_adj_4737), 
            .I3(GND_net), .O(n77110));   // verilog/motorControl.v(47[25:43])
    defparam i61275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4750), 
            .I3(GND_net), .O(n8_adj_4766));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4762), .I1(n535[22]), .I2(n45_adj_4729), 
            .I3(GND_net), .O(n24_adj_4767));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59586_4_lut (.I0(n43_adj_4730), .I1(n25_adj_4738), .I2(n23_adj_4737), 
            .I3(n75495), .O(n75421));
    defparam i59586_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61065_4_lut (.I0(n24_adj_4767), .I1(n8_adj_4766), .I2(n45_adj_4729), 
            .I3(n75410), .O(n76900));   // verilog/motorControl.v(47[25:43])
    defparam i61065_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59974_3_lut (.I0(n77110), .I1(n535[12]), .I2(n25_adj_4738), 
            .I3(GND_net), .O(n75809));   // verilog/motorControl.v(47[25:43])
    defparam i59974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4768));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_6250_3 (.CI(n58770), .I0(n15204[0]), .I1(n156_adj_4765), 
            .CO(n58771));
    SB_LUT4 add_6250_2_lut (.I0(GND_net), .I1(n14_adj_4769), .I2(n83_adj_4770), 
            .I3(GND_net), .O(n14365[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6250_2 (.CI(GND_net), .I0(n14_adj_4769), .I1(n83_adj_4770), 
            .CO(n58770));
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4772));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4773));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6601_5 (.CI(n59622), .I0(n20287[2]), .I1(n341_adj_4746), 
            .CO(n59623));
    SB_LUT4 add_6601_4_lut (.I0(GND_net), .I1(n20287[1]), .I2(n268_adj_4775), 
            .I3(n59621), .O(n20176[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4776));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6601_4 (.CI(n59621), .I0(n20287[1]), .I1(n268_adj_4775), 
            .CO(n59622));
    SB_LUT4 add_6601_3_lut (.I0(GND_net), .I1(n20287[0]), .I2(n195_adj_4777), 
            .I3(n59620), .O(n20176[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4778));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61272_3_lut (.I0(n4_adj_4768), .I1(n535[13]), .I2(n27_adj_4745), 
            .I3(GND_net), .O(n77107));   // verilog/motorControl.v(47[25:43])
    defparam i61272_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_16_8 (.CI(n58196), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n58197));
    SB_CARRY add_6601_3 (.CI(n59620), .I0(n20287[0]), .I1(n195_adj_4777), 
            .CO(n59621));
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4779));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61273_3_lut (.I0(n77107), .I1(n535[14]), .I2(n29_adj_4733), 
            .I3(GND_net), .O(n77108));   // verilog/motorControl.v(47[25:43])
    defparam i61273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6601_2_lut (.I0(GND_net), .I1(n53_adj_4780), .I2(n122_adj_4781), 
            .I3(GND_net), .O(n20176[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4782));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59609_4_lut (.I0(n33_adj_4748), .I1(n31_adj_4736), .I2(n29_adj_4733), 
            .I3(n75457), .O(n75444));
    defparam i59609_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6601_2 (.CI(GND_net), .I0(n53_adj_4780), .I1(n122_adj_4781), 
            .CO(n59620));
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4783));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i61612_4_lut (.I0(n30), .I1(n10_adj_4759), .I2(n35_adj_4739), 
            .I3(n75440), .O(n77447));   // verilog/motorControl.v(47[25:43])
    defparam i61612_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n350));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59976_3_lut (.I0(n77108), .I1(n535[15]), .I2(n31_adj_4736), 
            .I3(GND_net), .O(n75811));   // verilog/motorControl.v(47[25:43])
    defparam i59976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61772_4_lut (.I0(n75811), .I1(n77447), .I2(n35_adj_4739), 
            .I3(n75444), .O(n77607));   // verilog/motorControl.v(47[25:43])
    defparam i61772_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4785));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4617));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4786));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61773_3_lut (.I0(n77607), .I1(n535[18]), .I2(n37_adj_4731), 
            .I3(GND_net), .O(n77608));   // verilog/motorControl.v(47[25:43])
    defparam i61773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4787));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4616));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_13_lut (.I0(GND_net), .I1(n19538[10]), .I2(n910), 
            .I3(n59619), .O(n19254[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4615));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4788));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4791));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4793));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4794));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61722_3_lut (.I0(n77608), .I1(n535[19]), .I2(n39_adj_4728), 
            .I3(GND_net), .O(n77557));   // verilog/motorControl.v(47[25:43])
    defparam i61722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6520_12_lut (.I0(GND_net), .I1(n19538[9]), .I2(n837), 
            .I3(n59618), .O(n19254[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_12 (.CI(n59618), .I0(n19538[9]), .I1(n837), .CO(n59619));
    SB_LUT4 add_6520_11_lut (.I0(GND_net), .I1(n19538[8]), .I2(n764), 
            .I3(n59617), .O(n19254[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_11 (.CI(n59617), .I0(n19538[8]), .I1(n764), .CO(n59618));
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4795));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_10_lut (.I0(GND_net), .I1(n19538[7]), .I2(n691), 
            .I3(n59616), .O(n19254[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59592_4_lut (.I0(n43_adj_4730), .I1(n41_adj_4727), .I2(n39_adj_4728), 
            .I3(n77503), .O(n75427));
    defparam i59592_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6520_10 (.CI(n59616), .I0(n19538[7]), .I1(n691), .CO(n59617));
    SB_LUT4 add_6520_9_lut (.I0(GND_net), .I1(n19538[6]), .I2(n618), .I3(n59615), 
            .O(n19254[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_9 (.CI(n59615), .I0(n19538[6]), .I1(n618), .CO(n59616));
    SB_LUT4 add_6520_8_lut (.I0(GND_net), .I1(n19538[5]), .I2(n545), .I3(n59614), 
            .O(n19254[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61574_4_lut (.I0(n75809), .I1(n76900), .I2(n45_adj_4729), 
            .I3(n75421), .O(n77409));   // verilog/motorControl.v(47[25:43])
    defparam i61574_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59982_3_lut (.I0(n77557), .I1(n535[20]), .I2(n41_adj_4727), 
            .I3(GND_net), .O(n75817));   // verilog/motorControl.v(47[25:43])
    defparam i59982_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6520_8 (.CI(n59614), .I0(n19538[5]), .I1(n545), .CO(n59615));
    SB_LUT4 add_6520_7_lut (.I0(GND_net), .I1(n19538[4]), .I2(n472), .I3(n59613), 
            .O(n19254[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_7 (.CI(n59613), .I0(n19538[4]), .I1(n472), .CO(n59614));
    SB_LUT4 i61576_4_lut (.I0(n75817), .I1(n77409), .I2(n45_adj_4729), 
            .I3(n75427), .O(n77411));   // verilog/motorControl.v(47[25:43])
    defparam i61576_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6520_6_lut (.I0(GND_net), .I1(n19538[3]), .I2(n399), .I3(n59612), 
            .O(n19254[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_6 (.CI(n59612), .I0(n19538[3]), .I1(n399), .CO(n59613));
    SB_LUT4 add_6520_5_lut (.I0(GND_net), .I1(n19538[2]), .I2(n326), .I3(n59611), 
            .O(n19254[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_5 (.CI(n59611), .I0(n19538[2]), .I1(n326), .CO(n59612));
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6520_4_lut (.I0(GND_net), .I1(n19538[1]), .I2(n253), .I3(n59610), 
            .O(n19254[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4798));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6520_4 (.CI(n59610), .I0(n19538[1]), .I1(n253), .CO(n59611));
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4799));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_3_lut (.I0(GND_net), .I1(n19538[0]), .I2(n180), .I3(n59609), 
            .O(n19254[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_3 (.CI(n59609), .I0(n19538[0]), .I1(n180), .CO(n59610));
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4800));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6520_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n19254[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6520_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6520_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n59609));
    SB_LUT4 add_6542_12_lut (.I0(GND_net), .I1(n19776[9]), .I2(n840_adj_4461), 
            .I3(n59608), .O(n19538[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6542_11_lut (.I0(GND_net), .I1(n19776[8]), .I2(n767_adj_4460), 
            .I3(n59607), .O(n19538[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4802));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4803));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\control_mode[5] ), .I1(\control_mode[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4804));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h4444;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4614));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_11 (.CI(n59607), .I0(n19776[8]), .I1(n767_adj_4460), 
            .CO(n59608));
    SB_LUT4 add_6542_10_lut (.I0(GND_net), .I1(n19776[7]), .I2(n694_adj_4459), 
            .I3(n59606), .O(n19538[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_10_lut (.I0(GND_net), .I1(n20130[7]), .I2(n700), 
            .I3(n58749), .O(n19972[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_9_lut (.I0(GND_net), .I1(n20130[6]), .I2(n627), .I3(n58748), 
            .O(n19972[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4613));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_10 (.CI(n59606), .I0(n19776[7]), .I1(n694_adj_4459), 
            .CO(n59607));
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6580_9 (.CI(n58748), .I0(n20130[6]), .I1(n627), .CO(n58749));
    SB_LUT4 add_6542_9_lut (.I0(GND_net), .I1(n19776[6]), .I2(n621_adj_4458), 
            .I3(n59605), .O(n19538[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_9 (.CI(n59605), .I0(n19776[6]), .I1(n621_adj_4458), 
            .CO(n59606));
    SB_LUT4 add_6542_8_lut (.I0(GND_net), .I1(n19776[5]), .I2(n548_adj_4457), 
            .I3(n59604), .O(n19538[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_8_lut (.I0(GND_net), .I1(n20130[5]), .I2(n554), .I3(n58747), 
            .O(n19972[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4612));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4806));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6580_8 (.CI(n58747), .I0(n20130[5]), .I1(n554), .CO(n58748));
    SB_CARRY add_6542_8 (.CI(n59604), .I0(n19776[5]), .I1(n548_adj_4457), 
            .CO(n59605));
    SB_LUT4 add_6580_7_lut (.I0(GND_net), .I1(n20130[4]), .I2(n481), .I3(n58746), 
            .O(n19972[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4807));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4808));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6580_7 (.CI(n58746), .I0(n20130[4]), .I1(n481), .CO(n58747));
    SB_LUT4 add_6542_7_lut (.I0(GND_net), .I1(n19776[4]), .I2(n475_adj_4456), 
            .I3(n59603), .O(n19538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4809));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6580_6_lut (.I0(GND_net), .I1(n20130[3]), .I2(n408), .I3(n58745), 
            .O(n19972[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6542_7 (.CI(n59603), .I0(n19776[4]), .I1(n475_adj_4456), 
            .CO(n59604));
    SB_LUT4 add_6542_6_lut (.I0(GND_net), .I1(n19776[3]), .I2(n402_adj_4455), 
            .I3(n59602), .O(n19538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(\control_mode[1] ), .I1(\control_mode[6] ), .I2(\control_mode[7] ), 
            .I3(n6_adj_4804), .O(n65754));
    defparam i4_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6580_6 (.CI(n58745), .I0(n20130[3]), .I1(n408), .CO(n58746));
    SB_CARRY add_6542_6 (.CI(n59602), .I0(n19776[3]), .I1(n402_adj_4455), 
            .CO(n59603));
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6580_5_lut (.I0(GND_net), .I1(n20130[2]), .I2(n335), .I3(n58744), 
            .O(n19972[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6542_5_lut (.I0(GND_net), .I1(n19776[2]), .I2(n329_adj_4454), 
            .I3(n59601), .O(n19538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_5 (.CI(n58744), .I0(n20130[2]), .I1(n335), .CO(n58745));
    SB_CARRY add_6542_5 (.CI(n59601), .I0(n19776[2]), .I1(n329_adj_4454), 
            .CO(n59602));
    SB_LUT4 add_6580_4_lut (.I0(GND_net), .I1(n20130[1]), .I2(n262), .I3(n58743), 
            .O(n19972[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6542_4_lut (.I0(GND_net), .I1(n19776[1]), .I2(n256_adj_4453), 
            .I3(n59600), .O(n19538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_4 (.CI(n59600), .I0(n19776[1]), .I1(n256_adj_4453), 
            .CO(n59601));
    SB_CARRY add_6580_4 (.CI(n58743), .I0(n20130[1]), .I1(n262), .CO(n58744));
    SB_LUT4 add_6542_3_lut (.I0(GND_net), .I1(n19776[0]), .I2(n183_adj_4452), 
            .I3(n59599), .O(n19538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6580_3_lut (.I0(GND_net), .I1(n20130[0]), .I2(n189), .I3(n58742), 
            .O(n19972[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6542_3 (.CI(n59599), .I0(n19776[0]), .I1(n183_adj_4452), 
            .CO(n59600));
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4611));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6542_2_lut (.I0(GND_net), .I1(n41_adj_4450), .I2(n110), 
            .I3(GND_net), .O(n19538[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6542_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_3 (.CI(n58742), .I0(n20130[0]), .I1(n189), .CO(n58743));
    SB_LUT4 add_6580_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19972[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6580_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6542_2 (.CI(GND_net), .I0(n41_adj_4450), .I1(n110), .CO(n59599));
    SB_LUT4 add_6614_7_lut (.I0(GND_net), .I1(n68674), .I2(n490), .I3(n59598), 
            .O(n20287[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6580_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n58742));
    SB_LUT4 add_6614_6_lut (.I0(GND_net), .I1(n20370[3]), .I2(n417), .I3(n59597), 
            .O(n20287[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_6 (.CI(n59597), .I0(n20370[3]), .I1(n417), .CO(n59598));
    SB_LUT4 add_6614_5_lut (.I0(GND_net), .I1(n20370[2]), .I2(n344_adj_4443), 
            .I3(n59596), .O(n20287[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_20_lut (.I0(GND_net), .I1(n15963[17]), .I2(GND_net), 
            .I3(n58741), .O(n15204[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_5 (.CI(n59596), .I0(n20370[2]), .I1(n344_adj_4443), 
            .CO(n59597));
    SB_LUT4 add_6614_4_lut (.I0(GND_net), .I1(n20370[1]), .I2(n271), .I3(n59595), 
            .O(n20287[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_4 (.CI(n59595), .I0(n20370[1]), .I1(n271), .CO(n59596));
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6614_3_lut (.I0(GND_net), .I1(n20370[0]), .I2(n198), .I3(n59594), 
            .O(n20287[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_19_lut (.I0(GND_net), .I1(n15963[16]), .I2(GND_net), 
            .I3(n58740), .O(n15204[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6289_19 (.CI(n58740), .I0(n15963[16]), .I1(GND_net), 
            .CO(n58741));
    SB_CARRY add_6614_3 (.CI(n59594), .I0(n20370[0]), .I1(n198), .CO(n59595));
    SB_LUT4 add_6614_2_lut (.I0(GND_net), .I1(n56_c), .I2(n125), .I3(GND_net), 
            .O(n20287[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6614_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6614_2 (.CI(GND_net), .I0(n56_c), .I1(n125), .CO(n59594));
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4818));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_18_lut (.I0(GND_net), .I1(n15963[15]), .I2(GND_net), 
            .I3(n58739), .O(n15204[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_18 (.CI(n58739), .I0(n15963[15]), .I1(GND_net), 
            .CO(n58740));
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4997[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6289_17_lut (.I0(GND_net), .I1(n15963[14]), .I2(GND_net), 
            .I3(n58738), .O(n15204[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4821));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6289_17 (.CI(n58738), .I0(n15963[14]), .I1(GND_net), 
            .CO(n58739));
    SB_LUT4 LessThan_9_i43_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4822));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4823));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6289_16_lut (.I0(GND_net), .I1(n15963[13]), .I2(n1108), 
            .I3(n58737), .O(n15204[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4824));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6289_16 (.CI(n58737), .I0(n15963[13]), .I1(n1108), .CO(n58738));
    SB_LUT4 add_6289_15_lut (.I0(GND_net), .I1(n15963[12]), .I2(n1035), 
            .I3(n58736), .O(n15204[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n58195), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_15 (.CI(n58736), .I0(n15963[12]), .I1(n1035), .CO(n58737));
    SB_LUT4 add_6289_14_lut (.I0(GND_net), .I1(n15963[11]), .I2(n962), 
            .I3(n58735), .O(n15204[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_7 (.CI(n58195), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n58196));
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n58194), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n58382), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_14 (.CI(n58735), .I0(n15963[11]), .I1(n962), .CO(n58736));
    SB_LUT4 add_6289_13_lut (.I0(GND_net), .I1(n15963[10]), .I2(n889), 
            .I3(n58734), .O(n15204[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n58171), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n58381), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4827));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_4828));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_9_i8_3_lut (.I0(n6_adj_4829), .I1(setpoint[4]), .I2(n9), 
            .I3(GND_net), .O(n8_adj_4831));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4832));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61608_4_lut (.I0(n8_adj_4831), .I1(n4_adj_4828), .I2(n9), 
            .I3(n75597), .O(n77443));   // verilog/motorControl.v(45[16:33])
    defparam i61608_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6289_13 (.CI(n58734), .I0(n15963[10]), .I1(n889), .CO(n58735));
    SB_LUT4 add_6289_12_lut (.I0(GND_net), .I1(n15963[9]), .I2(n816), 
            .I3(n58733), .O(n15204[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_12 (.CI(n58733), .I0(n15963[9]), .I1(n816), .CO(n58734));
    SB_CARRY unary_minus_33_add_3_24 (.CI(n58381), .I0(GND_net), .I1(n1[22]), 
            .CO(n58382));
    SB_LUT4 i61609_3_lut (.I0(n77443), .I1(setpoint[5]), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n77444));   // verilog/motorControl.v(45[16:33])
    defparam i61609_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61489_3_lut (.I0(n77444), .I1(setpoint[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n77324));   // verilog/motorControl.v(45[16:33])
    defparam i61489_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6289_11_lut (.I0(GND_net), .I1(n15963[8]), .I2(n743), 
            .I3(n58732), .O(n15204[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n58380), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_11 (.CI(n58732), .I0(n15963[8]), .I1(n743), .CO(n58733));
    SB_LUT4 add_6289_10_lut (.I0(GND_net), .I1(n15963[7]), .I2(n670), 
            .I3(n58731), .O(n15204[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59968_3_lut (.I0(n77324), .I1(setpoint[7]), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(45[16:33])
    defparam i59968_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_6289_10 (.CI(n58731), .I0(n15963[7]), .I1(n670), .CO(n58732));
    SB_CARRY add_16_6 (.CI(n58194), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n58195));
    SB_LUT4 add_6289_9_lut (.I0(GND_net), .I1(n15963[6]), .I2(n597), .I3(n58730), 
            .O(n15204[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_23 (.CI(n58380), .I0(GND_net), .I1(n1[21]), 
            .CO(n58381));
    SB_CARRY add_6289_9 (.CI(n58730), .I0(n15963[6]), .I1(n597), .CO(n58731));
    SB_LUT4 add_6289_8_lut (.I0(GND_net), .I1(n15963[5]), .I2(n524), .I3(n58729), 
            .O(n15204[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n58379), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n58193), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_8 (.CI(n58729), .I0(n15963[5]), .I1(n524), .CO(n58730));
    SB_LUT4 add_6289_7_lut (.I0(GND_net), .I1(n15963[4]), .I2(n451), .I3(n58728), 
            .O(n15204[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n58379), .I0(GND_net), .I1(n1[20]), 
            .CO(n58380));
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n58378), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n58378), .I0(GND_net), .I1(n1[19]), 
            .CO(n58379));
    SB_CARRY add_6289_7 (.CI(n58728), .I0(n15963[4]), .I1(n451), .CO(n58729));
    SB_LUT4 LessThan_9_i20_3_lut (.I0(n34707), .I1(setpoint[9]), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6289_6_lut (.I0(GND_net), .I1(n15963[3]), .I2(n378), .I3(n58727), 
            .O(n15204[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_6 (.CI(n58727), .I0(n15963[3]), .I1(n378), .CO(n58728));
    SB_LUT4 add_6289_5_lut (.I0(GND_net), .I1(n15963[2]), .I2(n305_adj_4436), 
            .I3(n58726), .O(n15204[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_5 (.CI(n58726), .I0(n15963[2]), .I1(n305_adj_4436), 
            .CO(n58727));
    SB_LUT4 add_6289_4_lut (.I0(GND_net), .I1(n15963[1]), .I2(n232), .I3(n58725), 
            .O(n15204[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_4 (.CI(n58725), .I0(n15963[1]), .I1(n232), .CO(n58726));
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n58377), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_20 (.CI(n58377), .I0(GND_net), .I1(n1[18]), 
            .CO(n58378));
    SB_LUT4 add_6289_3_lut (.I0(GND_net), .I1(n15963[0]), .I2(n159), .I3(n58724), 
            .O(n15204[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_3 (.CI(n58724), .I0(n15963[0]), .I1(n159), .CO(n58725));
    SB_LUT4 add_6289_2_lut (.I0(GND_net), .I1(n17_adj_4435), .I2(n86), 
            .I3(GND_net), .O(n15204[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_2 (.CI(GND_net), .I0(n17_adj_4435), .I1(n86), .CO(n58724));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n58376), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n58376), .I0(GND_net), .I1(n1[17]), 
            .CO(n58377));
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4835));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n58375), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n58375), .I0(GND_net), .I1(n1[16]), 
            .CO(n58376));
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n58374), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4836));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i31_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4837));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i35_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4838));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4839));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59737_4_lut (.I0(n29_adj_4836), .I1(n27_adj_4835), .I2(n25), 
            .I3(n23_adj_4839), .O(n75572));
    defparam i59737_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59723_4_lut (.I0(n35_adj_4838), .I1(n33), .I2(n31_adj_4837), 
            .I3(n75572), .O(n75558));
    defparam i59723_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_33_add_3_17 (.CI(n58374), .I0(GND_net), .I1(n1[15]), 
            .CO(n58375));
    SB_LUT4 LessThan_9_i30_3_lut (.I0(n28), .I1(setpoint[16]), .I2(n33), 
            .I3(GND_net), .O(n30_adj_4842));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n58373), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_16 (.CI(n58373), .I0(GND_net), .I1(n1[14]), 
            .CO(n58374));
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n58372), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_15 (.CI(n58372), .I0(GND_net), .I1(n1[13]), 
            .CO(n58373));
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n58371), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_14 (.CI(n58371), .I0(GND_net), .I1(n1[12]), 
            .CO(n58372));
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n58370), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n58370), .I0(GND_net), .I1(n1[11]), 
            .CO(n58371));
    SB_CARRY add_16_5 (.CI(n58193), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n58194));
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n58369), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_12 (.CI(n58369), .I0(GND_net), .I1(n1[10]), 
            .CO(n58370));
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n58368), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_11 (.CI(n58368), .I0(GND_net), .I1(n1[9]), 
            .CO(n58369));
    SB_LUT4 add_6326_19_lut (.I0(GND_net), .I1(n16646[16]), .I2(GND_net), 
            .I3(n58704), .O(n15963[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_18_lut (.I0(GND_net), .I1(n16646[15]), .I2(GND_net), 
            .I3(n58703), .O(n15963[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_18 (.CI(n58703), .I0(n16646[15]), .I1(GND_net), 
            .CO(n58704));
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n58367), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_17_lut (.I0(GND_net), .I1(n16646[14]), .I2(GND_net), 
            .I3(n58702), .O(n15963[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_10 (.CI(n58367), .I0(GND_net), .I1(n1[8]), 
            .CO(n58368));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n58366), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_17 (.CI(n58702), .I0(n16646[14]), .I1(GND_net), 
            .CO(n58703));
    SB_CARRY unary_minus_33_add_3_9 (.CI(n58366), .I0(GND_net), .I1(n1[7]), 
            .CO(n58367));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n58192), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_16_lut (.I0(GND_net), .I1(n16646[13]), .I2(n1111), 
            .I3(n58701), .O(n15963[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_16 (.CI(n58701), .I0(n16646[13]), .I1(n1111), .CO(n58702));
    SB_LUT4 add_6326_15_lut (.I0(GND_net), .I1(n16646[12]), .I2(n1038), 
            .I3(n58700), .O(n15963[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n58365), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_15 (.CI(n58700), .I0(n16646[12]), .I1(n1038), .CO(n58701));
    SB_LUT4 add_6326_14_lut (.I0(GND_net), .I1(n16646[11]), .I2(n965), 
            .I3(n58699), .O(n15963[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_14 (.CI(n58699), .I0(n16646[11]), .I1(n965), .CO(n58700));
    SB_CARRY unary_minus_33_add_3_8 (.CI(n58365), .I0(GND_net), .I1(n1[6]), 
            .CO(n58366));
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n58364), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n58364), .I0(GND_net), .I1(n1[5]), 
            .CO(n58365));
    SB_LUT4 add_6326_13_lut (.I0(GND_net), .I1(n16646[10]), .I2(n892), 
            .I3(n58698), .O(n15963[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_13 (.CI(n58698), .I0(n16646[10]), .I1(n892), .CO(n58699));
    SB_CARRY add_16_4 (.CI(n58192), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n58193));
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n58191), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_6 (.CI(n58171), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n58172));
    SB_CARRY sub_15_add_2_5 (.CI(n58170), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n58171));
    SB_CARRY sub_15_add_2_4 (.CI(n58169), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n58170));
    SB_LUT4 add_6326_12_lut (.I0(GND_net), .I1(n16646[9]), .I2(n819), 
            .I3(n58697), .O(n15963[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n58363), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_3 (.CI(n58168), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n58169));
    SB_CARRY add_6326_12 (.CI(n58697), .I0(n16646[9]), .I1(n819), .CO(n58698));
    SB_LUT4 add_6326_11_lut (.I0(GND_net), .I1(n16646[8]), .I2(n746), 
            .I3(n58696), .O(n15963[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_3 (.CI(n58191), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n58192));
    SB_CARRY add_6326_11 (.CI(n58696), .I0(n16646[8]), .I1(n746), .CO(n58697));
    SB_LUT4 LessThan_9_i34_3_lut (.I0(n26_adj_4843), .I1(setpoint[18]), 
            .I2(n37), .I3(GND_net), .O(n34));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6326_10_lut (.I0(GND_net), .I1(n16646[7]), .I2(n673), 
            .I3(n58695), .O(n15963[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_6 (.CI(n58363), .I0(GND_net), .I1(n1[4]), 
            .CO(n58364));
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n58362), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_10 (.CI(n58695), .I0(n16646[7]), .I1(n673), .CO(n58696));
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n58191));
    SB_LUT4 i61610_4_lut (.I0(n34), .I1(n24_adj_4845), .I2(n37), .I3(n75556), 
            .O(n77445));   // verilog/motorControl.v(45[16:33])
    defparam i61610_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6326_9_lut (.I0(GND_net), .I1(n16646[6]), .I2(n600), .I3(n58694), 
            .O(n15963[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61611_3_lut (.I0(n77445), .I1(setpoint[19]), .I2(n39_adj_4824), 
            .I3(GND_net), .O(n77446));   // verilog/motorControl.v(45[16:33])
    defparam i61611_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6326_9 (.CI(n58694), .I0(n16646[6]), .I1(n600), .CO(n58695));
    SB_LUT4 add_6326_8_lut (.I0(GND_net), .I1(n16646[5]), .I2(n527), .I3(n58693), 
            .O(n15963[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_5 (.CI(n58362), .I0(GND_net), .I1(n1[3]), 
            .CO(n58363));
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n58190), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_8 (.CI(n58693), .I0(n16646[5]), .I1(n527), .CO(n58694));
    SB_LUT4 add_6326_7_lut (.I0(GND_net), .I1(n16646[4]), .I2(n454), .I3(n58692), 
            .O(n15963[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_7 (.CI(n58692), .I0(n16646[4]), .I1(n454), .CO(n58693));
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n58361), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_4 (.CI(n58361), .I0(GND_net), .I1(n1[2]), 
            .CO(n58362));
    SB_LUT4 i61487_3_lut (.I0(n77446), .I1(setpoint[20]), .I2(n41), .I3(GND_net), 
            .O(n77322));   // verilog/motorControl.v(45[16:33])
    defparam i61487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n58360), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6326_6_lut (.I0(GND_net), .I1(n16646[3]), .I2(n381_adj_4832), 
            .I3(n58691), .O(n15963[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6326_6 (.CI(n58691), .I0(n16646[3]), .I1(n381_adj_4832), 
            .CO(n58692));
    SB_LUT4 add_6326_5_lut (.I0(GND_net), .I1(n16646[2]), .I2(n308_adj_4827), 
            .I3(n58690), .O(n15963[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_3 (.CI(n58360), .I0(GND_net), .I1(n1[1]), 
            .CO(n58361));
    SB_CARRY add_6326_5 (.CI(n58690), .I0(n16646[2]), .I1(n308_adj_4827), 
            .CO(n58691));
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61342_4_lut (.I0(n41), .I1(n39_adj_4824), .I2(n37), .I3(n75558), 
            .O(n77177));
    defparam i61342_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n58189), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61508_4_lut (.I0(n30_adj_4842), .I1(n22_adj_1), .I2(n33), 
            .I3(n75566), .O(n77343));   // verilog/motorControl.v(45[16:33])
    defparam i61508_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_6326_4_lut (.I0(GND_net), .I1(n16646[1]), .I2(n235_adj_4823), 
            .I3(n58689), .O(n15963[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59972_3_lut (.I0(n77322), .I1(setpoint[21]), .I2(n43_adj_4822), 
            .I3(GND_net), .O(n75807));   // verilog/motorControl.v(45[16:33])
    defparam i59972_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6326_4 (.CI(n58689), .I0(n16646[1]), .I1(n235_adj_4823), 
            .CO(n58690));
    SB_LUT4 add_6326_3_lut (.I0(GND_net), .I1(n16646[0]), .I2(n162_adj_4821), 
            .I3(n58688), .O(n15963[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n58360));
    SB_CARRY add_6326_3 (.CI(n58688), .I0(n16646[0]), .I1(n162_adj_4821), 
            .CO(n58689));
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_4997[23]), 
            .I3(n58359), .O(n47_adj_4849)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6326_2_lut (.I0(GND_net), .I1(n20_adj_4819), .I2(n89_adj_4818), 
            .I3(GND_net), .O(n15963[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6326_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61652_4_lut (.I0(n75807), .I1(n77343), .I2(n43_adj_4822), 
            .I3(n77177), .O(n77487));   // verilog/motorControl.v(45[16:33])
    defparam i61652_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6326_2 (.CI(GND_net), .I0(n20_adj_4819), .I1(n89_adj_4818), 
            .CO(n58688));
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[22]), 
            .I3(n58358), .O(n48[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61653_3_lut (.I0(n77487), .I1(setpoint[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n77488));   // verilog/motorControl.v(45[16:33])
    defparam i61653_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61383_3_lut (.I0(n77488), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i61383_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n58358), .I0(GND_net), .I1(n1_adj_4997[22]), 
            .CO(n58359));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[21]), 
            .I3(n58357), .O(n48[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_24 (.CI(n58189), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n58190));
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n58188), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n58168));
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4851));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n58357), .I0(GND_net), .I1(n1_adj_4997[21]), 
            .CO(n58358));
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4852));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[20]), 
            .I3(n58356), .O(n48[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_23 (.CI(n58188), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n58189));
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4853));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4854));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_27_add_3_22 (.CI(n58356), .I0(GND_net), .I1(n1_adj_4997[20]), 
            .CO(n58357));
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4855));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4856));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i7_2_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4857));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[19]), 
            .I3(n58355), .O(n486)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_21 (.CI(n58355), .I0(GND_net), .I1(n1_adj_4997[19]), 
            .CO(n58356));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[18]), 
            .I3(n58354), .O(n48[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4859));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i5_2_lut (.I0(PWMLimit[2]), .I1(n455[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4860));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_27_add_3_20 (.CI(n58354), .I0(GND_net), .I1(n1_adj_4997[18]), 
            .CO(n58355));
    SB_LUT4 i59305_4_lut (.I0(n11_adj_4859), .I1(n35808), .I2(n7_adj_4857), 
            .I3(n5_adj_4860), .O(n75140));
    defparam i59305_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[17]), 
            .I3(n58353), .O(n48[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n58187), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n475), .I1(n455[8]), .I2(n17_adj_4856), 
            .I3(GND_net), .O(n8_adj_4861));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6596_9_lut (.I0(GND_net), .I1(n20254[6]), .I2(n630_adj_4810), 
            .I3(n58669), .O(n20130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6596_8_lut (.I0(GND_net), .I1(n20254[5]), .I2(n557_adj_4809), 
            .I3(n58668), .O(n20130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_8 (.CI(n58668), .I0(n20254[5]), .I1(n557_adj_4809), 
            .CO(n58669));
    SB_LUT4 add_6596_7_lut (.I0(GND_net), .I1(n20254[4]), .I2(n484_adj_4808), 
            .I3(n58667), .O(n20130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_7 (.CI(n58667), .I0(n20254[4]), .I1(n484_adj_4808), 
            .CO(n58668));
    SB_LUT4 add_6596_6_lut (.I0(GND_net), .I1(n20254[3]), .I2(n411_adj_4807), 
            .I3(n58666), .O(n20130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i6_3_lut (.I0(n455[2]), .I1(n455[3]), .I2(n7_adj_4857), 
            .I3(GND_net), .O(n6_adj_4862));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6596_6 (.CI(n58666), .I0(n20254[3]), .I1(n411_adj_4807), 
            .CO(n58667));
    SB_LUT4 add_6596_5_lut (.I0(GND_net), .I1(n20254[2]), .I2(n338_adj_4806), 
            .I3(n58665), .O(n20130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n58353), .I0(GND_net), .I1(n1_adj_4997[17]), 
            .CO(n58354));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[16]), 
            .I3(n58352), .O(n48[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_5 (.CI(n58665), .I0(n20254[2]), .I1(n338_adj_4806), 
            .CO(n58666));
    SB_CARRY unary_minus_27_add_3_18 (.CI(n58352), .I0(GND_net), .I1(n1_adj_4997[16]), 
            .CO(n58353));
    SB_LUT4 add_6596_4_lut (.I0(GND_net), .I1(n20254[1]), .I2(n265_adj_4803), 
            .I3(n58664), .O(n20130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_4 (.CI(n58664), .I0(n20254[1]), .I1(n265_adj_4803), 
            .CO(n58665));
    SB_LUT4 add_6596_3_lut (.I0(GND_net), .I1(n20254[0]), .I2(n192_adj_4802), 
            .I3(n58663), .O(n20130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n8_adj_4861), .I1(n455[9]), .I2(n19_adj_4855), 
            .I3(GND_net), .O(n16_adj_4863));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4865));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_CARRY add_6596_3 (.CI(n58663), .I0(n20254[0]), .I1(n192_adj_4802), 
            .CO(n58664));
    SB_LUT4 add_6596_2_lut (.I0(GND_net), .I1(n50_adj_4800), .I2(n119_adj_4799), 
            .I3(GND_net), .O(n20130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6596_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6596_2 (.CI(GND_net), .I0(n50_adj_4800), .I1(n119_adj_4799), 
            .CO(n58663));
    SB_LUT4 add_6361_18_lut (.I0(GND_net), .I1(n17257[15]), .I2(GND_net), 
            .I3(n58662), .O(n16646[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_17_lut (.I0(GND_net), .I1(n17257[14]), .I2(GND_net), 
            .I3(n58661), .O(n16646[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_17 (.CI(n58661), .I0(n17257[14]), .I1(GND_net), 
            .CO(n58662));
    SB_LUT4 add_6361_16_lut (.I0(GND_net), .I1(n17257[13]), .I2(n1114_adj_4798), 
            .I3(n58660), .O(n16646[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_16 (.CI(n58660), .I0(n17257[13]), .I1(n1114_adj_4798), 
            .CO(n58661));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[15]), 
            .I3(n58351), .O(n48[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_17 (.CI(n58351), .I0(GND_net), .I1(n1_adj_4997[15]), 
            .CO(n58352));
    SB_CARRY sub_15_add_2_22 (.CI(n58187), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n58188));
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n58186), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[14]), 
            .I3(n58350), .O(n48[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n58350), .I0(GND_net), .I1(n1_adj_4997[14]), 
            .CO(n58351));
    SB_LUT4 i61199_3_lut (.I0(n4_adj_4865), .I1(n455[5]), .I2(n11_adj_4859), 
            .I3(GND_net), .O(n77034));   // verilog/motorControl.v(63[16:31])
    defparam i61199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6361_15_lut (.I0(GND_net), .I1(n17257[12]), .I2(n1041_adj_4795), 
            .I3(n58659), .O(n16646[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_15 (.CI(n58659), .I0(n17257[12]), .I1(n1041_adj_4795), 
            .CO(n58660));
    SB_LUT4 add_6361_14_lut (.I0(GND_net), .I1(n17257[11]), .I2(n968_adj_4794), 
            .I3(n58658), .O(n16646[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_14 (.CI(n58658), .I0(n17257[11]), .I1(n968_adj_4794), 
            .CO(n58659));
    SB_LUT4 add_6361_13_lut (.I0(GND_net), .I1(n17257[10]), .I2(n895_adj_4793), 
            .I3(n58657), .O(n16646[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_13 (.CI(n58657), .I0(n17257[10]), .I1(n895_adj_4793), 
            .CO(n58658));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[13]), 
            .I3(n58349), .O(n48[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_12_lut (.I0(GND_net), .I1(n17257[9]), .I2(n822_adj_4791), 
            .I3(n58656), .O(n16646[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_15 (.CI(n58349), .I0(GND_net), .I1(n1_adj_4997[13]), 
            .CO(n58350));
    SB_CARRY add_6361_12 (.CI(n58656), .I0(n17257[9]), .I1(n822_adj_4791), 
            .CO(n58657));
    SB_CARRY sub_15_add_2_21 (.CI(n58186), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n58187));
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n58185), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[12]), 
            .I3(n58348), .O(n48[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61200_3_lut (.I0(n77034), .I1(n455[6]), .I2(n13_adj_4853), 
            .I3(GND_net), .O(n77035));   // verilog/motorControl.v(63[16:31])
    defparam i61200_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n58348), .I0(GND_net), .I1(n1_adj_4997[12]), 
            .CO(n58349));
    SB_LUT4 i59301_4_lut (.I0(n17_adj_4856), .I1(n15_adj_4854), .I2(n13_adj_4853), 
            .I3(n75140), .O(n75136));
    defparam i59301_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[11]), 
            .I3(n58347), .O(n48[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_11_lut (.I0(GND_net), .I1(n17257[8]), .I2(n749_adj_4788), 
            .I3(n58655), .O(n16646[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_11 (.CI(n58655), .I0(n17257[8]), .I1(n749_adj_4788), 
            .CO(n58656));
    SB_LUT4 add_6361_10_lut (.I0(GND_net), .I1(n17257[7]), .I2(n676_adj_4787), 
            .I3(n58654), .O(n16646[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_10 (.CI(n58654), .I0(n17257[7]), .I1(n676_adj_4787), 
            .CO(n58655));
    SB_LUT4 add_6361_9_lut (.I0(GND_net), .I1(n17257[6]), .I2(n603_adj_4786), 
            .I3(n58653), .O(n16646[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_9 (.CI(n58653), .I0(n17257[6]), .I1(n603_adj_4786), 
            .CO(n58654));
    SB_CARRY unary_minus_27_add_3_13 (.CI(n58347), .I0(GND_net), .I1(n1_adj_4997[11]), 
            .CO(n58348));
    SB_LUT4 add_6361_8_lut (.I0(GND_net), .I1(n17257[5]), .I2(n530_adj_4785), 
            .I3(n58652), .O(n16646[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_8 (.CI(n58652), .I0(n17257[5]), .I1(n530_adj_4785), 
            .CO(n58653));
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[10]), 
            .I3(n58346), .O(n48[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6361_7_lut (.I0(GND_net), .I1(n17257[4]), .I2(n457_adj_4783), 
            .I3(n58651), .O(n16646[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61496_4_lut (.I0(n16_adj_4863), .I1(n6_adj_4862), .I2(n19_adj_4855), 
            .I3(n75134), .O(n77331));   // verilog/motorControl.v(63[16:31])
    defparam i61496_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6361_7 (.CI(n58651), .I0(n17257[4]), .I1(n457_adj_4783), 
            .CO(n58652));
    SB_LUT4 add_6361_6_lut (.I0(GND_net), .I1(n17257[3]), .I2(n384_adj_4782), 
            .I3(n58650), .O(n16646[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_6 (.CI(n58650), .I0(n17257[3]), .I1(n384_adj_4782), 
            .CO(n58651));
    SB_LUT4 add_6361_5_lut (.I0(GND_net), .I1(n17257[2]), .I2(n311_adj_4779), 
            .I3(n58649), .O(n16646[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_5 (.CI(n58649), .I0(n17257[2]), .I1(n311_adj_4779), 
            .CO(n58650));
    SB_CARRY sub_15_add_2_20 (.CI(n58185), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n58186));
    SB_LUT4 add_6361_4_lut (.I0(GND_net), .I1(n17257[1]), .I2(n238_adj_4778), 
            .I3(n58648), .O(n16646[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_4 (.CI(n58648), .I0(n17257[1]), .I1(n238_adj_4778), 
            .CO(n58649));
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n58184), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n58346), .I0(GND_net), .I1(n1_adj_4997[10]), 
            .CO(n58347));
    SB_LUT4 add_6361_3_lut (.I0(GND_net), .I1(n17257[0]), .I2(n165_adj_4776), 
            .I3(n58647), .O(n16646[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[9]), 
            .I3(n58345), .O(n48[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6361_3 (.CI(n58647), .I0(n17257[0]), .I1(n165_adj_4776), 
            .CO(n58648));
    SB_LUT4 i60024_3_lut (.I0(n77035), .I1(n455[7]), .I2(n15_adj_4854), 
            .I3(GND_net), .O(n75859));   // verilog/motorControl.v(63[16:31])
    defparam i60024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6361_2_lut (.I0(GND_net), .I1(n23_adj_4773), .I2(n92_adj_4772), 
            .I3(GND_net), .O(n16646[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6361_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_11 (.CI(n58345), .I0(GND_net), .I1(n1_adj_4997[9]), 
            .CO(n58346));
    SB_CARRY add_6361_2 (.CI(GND_net), .I0(n23_adj_4773), .I1(n92_adj_4772), 
            .CO(n58647));
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[8]), 
            .I3(n58344), .O(n48[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61733_4_lut (.I0(n75859), .I1(n77331), .I2(n19_adj_4855), 
            .I3(n75136), .O(n77568));   // verilog/motorControl.v(63[16:31])
    defparam i61733_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61734_3_lut (.I0(n77568), .I1(n455[10]), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n77569));   // verilog/motorControl.v(63[16:31])
    defparam i61734_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_15_add_2_19 (.CI(n58184), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n58185));
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n58183), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n58344), .I0(GND_net), .I1(n1_adj_4997[8]), 
            .CO(n58345));
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[7]), 
            .I3(n58343), .O(n48[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n58343), .I0(GND_net), .I1(n1_adj_4997[7]), 
            .CO(n58344));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[6]), 
            .I3(n58342), .O(n48[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n58342), .I0(GND_net), .I1(n1_adj_4997[6]), 
            .CO(n58343));
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[5]), 
            .I3(n58341), .O(n48[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n58341), .I0(GND_net), .I1(n1_adj_4997[5]), 
            .CO(n58342));
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[4]), 
            .I3(n58340), .O(n48[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n58183), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n58184));
    SB_CARRY unary_minus_27_add_3_6 (.CI(n58340), .I0(GND_net), .I1(n1_adj_4997[4]), 
            .CO(n58341));
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[3]), 
            .I3(n58339), .O(n48[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61684_3_lut (.I0(n77569), .I1(n455[11]), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(63[16:31])
    defparam i61684_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n58339), .I0(GND_net), .I1(n1_adj_4997[3]), 
            .CO(n58340));
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[2]), 
            .I3(n58338), .O(n48[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_4 (.CI(n58338), .I0(GND_net), .I1(n1_adj_4997[2]), 
            .CO(n58339));
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4997[1]), 
            .I3(n58337), .O(n48[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n58337), .I0(GND_net), .I1(n1_adj_4997[1]), 
            .CO(n58338));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n45170), .I1(GND_net), .I2(n1_adj_4997[0]), 
            .I3(VCC_net), .O(n74481)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n58182), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4997[0]), 
            .CO(n58337));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[23]), 
            .I3(n58336), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[22]), 
            .I3(n58335), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n58335), .I0(GND_net), .I1(n1_adj_4996[22]), 
            .CO(n58336));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[21]), 
            .I3(n58334), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n58182), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n58183));
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n58181), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n58334), .I0(GND_net), .I1(n1_adj_4996[21]), 
            .CO(n58335));
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4868));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n460), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4869));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4870));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[20]), 
            .I3(n58333), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n58333), .I0(GND_net), .I1(n1_adj_4996[20]), 
            .CO(n58334));
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4871));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[19]), 
            .I3(n58332), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n58332), .I0(GND_net), .I1(n1_adj_4996[19]), 
            .CO(n58333));
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4872));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6394_17_lut (.I0(GND_net), .I1(n17800[14]), .I2(GND_net), 
            .I3(n58629), .O(n17257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6394_16_lut (.I0(GND_net), .I1(n17800[13]), .I2(n1117_adj_4638), 
            .I3(n58628), .O(n17257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4873));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59291_4_lut (.I0(n33_adj_4872), .I1(n31_adj_4871), .I2(n29_adj_4870), 
            .I3(n27_adj_4873), .O(n75126));
    defparam i59291_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n455[15]), .I1(n460), .I2(n39_adj_4869), 
            .I3(GND_net), .O(n30_adj_4874));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i28_3_lut (.I0(n455[13]), .I1(n455[14]), .I2(n29_adj_4870), 
            .I3(GND_net), .O(n28_adj_4875));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6394_16 (.CI(n58628), .I0(n17800[13]), .I1(n1117_adj_4638), 
            .CO(n58629));
    SB_LUT4 add_6394_15_lut (.I0(GND_net), .I1(n17800[12]), .I2(n1044_adj_4637), 
            .I3(n58627), .O(n17257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i38_3_lut (.I0(n30_adj_4874), .I1(n455[20]), .I2(n41_adj_4868), 
            .I3(GND_net), .O(n38_adj_4876));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6394_15 (.CI(n58627), .I0(n17800[12]), .I1(n1044_adj_4637), 
            .CO(n58628));
    SB_LUT4 add_6394_14_lut (.I0(GND_net), .I1(n17800[11]), .I2(n971_adj_4636), 
            .I3(n58626), .O(n17257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_14 (.CI(n58626), .I0(n17800[11]), .I1(n971_adj_4636), 
            .CO(n58627));
    SB_LUT4 add_6394_13_lut (.I0(GND_net), .I1(n17800[10]), .I2(n898_adj_4635), 
            .I3(n58625), .O(n17257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_13 (.CI(n58625), .I0(n17800[10]), .I1(n898_adj_4635), 
            .CO(n58626));
    SB_LUT4 add_6394_12_lut (.I0(GND_net), .I1(n17800[9]), .I2(n825_adj_4634), 
            .I3(n58624), .O(n17257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61195_3_lut (.I0(n36173), .I1(n455[16]), .I2(n33_adj_4872), 
            .I3(GND_net), .O(n77030));   // verilog/motorControl.v(63[16:31])
    defparam i61195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61196_3_lut (.I0(n77030), .I1(n455[17]), .I2(n35_adj_4852), 
            .I3(GND_net), .O(n77031));   // verilog/motorControl.v(63[16:31])
    defparam i61196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59285_4_lut (.I0(n39_adj_4869), .I1(n37_adj_4851), .I2(n35_adj_4852), 
            .I3(n75126), .O(n75120));
    defparam i59285_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6394_12 (.CI(n58624), .I0(n17800[9]), .I1(n825_adj_4634), 
            .CO(n58625));
    SB_LUT4 add_6394_11_lut (.I0(GND_net), .I1(n17800[8]), .I2(n752_adj_4633), 
            .I3(n58623), .O(n17257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_11 (.CI(n58623), .I0(n17800[8]), .I1(n752_adj_4633), 
            .CO(n58624));
    SB_LUT4 add_6394_10_lut (.I0(GND_net), .I1(n17800[7]), .I2(n679_adj_4632), 
            .I3(n58622), .O(n17257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61622_4_lut (.I0(n38_adj_4876), .I1(n28_adj_4875), .I2(n41_adj_4868), 
            .I3(n75118), .O(n77457));   // verilog/motorControl.v(63[16:31])
    defparam i61622_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6394_10 (.CI(n58622), .I0(n17800[7]), .I1(n679_adj_4632), 
            .CO(n58623));
    SB_LUT4 add_6394_9_lut (.I0(GND_net), .I1(n17800[6]), .I2(n606_adj_4631), 
            .I3(n58621), .O(n17257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_9 (.CI(n58621), .I0(n17800[6]), .I1(n606_adj_4631), 
            .CO(n58622));
    SB_LUT4 i60026_3_lut (.I0(n77031), .I1(n455[18]), .I2(n37_adj_4851), 
            .I3(GND_net), .O(n75861));   // verilog/motorControl.v(63[16:31])
    defparam i60026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61762_4_lut (.I0(n75861), .I1(n77457), .I2(n41_adj_4868), 
            .I3(n75120), .O(n77597));   // verilog/motorControl.v(63[16:31])
    defparam i61762_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_6394_8_lut (.I0(GND_net), .I1(n17800[5]), .I2(n533_adj_4630), 
            .I3(n58620), .O(n17257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_8 (.CI(n58620), .I0(n17800[5]), .I1(n533_adj_4630), 
            .CO(n58621));
    SB_LUT4 i61763_3_lut (.I0(n77597), .I1(n455[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n77598));   // verilog/motorControl.v(63[16:31])
    defparam i61763_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61713_3_lut (.I0(n77598), .I1(n455[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n77548));   // verilog/motorControl.v(63[16:31])
    defparam i61713_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6394_7_lut (.I0(GND_net), .I1(n17800[4]), .I2(n460_adj_4602), 
            .I3(n58619), .O(n17257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_7 (.CI(n58619), .I0(n17800[4]), .I1(n460_adj_4602), 
            .CO(n58620));
    SB_LUT4 add_6394_6_lut (.I0(GND_net), .I1(n17800[3]), .I2(n387_adj_4601), 
            .I3(n58618), .O(n17257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_16 (.CI(n58181), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n58182));
    SB_CARRY add_6394_6 (.CI(n58618), .I0(n17800[3]), .I1(n387_adj_4601), 
            .CO(n58619));
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n58180), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n58180), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n58181));
    SB_LUT4 add_6394_5_lut (.I0(GND_net), .I1(n17800[2]), .I2(n314_adj_4590), 
            .I3(n58617), .O(n17257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n58179), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n58179), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n58180));
    SB_CARRY add_6394_5 (.CI(n58617), .I0(n17800[2]), .I1(n314_adj_4590), 
            .CO(n58618));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n58178), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n58178), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n58179));
    SB_LUT4 add_6394_4_lut (.I0(GND_net), .I1(n17800[1]), .I2(n241_adj_4583), 
            .I3(n58616), .O(n17257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n58177), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_4 (.CI(n58616), .I0(n17800[1]), .I1(n241_adj_4583), 
            .CO(n58617));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[18]), 
            .I3(n58331), .O(n291)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(control_update), .I1(n25794), .I2(n105), .I3(GND_net), 
            .O(n7054));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 LessThan_28_i35_2_lut (.I0(n455[17]), .I1(n48[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4877));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i7_2_lut (.I0(n455[3]), .I1(n48[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4878));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6394_3_lut (.I0(GND_net), .I1(n17800[0]), .I2(n168), .I3(n58615), 
            .O(n17257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_3 (.CI(n58615), .I0(n17800[0]), .I1(n168), .CO(n58616));
    SB_LUT4 add_6394_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6394_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6394_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n58615));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n58331), .I0(GND_net), .I1(n1_adj_4996[18]), 
            .CO(n58332));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[17]), 
            .I3(n58330), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i9_2_lut (.I0(n475), .I1(n48[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4879));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4610));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i31_2_lut (.I0(n455[15]), .I1(n48[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4880));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n58330), .I0(GND_net), .I1(n1_adj_4996[17]), 
            .CO(n58331));
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4609));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[16]), 
            .I3(n58329), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i23_2_lut (.I0(n455[11]), .I1(n48[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4881));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n58329), .I0(GND_net), .I1(n1_adj_4996[16]), 
            .CO(n58330));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[15]), 
            .I3(n58328), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i25_2_lut (.I0(n467), .I1(n48[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4882));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4608));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_17 (.CI(n58328), .I0(GND_net), .I1(n1_adj_4996[15]), 
            .CO(n58329));
    SB_LUT4 LessThan_28_i33_2_lut (.I0(n455[16]), .I1(n48[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4883));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4607));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i29_2_lut (.I0(n455[14]), .I1(n48[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4884));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i27_2_lut (.I0(n455[13]), .I1(n48[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4885));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i17_2_lut (.I0(n455[8]), .I1(n48[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4886));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i19_2_lut (.I0(n455[9]), .I1(n48[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4887));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i21_2_lut (.I0(n455[10]), .I1(n48[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4888));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i11_2_lut (.I0(n455[5]), .I1(n48[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4889));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i13_2_lut (.I0(n455[6]), .I1(n48[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4890));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i15_2_lut (.I0(n455[7]), .I1(n48[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4891));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4604));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59323_4_lut (.I0(n27_adj_4885), .I1(n15_adj_4891), .I2(n13_adj_4890), 
            .I3(n11_adj_4889), .O(n75158));
    defparam i59323_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i60320_4_lut (.I0(n9_adj_4879), .I1(n7_adj_4878), .I2(n455[2]), 
            .I3(n48[2]), .O(n76155));
    defparam i60320_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i60843_4_lut (.I0(n15_adj_4891), .I1(n13_adj_4890), .I2(n11_adj_4889), 
            .I3(n76155), .O(n76678));
    defparam i60843_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i60841_4_lut (.I0(n21_adj_4888), .I1(n19_adj_4887), .I2(n17_adj_4886), 
            .I3(n76678), .O(n76676));
    defparam i60841_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59327_4_lut (.I0(n27_adj_4885), .I1(n25_adj_4882), .I2(n23_adj_4881), 
            .I3(n76676), .O(n75162));
    defparam i59327_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59216_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n75051));
    defparam i59216_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n48[7]), .I1(n48[16]), .I2(n33_adj_4883), 
            .I3(GND_net), .O(n12_adj_4892));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4599));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n74481), .I1(n48[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_4893));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61201_3_lut (.I0(n4_adj_4893), .I1(n48[13]), .I2(n27_adj_4885), 
            .I3(GND_net), .O(n77036));   // verilog/motorControl.v(62[35:55])
    defparam i61201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4598));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61202_3_lut (.I0(n77036), .I1(n48[14]), .I2(n29_adj_4884), 
            .I3(GND_net), .O(n77037));   // verilog/motorControl.v(62[35:55])
    defparam i61202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n48[5]), .I1(n48[6]), .I2(n13_adj_4890), 
            .I3(GND_net), .O(n10_adj_4894));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n351));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4596));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_4892), .I1(n48[17]), .I2(n35_adj_4877), 
            .I3(GND_net), .O(n30_adj_4896));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59319_4_lut (.I0(n33_adj_4883), .I1(n31_adj_4880), .I2(n29_adj_4884), 
            .I3(n75158), .O(n75154));
    defparam i59319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4595));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61073_4_lut (.I0(n30_adj_4896), .I1(n10_adj_4894), .I2(n35_adj_4877), 
            .I3(n75152), .O(n76908));   // verilog/motorControl.v(62[35:55])
    defparam i61073_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_12 (.CI(n58177), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n58178));
    SB_LUT4 i60022_3_lut (.I0(n77037), .I1(n48[15]), .I2(n31_adj_4880), 
            .I3(GND_net), .O(n75857));   // verilog/motorControl.v(62[35:55])
    defparam i60022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n48[4]), .I1(n48[8]), .I2(n17_adj_4886), 
            .I3(GND_net), .O(n8_adj_4897));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4592));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i6_3_lut (.I0(n48[2]), .I1(n48[3]), .I2(n7_adj_4878), 
            .I3(GND_net), .O(n6_adj_4898));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[14]), 
            .I3(n58327), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6610_8_lut (.I0(GND_net), .I1(n20348[5]), .I2(n560), .I3(n58598), 
            .O(n20254[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n8_adj_4897), .I1(n48[9]), .I2(n19_adj_4887), 
            .I3(GND_net), .O(n16_adj_4899));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6610_7_lut (.I0(GND_net), .I1(n20348[4]), .I2(n487), .I3(n58597), 
            .O(n20254[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61620_4_lut (.I0(n16_adj_4899), .I1(n6_adj_4898), .I2(n19_adj_4887), 
            .I3(n75200), .O(n77455));   // verilog/motorControl.v(62[35:55])
    defparam i61620_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_6610_7 (.CI(n58597), .I0(n20348[4]), .I1(n487), .CO(n58598));
    SB_LUT4 i61621_3_lut (.I0(n77455), .I1(n48[10]), .I2(n21_adj_4888), 
            .I3(GND_net), .O(n77456));   // verilog/motorControl.v(62[35:55])
    defparam i61621_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n58327), .I0(GND_net), .I1(n1_adj_4996[14]), 
            .CO(n58328));
    SB_LUT4 i61469_3_lut (.I0(n77456), .I1(n48[11]), .I2(n23_adj_4881), 
            .I3(GND_net), .O(n77304));   // verilog/motorControl.v(62[35:55])
    defparam i61469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[13]), 
            .I3(n58326), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n460_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6610_6_lut (.I0(GND_net), .I1(n20348[3]), .I2(n414), .I3(n58596), 
            .O(n20254[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n58326), .I0(GND_net), .I1(n1_adj_4996[13]), 
            .CO(n58327));
    SB_CARRY add_6610_6 (.CI(n58596), .I0(n20348[3]), .I1(n414), .CO(n58597));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[12]), 
            .I3(n58325), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n58325), .I0(GND_net), .I1(n1_adj_4996[12]), 
            .CO(n58326));
    SB_LUT4 add_6610_5_lut (.I0(GND_net), .I1(n20348[2]), .I2(n341), .I3(n58595), 
            .O(n20254[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6610_5 (.CI(n58595), .I0(n20348[2]), .I1(n341), .CO(n58596));
    SB_LUT4 add_6610_4_lut (.I0(GND_net), .I1(n20348[1]), .I2(n268), .I3(n58594), 
            .O(n20254[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61268_4_lut (.I0(n33_adj_4883), .I1(n31_adj_4880), .I2(n29_adj_4884), 
            .I3(n75162), .O(n77103));
    defparam i61268_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_6610_4 (.CI(n58594), .I0(n20348[1]), .I1(n268), .CO(n58595));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[11]), 
            .I3(n58324), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6610_3_lut (.I0(GND_net), .I1(n20348[0]), .I2(n195), .I3(n58593), 
            .O(n20254[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n58324), .I0(GND_net), .I1(n1_adj_4996[11]), 
            .CO(n58325));
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6610_3 (.CI(n58593), .I0(n20348[0]), .I1(n195), .CO(n58594));
    SB_LUT4 add_6610_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20254[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6610_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6610_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n58593));
    SB_LUT4 add_6425_16_lut (.I0(GND_net), .I1(n18279[13]), .I2(n1120), 
            .I3(n58592), .O(n17800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[10]), 
            .I3(n58323), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61586_4_lut (.I0(n75857), .I1(n76908), .I2(n35_adj_4877), 
            .I3(n75154), .O(n77421));   // verilog/motorControl.v(62[35:55])
    defparam i61586_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n58323), .I0(GND_net), .I1(n1_adj_4996[10]), 
            .CO(n58324));
    SB_LUT4 i60020_3_lut (.I0(n77304), .I1(n48[12]), .I2(n25_adj_4882), 
            .I3(GND_net), .O(n75855));   // verilog/motorControl.v(62[35:55])
    defparam i60020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61588_4_lut (.I0(n75855), .I1(n77421), .I2(n35_adj_4877), 
            .I3(n77103), .O(n77423));   // verilog/motorControl.v(62[35:55])
    defparam i61588_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_28_i38_3_lut (.I0(n77423), .I1(n48[18]), .I2(n455[18]), 
            .I3(GND_net), .O(n38_adj_2));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6425_15_lut (.I0(GND_net), .I1(n18279[12]), .I2(n1047), 
            .I3(n58591), .O(n17800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_15 (.CI(n58591), .I0(n18279[12]), .I1(n1047), .CO(n58592));
    SB_LUT4 LessThan_26_i37_2_lut (.I0(deadband[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4903));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6425_14_lut (.I0(GND_net), .I1(n18279[11]), .I2(n974), 
            .I3(n58590), .O(n17800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n11920[0]), .I2(n12496[0]), 
            .I3(n58236), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(deadband[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4904));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6425_14 (.CI(n58590), .I0(n18279[11]), .I1(n974), .CO(n58591));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[9]), 
            .I3(n58322), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4905));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n58322), .I0(GND_net), .I1(n1_adj_4996[9]), 
            .CO(n58323));
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n46[22]), 
            .I3(n58235), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6425_13_lut (.I0(GND_net), .I1(n18279[10]), .I2(n901), 
            .I3(n58589), .O(n17800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(deadband[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4906));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6425_13 (.CI(n58589), .I0(n18279[10]), .I1(n901), .CO(n58590));
    SB_LUT4 add_6425_12_lut (.I0(GND_net), .I1(n18279[9]), .I2(n828), 
            .I3(n58588), .O(n17800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(deadband[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4907));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6425_12 (.CI(n58588), .I0(n18279[9]), .I1(n828), .CO(n58589));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[8]), 
            .I3(n58321), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n58321), .I0(GND_net), .I1(n1_adj_4996[8]), 
            .CO(n58322));
    SB_LUT4 add_6425_11_lut (.I0(GND_net), .I1(n18279[8]), .I2(n755), 
            .I3(n58587), .O(n17800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_11 (.CI(n58587), .I0(n18279[8]), .I1(n755), .CO(n58588));
    SB_LUT4 add_6425_10_lut (.I0(GND_net), .I1(n18279[7]), .I2(n682), 
            .I3(n58586), .O(n17800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_10 (.CI(n58586), .I0(n18279[7]), .I1(n682), .CO(n58587));
    SB_CARRY add_25_24 (.CI(n58235), .I0(n360[22]), .I1(n46[22]), .CO(n58236));
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n46[21]), 
            .I3(n58234), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_9_lut (.I0(GND_net), .I1(n18279[6]), .I2(n609), .I3(n58585), 
            .O(n17800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_9 (.CI(n58585), .I0(n18279[6]), .I1(n609), .CO(n58586));
    SB_LUT4 add_6425_8_lut (.I0(GND_net), .I1(n18279[5]), .I2(n536), .I3(n58584), 
            .O(n17800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n58234), .I0(n360[21]), .I1(n46[21]), .CO(n58235));
    SB_LUT4 LessThan_26_i33_2_lut (.I0(deadband[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4908));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_4909));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_6425_8 (.CI(n58584), .I0(n18279[5]), .I1(n536), .CO(n58585));
    SB_LUT4 add_6425_7_lut (.I0(GND_net), .I1(n18279[4]), .I2(n463), .I3(n58583), 
            .O(n17800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_7 (.CI(n58583), .I0(n18279[4]), .I1(n463), .CO(n58584));
    SB_LUT4 add_6425_6_lut (.I0(GND_net), .I1(n18279[3]), .I2(n390_adj_4549), 
            .I3(n58582), .O(n17800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i61071_3_lut (.I0(n4_adj_4909), .I1(n455[2]), .I2(deadband[2]), 
            .I3(GND_net), .O(n76906));   // verilog/motorControl.v(62[14:31])
    defparam i61071_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61072_3_lut (.I0(n76906), .I1(n455[3]), .I2(deadband[3]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(62[14:31])
    defparam i61072_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4911));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6425_6 (.CI(n58582), .I0(n18279[3]), .I1(n390_adj_4549), 
            .CO(n58583));
    SB_LUT4 add_6425_5_lut (.I0(GND_net), .I1(n18279[2]), .I2(n317_adj_4548), 
            .I3(n58581), .O(n17800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_5 (.CI(n58581), .I0(n18279[2]), .I1(n317_adj_4548), 
            .CO(n58582));
    SB_LUT4 add_6425_4_lut (.I0(GND_net), .I1(n18279[1]), .I2(n244_adj_4546), 
            .I3(n58580), .O(n17800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n59529), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n59528), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_4 (.CI(n58580), .I0(n18279[1]), .I1(n244_adj_4546), 
            .CO(n58581));
    SB_LUT4 add_6425_3_lut (.I0(GND_net), .I1(n18279[0]), .I2(n171), .I3(n58579), 
            .O(n17800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_3 (.CI(n58579), .I0(n18279[0]), .I1(n171), .CO(n58580));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n46[20]), 
            .I3(n58233), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6425_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n17800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6425_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6425_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n58579));
    SB_CARRY add_25_22 (.CI(n58233), .I0(n360[20]), .I1(n46[20]), .CO(n58234));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n46[19]), 
            .I3(n58232), .O(n460)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n58232), .I0(n360[19]), .I1(n46[19]), .CO(n58233));
    SB_CARRY counter_2045_2046_add_4_14 (.CI(n59528), .I0(GND_net), .I1(counter[12]), 
            .CO(n59529));
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n46[18]), 
            .I3(n58231), .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n58231), .I0(n360[18]), .I1(n46[18]), .CO(n58232));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n46[17]), 
            .I3(n58230), .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n58230), .I0(n360[17]), .I1(n46[17]), .CO(n58231));
    SB_LUT4 counter_2045_2046_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n59527), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(deadband[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4912));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4913));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4914));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n46[16]), 
            .I3(n58229), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59240_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n75075));
    defparam i59240_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_25_18 (.CI(n58229), .I0(n360[16]), .I1(n46[16]), .CO(n58230));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n46[15]), 
            .I3(n58228), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4915));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_25_17 (.CI(n58228), .I0(n360[15]), .I1(n46[15]), .CO(n58229));
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n46[14]), 
            .I3(n58227), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_15_lut (.I0(GND_net), .I1(n18698[12]), .I2(n1050), 
            .I3(n58563), .O(n18279[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_13 (.CI(n59527), .I0(GND_net), .I1(counter[11]), 
            .CO(n59528));
    SB_LUT4 add_6454_14_lut (.I0(GND_net), .I1(n18698[11]), .I2(n977), 
            .I3(n58562), .O(n18279[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n59526), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_12 (.CI(n59526), .I0(GND_net), .I1(counter[10]), 
            .CO(n59527));
    SB_CARRY add_25_16 (.CI(n58227), .I0(n360[14]), .I1(n46[14]), .CO(n58228));
    SB_CARRY add_6454_14 (.CI(n58562), .I0(n18698[11]), .I1(n977), .CO(n58563));
    SB_LUT4 add_6454_13_lut (.I0(GND_net), .I1(n18698[10]), .I2(n904_adj_4540), 
            .I3(n58561), .O(n18279[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n46[13]), 
            .I3(n58226), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_13 (.CI(n58561), .I0(n18698[10]), .I1(n904_adj_4540), 
            .CO(n58562));
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n59525), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4916));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6454_12_lut (.I0(GND_net), .I1(n18698[9]), .I2(n831_adj_4539), 
            .I3(n58560), .O(n18279[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_12 (.CI(n58560), .I0(n18698[9]), .I1(n831_adj_4539), 
            .CO(n58561));
    SB_CARRY counter_2045_2046_add_4_11 (.CI(n59525), .I0(GND_net), .I1(counter[9]), 
            .CO(n59526));
    SB_LUT4 i59416_2_lut_4_lut (.I0(deadband[11]), .I1(n455[11]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n75251));
    defparam i59416_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4917));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 counter_2045_2046_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n59524), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_11_lut (.I0(GND_net), .I1(n18698[8]), .I2(n758_adj_4538), 
            .I3(n58559), .O(n18279[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_10 (.CI(n59524), .I0(GND_net), .I1(counter[8]), 
            .CO(n59525));
    SB_LUT4 counter_2045_2046_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n59523), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_11 (.CI(n58559), .I0(n18698[8]), .I1(n758_adj_4538), 
            .CO(n58560));
    SB_LUT4 i60366_4_lut (.I0(n15_adj_4917), .I1(n13_adj_4916), .I2(deadband[5]), 
            .I3(n455[5]), .O(n76201));
    defparam i60366_4_lut.LUT_INIT = 16'heffe;
    SB_CARRY counter_2045_2046_add_4_9 (.CI(n59523), .I0(GND_net), .I1(counter[7]), 
            .CO(n59524));
    SB_LUT4 i60871_4_lut (.I0(n21_adj_4915), .I1(n19_adj_4914), .I2(n17_adj_4913), 
            .I3(n76201), .O(n76706));
    defparam i60871_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 counter_2045_2046_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n59522), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_10_lut (.I0(GND_net), .I1(n18698[7]), .I2(n685_adj_4535), 
            .I3(n58558), .O(n18279[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_8 (.CI(n59522), .I0(GND_net), .I1(counter[6]), 
            .CO(n59523));
    SB_CARRY add_6454_10 (.CI(n58558), .I0(n18698[7]), .I1(n685_adj_4535), 
            .CO(n58559));
    SB_LUT4 counter_2045_2046_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n59521), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_9_lut (.I0(GND_net), .I1(n18698[6]), .I2(n612_adj_4534), 
            .I3(n58557), .O(n18279[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_7 (.CI(n59521), .I0(GND_net), .I1(counter[5]), 
            .CO(n59522));
    SB_CARRY add_6454_9 (.CI(n58557), .I0(n18698[6]), .I1(n612_adj_4534), 
            .CO(n58558));
    SB_LUT4 add_6454_8_lut (.I0(GND_net), .I1(n18698[5]), .I2(n539_adj_4533), 
            .I3(n58556), .O(n18279[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n58226), .I0(n360[13]), .I1(n46[13]), .CO(n58227));
    SB_CARRY add_6454_8 (.CI(n58556), .I0(n18698[5]), .I1(n539_adj_4533), 
            .CO(n58557));
    SB_LUT4 add_6454_7_lut (.I0(GND_net), .I1(n18698[4]), .I2(n466_adj_4531), 
            .I3(n58555), .O(n18279[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n46[12]), 
            .I3(n58225), .O(n467)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n59520), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i60869_4_lut (.I0(n27_adj_4912), .I1(n25_adj_3), .I2(n23_adj_4911), 
            .I3(n76706), .O(n76704));
    defparam i60869_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i59402_4_lut (.I0(n33_adj_4908), .I1(n31_adj_4907), .I2(n29_adj_4906), 
            .I3(n76704), .O(n75237));
    defparam i59402_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY counter_2045_2046_add_4_6 (.CI(n59520), .I0(GND_net), .I1(counter[4]), 
            .CO(n59521));
    SB_LUT4 counter_2045_2046_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n59519), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_7 (.CI(n58555), .I0(n18698[4]), .I1(n466_adj_4531), 
            .CO(n58556));
    SB_LUT4 add_6454_6_lut (.I0(GND_net), .I1(n18698[3]), .I2(n393_adj_4530), 
            .I3(n58554), .O(n18279[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n58225), .I0(n360[12]), .I1(n46[12]), .CO(n58226));
    SB_CARRY add_6454_6 (.CI(n58554), .I0(n18698[3]), .I1(n393_adj_4530), 
            .CO(n58555));
    SB_LUT4 add_6454_5_lut (.I0(GND_net), .I1(n18698[2]), .I2(n320_adj_4529), 
            .I3(n58553), .O(n18279[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_5 (.CI(n59519), .I0(GND_net), .I1(counter[3]), 
            .CO(n59520));
    SB_LUT4 counter_2045_2046_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n59518), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n46[11]), 
            .I3(n58224), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6454_5 (.CI(n58553), .I0(n18698[2]), .I1(n320_adj_4529), 
            .CO(n58554));
    SB_LUT4 add_6454_4_lut (.I0(GND_net), .I1(n18698[1]), .I2(n247_adj_4527), 
            .I3(n58552), .O(n18279[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n58224), .I0(n360[11]), .I1(n46[11]), .CO(n58225));
    SB_CARRY add_6454_4 (.CI(n58552), .I0(n18698[1]), .I1(n247_adj_4527), 
            .CO(n58553));
    SB_CARRY counter_2045_2046_add_4_4 (.CI(n59518), .I0(GND_net), .I1(counter[2]), 
            .CO(n59519));
    SB_LUT4 i61225_3_lut (.I0(n10), .I1(n455[16]), .I2(n33_adj_4908), 
            .I3(GND_net), .O(n77060));   // verilog/motorControl.v(62[14:31])
    defparam i61225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2045_2046_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n59517), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i59390_2_lut_4_lut (.I0(deadband[19]), .I1(n460), .I2(deadband[10]), 
            .I3(n455[10]), .O(n75225));
    defparam i59390_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_6454_3_lut (.I0(GND_net), .I1(n18698[0]), .I2(n174_adj_4525), 
            .I3(n58551), .O(n18279[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_3 (.CI(n59517), .I0(GND_net), .I1(counter[1]), 
            .CO(n59518));
    SB_CARRY add_6454_3 (.CI(n58551), .I0(n18698[0]), .I1(n174_adj_4525), 
            .CO(n58552));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n46[10]), 
            .I3(n58223), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6454_2_lut (.I0(GND_net), .I1(n32_adj_4523), .I2(n101_adj_4522), 
            .I3(GND_net), .O(n18279[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6454_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i18_3_lut (.I0(n455[10]), .I1(n460), .I2(n39), 
            .I3(GND_net), .O(n18_adj_4921));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6454_2 (.CI(GND_net), .I0(n32_adj_4523), .I1(n101_adj_4522), 
            .CO(n58551));
    SB_CARRY add_25_12 (.CI(n58223), .I0(n360[10]), .I1(n46[10]), .CO(n58224));
    SB_LUT4 counter_2045_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n59517));
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[8]), .I1(n455[9]), .I2(n19_adj_4914), 
            .I3(GND_net), .O(n16_adj_4922));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n46[9]), .I3(n58222), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_11 (.CI(n58222), .I0(n360[9]), .I1(n46[9]), .CO(n58223));
    SB_LUT4 i59365_2_lut_4_lut (.I0(n455[8]), .I1(n48[8]), .I2(n475), 
            .I3(n48[4]), .O(n75200));
    defparam i59365_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n46[8]), .I3(n58221), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_10 (.CI(n58221), .I0(n360[8]), .I1(n46[8]), .CO(n58222));
    SB_LUT4 i59317_2_lut_4_lut (.I0(n455[16]), .I1(n48[16]), .I2(n455[7]), 
            .I3(n48[7]), .O(n75152));
    defparam i59317_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n46[7]), .I3(n58220), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_9 (.CI(n58220), .I0(n360[7]), .I1(n46[7]), .CO(n58221));
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n46[6]), .I3(n58219), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11880_bdd_4_lut_62795 (.I0(n11880), .I1(n74594), .I2(setpoint[2]), 
            .I3(n4734), .O(n78657));
    defparam n11880_bdd_4_lut_62795.LUT_INIT = 16'he4aa;
    SB_CARRY add_25_8 (.CI(n58219), .I0(n360[6]), .I1(n46[6]), .CO(n58220));
    SB_LUT4 n78657_bdd_4_lut (.I0(n78657), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4734), .O(n78660));
    defparam n78657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4996[7]), 
            .I3(n58320), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n46[5]), .I3(n58218), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n58320), .I0(GND_net), .I1(n1_adj_4996[7]), 
            .CO(n58321));
    SB_LUT4 add_6622_7_lut (.I0(GND_net), .I1(n69074), .I2(n490_adj_4496), 
            .I3(n58536), .O(n20348[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i36_3_lut (.I0(n18_adj_4921), .I1(n455[20]), .I2(n41_adj_4905), 
            .I3(GND_net), .O(n36));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59400_4_lut (.I0(n33_adj_4908), .I1(n21_adj_4915), .I2(n19_adj_4914), 
            .I3(n17_adj_4913), .O(n75235));
    defparam i59400_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6622_6_lut (.I0(GND_net), .I1(n20416[3]), .I2(n417_adj_4486), 
            .I3(n58535), .O(n20348[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_6 (.CI(n58535), .I0(n20416[3]), .I1(n417_adj_4486), 
            .CO(n58536));
    SB_LUT4 add_6622_5_lut (.I0(GND_net), .I1(n20419), .I2(n344_adj_4485), 
            .I3(n58534), .O(n20348[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_5 (.CI(n58534), .I0(n20419), .I1(n344_adj_4485), 
            .CO(n58535));
    SB_LUT4 add_6622_4_lut (.I0(GND_net), .I1(n20420), .I2(n271_adj_4484), 
            .I3(n58533), .O(n20348[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_4 (.CI(n58533), .I0(n20420), .I1(n271_adj_4484), 
            .CO(n58534));
    SB_LUT4 i61226_3_lut (.I0(n77060), .I1(n455[17]), .I2(n35_adj_4904), 
            .I3(GND_net), .O(n77061));   // verilog/motorControl.v(62[14:31])
    defparam i61226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6622_3_lut (.I0(GND_net), .I1(n20416[0]), .I2(n198_adj_4483), 
            .I3(n58532), .O(n20348[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6622_3 (.CI(n58532), .I0(n20416[0]), .I1(n198_adj_4483), 
            .CO(n58533));
    SB_LUT4 i59392_4_lut (.I0(n39), .I1(n37_adj_4903), .I2(n35_adj_4904), 
            .I3(n75235), .O(n75227));
    defparam i59392_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6622_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_4482), 
            .I3(GND_net), .O(n20348[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6622_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_7 (.CI(n58218), .I0(n360[5]), .I1(n46[5]), .CO(n58219));
    SB_CARRY add_6622_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_4482), .CO(n58532));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n46[4]), .I3(n58217), 
            .O(n475)) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_14_lut (.I0(GND_net), .I1(n19061[11]), .I2(n980_adj_4481), 
            .I3(n58531), .O(n18698[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_13_lut (.I0(GND_net), .I1(n19061[10]), .I2(n907_adj_4480), 
            .I3(n58530), .O(n18698[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n58217), .I0(n360[4]), .I1(n46[4]), .CO(n58218));
    SB_CARRY add_6481_13 (.CI(n58530), .I0(n19061[10]), .I1(n907_adj_4480), 
            .CO(n58531));
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n46[3]), .I3(n58216), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6481_12_lut (.I0(GND_net), .I1(n19061[9]), .I2(n834_adj_4479), 
            .I3(n58529), .O(n18698[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_12 (.CI(n58529), .I0(n19061[9]), .I1(n834_adj_4479), 
            .CO(n58530));
    SB_CARRY add_25_5 (.CI(n58216), .I0(n360[3]), .I1(n46[3]), .CO(n58217));
    SB_LUT4 add_6481_11_lut (.I0(GND_net), .I1(n19061[8]), .I2(n761_adj_4478), 
            .I3(n58528), .O(n18698[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n46[2]), .I3(n58215), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_11 (.CI(n58528), .I0(n19061[8]), .I1(n761_adj_4478), 
            .CO(n58529));
    SB_LUT4 i61618_4_lut (.I0(n36), .I1(n16_adj_4922), .I2(n41_adj_4905), 
            .I3(n75225), .O(n77453));   // verilog/motorControl.v(62[14:31])
    defparam i61618_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60008_3_lut (.I0(n77061), .I1(n455[18]), .I2(n37_adj_4903), 
            .I3(GND_net), .O(n75843));   // verilog/motorControl.v(62[14:31])
    defparam i60008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6481_10_lut (.I0(GND_net), .I1(n19061[7]), .I2(n688_adj_4477), 
            .I3(n58527), .O(n18698[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_4 (.CI(n58215), .I0(n360[2]), .I1(n46[2]), .CO(n58216));
    SB_CARRY add_6481_10 (.CI(n58527), .I0(n19061[7]), .I1(n688_adj_4477), 
            .CO(n58528));
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n46[1]), .I3(n58214), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i42_3_lut (.I0(n48[20]), .I1(n48[21]), .I2(n455[21]), 
            .I3(GND_net), .O(n42));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_6481_9_lut (.I0(GND_net), .I1(n19061[6]), .I2(n615), .I3(n58526), 
            .O(n18698[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_9 (.CI(n58526), .I0(n19061[6]), .I1(n615), .CO(n58527));
    SB_LUT4 i59313_4_lut (.I0(n455[21]), .I1(n455[20]), .I2(n48[21]), 
            .I3(n48[20]), .O(n75148));
    defparam i59313_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 add_6481_8_lut (.I0(GND_net), .I1(n19061[5]), .I2(n542), .I3(n58525), 
            .O(n18698[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i45_rep_158_2_lut (.I0(n455[22]), .I1(n48[22]), 
            .I2(GND_net), .I3(GND_net), .O(n79219));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_rep_158_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6481_8 (.CI(n58525), .I0(n19061[5]), .I1(n542), .CO(n58526));
    SB_LUT4 add_6481_7_lut (.I0(GND_net), .I1(n19061[4]), .I2(n469_adj_4476), 
            .I3(n58524), .O(n18698[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_7 (.CI(n58524), .I0(n19061[4]), .I1(n469_adj_4476), 
            .CO(n58525));
    SB_LUT4 add_6481_6_lut (.I0(GND_net), .I1(n19061[3]), .I2(n396), .I3(n58523), 
            .O(n18698[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6481_6 (.CI(n58523), .I0(n19061[3]), .I1(n396), .CO(n58524));
    SB_LUT4 add_6481_5_lut (.I0(GND_net), .I1(n19061[2]), .I2(n323), .I3(n58522), 
            .O(n18698[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6481_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i44_3_lut (.I0(n42), .I1(n48[22]), .I2(n455[22]), 
            .I3(GND_net), .O(n44_adj_4924));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i44_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61075_4_lut (.I0(n44_adj_4924), .I1(n40), .I2(n79219), .I3(n75148), 
            .O(n76910));   // verilog/motorControl.v(62[35:55])
    defparam i61075_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 LessThan_26_i14_3_lut (.I0(n455[7]), .I1(n455[11]), .I2(n23_adj_4911), 
            .I3(GND_net), .O(n14_adj_4925));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59283_2_lut_4_lut (.I0(PWMLimit[19]), .I1(n460), .I2(PWMLimit[15]), 
            .I3(n455[15]), .O(n75118));
    defparam i59283_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4916), 
            .I3(GND_net), .O(n12_adj_4926));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i22_3_lut (.I0(n14_adj_4925), .I1(n467), .I2(n25_adj_3), 
            .I3(GND_net), .O(n22_adj_4927));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61616_4_lut (.I0(n22_adj_4927), .I1(n12_adj_4926), .I2(n25_adj_3), 
            .I3(n75251), .O(n77451));   // verilog/motorControl.v(62[14:31])
    defparam i61616_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i61617_3_lut (.I0(n77451), .I1(n455[13]), .I2(n27_adj_4912), 
            .I3(GND_net), .O(n77452));   // verilog/motorControl.v(62[14:31])
    defparam i61617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61477_3_lut (.I0(n77452), .I1(n455[14]), .I2(n29_adj_4906), 
            .I3(GND_net), .O(n77312));   // verilog/motorControl.v(62[14:31])
    defparam i61477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61292_4_lut (.I0(n39), .I1(n37_adj_4903), .I2(n35_adj_4904), 
            .I3(n75237), .O(n77127));
    defparam i61292_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i61760_4_lut (.I0(n75843), .I1(n77453), .I2(n41_adj_4905), 
            .I3(n75227), .O(n77595));   // verilog/motorControl.v(62[14:31])
    defparam i61760_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60006_3_lut (.I0(n77312), .I1(n455[15]), .I2(n31_adj_4907), 
            .I3(GND_net), .O(n75841));   // verilog/motorControl.v(62[14:31])
    defparam i60006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61808_4_lut (.I0(n75841), .I1(n77595), .I2(n41_adj_4905), 
            .I3(n77127), .O(n77643));   // verilog/motorControl.v(62[14:31])
    defparam i61808_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i59299_2_lut_4_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(PWMLimit[4]), 
            .I3(n475), .O(n75134));
    defparam i59299_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61809_3_lut (.I0(n77643), .I1(n455[21]), .I2(deadband[21]), 
            .I3(GND_net), .O(n77644));   // verilog/motorControl.v(62[14:31])
    defparam i61809_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i61076_3_lut (.I0(n76910), .I1(n455[23]), .I2(n47_adj_4849), 
            .I3(GND_net), .O(n76911));   // verilog/motorControl.v(62[35:55])
    defparam i61076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61807_3_lut (.I0(n77644), .I1(n455[22]), .I2(deadband[22]), 
            .I3(GND_net), .O(n77642));   // verilog/motorControl.v(62[14:31])
    defparam i61807_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30514_4_lut (.I0(n77642), .I1(n76911), .I2(deadband[23]), 
            .I3(n455[23]), .O(n44588));
    defparam i30514_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 n11880_bdd_4_lut_63013 (.I0(n11880), .I1(n74632), .I2(setpoint[22]), 
            .I3(n4734), .O(n78903));
    defparam n11880_bdd_4_lut_63013.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_9_i24_3_lut_3_lut (.I0(setpoint[11]), .I1(setpoint[12]), 
            .I2(PWMLimit[12]), .I3(GND_net), .O(n24_adj_4845));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut_adj_957 (.I0(n7052), .I1(n7054), .I2(n25756), .I3(n67040), 
            .O(n4734));
    defparam i3_4_lut_adj_957.LUT_INIT = 16'hefff;
    SB_LUT4 i59721_2_lut_4_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), .I2(PWMLimit[13]), 
            .I3(setpoint[13]), .O(n75556));
    defparam i59721_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i59246_4_lut (.I0(n27), .I1(n15_adj_4722), .I2(n13_adj_4723), 
            .I3(n11_adj_4721), .O(n75081));
    defparam i59246_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_c), 
            .I3(GND_net), .O(n12_adj_4928));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4723), 
            .I3(GND_net), .O(n10_adj_4929));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_4928), .I1(n535[17]), .I2(n35_adj_4719), 
            .I3(GND_net), .O(n30_adj_4930));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i26_3_lut_3_lut (.I0(setpoint[13]), .I1(setpoint[17]), 
            .I2(PWMLimit[17]), .I3(GND_net), .O(n26_adj_4843));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i60240_4_lut (.I0(n13_adj_4723), .I1(n11_adj_4721), .I2(n9_adj_4716), 
            .I3(n75112), .O(n76075));
    defparam i60240_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60236_4_lut (.I0(n19_adj_4715), .I1(n17_adj_4714), .I2(n15_adj_4722), 
            .I3(n76075), .O(n76071));
    defparam i60236_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61466_4_lut (.I0(n25_adj_4713), .I1(n23_adj_4712), .I2(n21_adj_4711), 
            .I3(n76071), .O(n77301));
    defparam i61466_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i60793_4_lut (.I0(n31), .I1(n29_adj_4709), .I2(n27), .I3(n77301), 
            .O(n76628));
    defparam i60793_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61640_4_lut (.I0(n37_c), .I1(n35_adj_4719), .I2(n33_c), .I3(n76628), 
            .O(n77475));
    defparam i61640_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i61191_3_lut (.I0(n6_adj_4931), .I1(n535[10]), .I2(n21_adj_4711), 
            .I3(GND_net), .O(n77026));   // verilog/motorControl.v(65[25:41])
    defparam i61191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61192_3_lut (.I0(n77026), .I1(n535[11]), .I2(n23_adj_4712), 
            .I3(GND_net), .O(n77027));   // verilog/motorControl.v(65[25:41])
    defparam i61192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4932));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4714), 
            .I3(GND_net), .O(n8_adj_4933));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_4932), .I1(n535[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4934));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59260_4_lut (.I0(n21_adj_4711), .I1(n19_adj_4715), .I2(n17_adj_4714), 
            .I3(n9_adj_4716), .O(n75095));
    defparam i59260_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59222_4_lut (.I0(n43), .I1(n25_adj_4713), .I2(n23_adj_4712), 
            .I3(n75095), .O(n75057));
    defparam i59222_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61079_4_lut (.I0(n24_adj_4934), .I1(n8_adj_4933), .I2(n45), 
            .I3(n75051), .O(n76914));   // verilog/motorControl.v(65[25:41])
    defparam i61079_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60034_3_lut (.I0(n77027), .I1(n535[12]), .I2(n25_adj_4713), 
            .I3(GND_net), .O(n75869));   // verilog/motorControl.v(65[25:41])
    defparam i60034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_4935));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i60791_3_lut (.I0(n4_adj_4935), .I1(n535[13]), .I2(n27), .I3(GND_net), 
            .O(n76626));   // verilog/motorControl.v(65[25:41])
    defparam i60791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60792_3_lut (.I0(n76626), .I1(n535[14]), .I2(n29_adj_4709), 
            .I3(GND_net), .O(n76627));   // verilog/motorControl.v(65[25:41])
    defparam i60792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59731_2_lut_4_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), .I2(PWMLimit[14]), 
            .I3(setpoint[14]), .O(n75566));
    defparam i59731_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i28_3_lut_3_lut (.I0(setpoint[14]), .I1(setpoint[15]), 
            .I2(PWMLimit[15]), .I3(GND_net), .O(n28));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i59242_4_lut (.I0(n33_c), .I1(n31), .I2(n29_adj_4709), .I3(n75081), 
            .O(n75077));
    defparam i59242_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61430_4_lut (.I0(n30_adj_4930), .I1(n10_adj_4929), .I2(n35_adj_4719), 
            .I3(n75075), .O(n77265));   // verilog/motorControl.v(65[25:41])
    defparam i61430_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i60036_3_lut (.I0(n76627), .I1(n535[15]), .I2(n31), .I3(GND_net), 
            .O(n75871));   // verilog/motorControl.v(65[25:41])
    defparam i60036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61697_4_lut (.I0(n75871), .I1(n77265), .I2(n35_adj_4719), 
            .I3(n75077), .O(n77532));   // verilog/motorControl.v(65[25:41])
    defparam i61697_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61698_3_lut (.I0(n77532), .I1(n535[18]), .I2(n37_c), .I3(GND_net), 
            .O(n77533));   // verilog/motorControl.v(65[25:41])
    defparam i61698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61643_3_lut (.I0(n77533), .I1(n535[19]), .I2(n39_c), .I3(GND_net), 
            .O(n77478));   // verilog/motorControl.v(65[25:41])
    defparam i61643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59230_4_lut (.I0(n43), .I1(n41_adj_4705), .I2(n39_c), .I3(n77475), 
            .O(n75065));
    defparam i59230_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59575_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n75410));
    defparam i59575_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61386_4_lut (.I0(n75869), .I1(n76914), .I2(n45), .I3(n75057), 
            .O(n77221));   // verilog/motorControl.v(65[25:41])
    defparam i61386_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60042_3_lut (.I0(n77478), .I1(n535[20]), .I2(n41_adj_4705), 
            .I3(GND_net), .O(n75877));   // verilog/motorControl.v(65[25:41])
    defparam i60042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59605_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n75440));
    defparam i59605_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i61589_4_lut (.I0(n75877), .I1(n77221), .I2(n45), .I3(n75065), 
            .O(n77424));   // verilog/motorControl.v(65[25:41])
    defparam i61589_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n11880_bdd_4_lut_62790 (.I0(n11880), .I1(n74593), .I2(setpoint[1]), 
            .I3(n4734), .O(n78651));
    defparam n11880_bdd_4_lut_62790.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut (.I0(n77424), .I1(n4_adj_4936), .I2(n455[23]), .I3(n535[23]), 
            .O(n68521));
    defparam i2_4_lut.LUT_INIT = 16'hdfcd;
    SB_LUT4 n78651_bdd_4_lut (.I0(n78651), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4734), .O(n78654));
    defparam n78651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6058_4_lut (.I0(n7052), .I1(n4734), .I2(n68521), .I3(n25798), 
            .O(n11880));
    defparam i6058_4_lut.LUT_INIT = 16'hbbab;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_adj_4937));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59571_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n75406));   // verilog/motorControl.v(56[14:36])
    defparam i59571_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59503_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n75338));   // verilog/motorControl.v(58[23:46])
    defparam i59503_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4588));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4938));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4587));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4586));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4584));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78903_bdd_4_lut (.I0(n78903), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4734), .O(n78906));
    defparam n78903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4582));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4580));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4579));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4578));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4577));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4576));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n346));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4575));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4574));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4570));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4569));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4781));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4780));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4777));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4775));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4564));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4769));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4563));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4765));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n353));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4764));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4561));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4559));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4760));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4557));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4757));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4555));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4553));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4552));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4756));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4551));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4550));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4754));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4544));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4746));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4744));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4543));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4741));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4735));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4541));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4537));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4734));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4732));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4532));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44015_2_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(\Ki[1] ), 
            .I3(n340), .O(n20466));   // verilog/motorControl.v(61[29:40])
    defparam i44015_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4528));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4524));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4521));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4519));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n354));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4517));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4516));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4703));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4702));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4701));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4699));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4514));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62993 (.I0(n11880), .I1(n74631), .I2(setpoint[21]), 
            .I3(n4734), .O(n78891));
    defparam n11880_bdd_4_lut_62993.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4698));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4697));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4696));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78891_bdd_4_lut (.I0(n78891), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4734), .O(n78894));
    defparam n78891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4695));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4513));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4693));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62983 (.I0(n11880), .I1(n74630), .I2(setpoint[20]), 
            .I3(n4734), .O(n78885));
    defparam n11880_bdd_4_lut_62983.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4512));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4510));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4509));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4692));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78885_bdd_4_lut (.I0(n78885), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4734), .O(n78888));
    defparam n78885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4690));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4508));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4506));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4505));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62978 (.I0(n11880), .I1(n74629), .I2(setpoint[19]), 
            .I3(n4734), .O(n78879));
    defparam n11880_bdd_4_lut_62978.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4689));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4503));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4688));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4501));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4500));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4499));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4498));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4687));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4686));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4495));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78879_bdd_4_lut (.I0(n78879), .I1(n535[19]), .I2(n460), .I3(n4734), 
            .O(n78882));
    defparam n78879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4685));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4494));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4684));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4493));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4683));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4681));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4680));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4492));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4488));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62973 (.I0(n11880), .I1(n74628), .I2(setpoint[18]), 
            .I3(n4734), .O(n78873));
    defparam n11880_bdd_4_lut_62973.LUT_INIT = 16'he4aa;
    SB_LUT4 n78873_bdd_4_lut (.I0(n78873), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4734), .O(n78876));
    defparam n78873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11880_bdd_4_lut_62968 (.I0(n11880), .I1(n74627), .I2(setpoint[17]), 
            .I3(n4734), .O(n78867));
    defparam n11880_bdd_4_lut_62968.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4677));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78867_bdd_4_lut (.I0(n78867), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4734), .O(n78870));
    defparam n78867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4675));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4674));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62963 (.I0(n11880), .I1(n74626), .I2(setpoint[16]), 
            .I3(n4734), .O(n78855));
    defparam n11880_bdd_4_lut_62963.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut (.I0(n25794), .I1(control_update), .I2(n44588), 
            .I3(GND_net), .O(n25754));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i51255_2_lut_3_lut (.I0(n25794), .I1(control_update), .I2(n44588), 
            .I3(GND_net), .O(n67040));
    defparam i51255_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4673));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4672));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4671));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4670));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4669));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4668));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n78855_bdd_4_lut (.I0(n78855), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4734), .O(n78858));
    defparam n78855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4667));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4666));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4665));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4664));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62785 (.I0(n11880), .I1(n74592), .I2(setpoint[0]), 
            .I3(n4734), .O(n78627));
    defparam n11880_bdd_4_lut_62785.LUT_INIT = 16'he4aa;
    SB_LUT4 n78627_bdd_4_lut (.I0(n78627), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4734), .O(n78630));
    defparam n78627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4663));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4662));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(n77548), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n25754), .O(n25756));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff71;
    SB_LUT4 i1_2_lut_4_lut_adj_958 (.I0(n77548), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n25754), .O(n4_adj_4936));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_958.LUT_INIT = 16'hff8e;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), 
            .I2(setpoint[2]), .I3(GND_net), .O(n6_adj_4829));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59762_3_lut_4_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(setpoint[2]), 
            .I3(PWMLimit[2]), .O(n75597));   // verilog/motorControl.v(45[16:33])
    defparam i59762_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_959 (.I0(n77411), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n25796), .O(n7052));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut_adj_959.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_4_lut_adj_960 (.I0(n77411), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n25796), .O(n25798));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut_adj_960.LUT_INIT = 16'h8e00;
    SB_LUT4 i59676_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n75511));   // verilog/motorControl.v(47[25:43])
    defparam i59676_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_4763));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59267_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n74624));
    defparam i59267_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59150_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[15]), 
            .I3(GND_net), .O(n74625));
    defparam i59150_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59270_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[0]), 
            .I3(GND_net), .O(n74592));
    defparam i59270_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59149_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n74626));
    defparam i59149_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59176_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n74627));
    defparam i59176_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59148_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n74628));
    defparam i59148_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59152_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n74604));
    defparam i59152_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59002_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n74603));
    defparam i59002_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59171_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n74601));
    defparam i59171_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59154_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n74600));
    defparam i59154_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59153_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n74602));
    defparam i59153_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59021_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n74599));
    defparam i59021_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i59147_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[20]), 
            .I3(GND_net), .O(n74630));
    defparam i59147_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59112_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n74615));
    defparam i59112_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59133_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n74631));
    defparam i59133_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59014_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n74593));
    defparam i59014_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59146_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n74632));
    defparam i59146_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59157_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n74594));
    defparam i59157_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4661));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59701_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[23]), 
            .I3(GND_net), .O(n74663));
    defparam i59701_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4660));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4659));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4658));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59018_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n74595));
    defparam i59018_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4657));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i59156_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[4]), 
            .I3(GND_net), .O(n74596));
    defparam i59156_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59019_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n74597));
    defparam i59019_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59155_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n74598));
    defparam i59155_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i59003_2_lut_3_lut (.I0(n7054), .I1(n25756), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n74629));
    defparam i59003_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4931));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i59277_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n75112));   // verilog/motorControl.v(65[25:41])
    defparam i59277_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i44054_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n58123));   // verilog/motorControl.v(61[20:26])
    defparam i44054_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 n11880_bdd_4_lut_62953 (.I0(n11880), .I1(n74625), .I2(setpoint[15]), 
            .I3(n4734), .O(n78843));
    defparam n11880_bdd_4_lut_62953.LUT_INIT = 16'he4aa;
    SB_LUT4 n78843_bdd_4_lut (.I0(n78843), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4734), .O(n78846));
    defparam n78843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4656));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i43865_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n57908));   // verilog/motorControl.v(61[20:26])
    defparam i43865_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i55520_2_lut (.I0(counter[13]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n71340));
    defparam i55520_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(counter[5]), .I1(counter[4]), .I2(counter[3]), 
            .I3(counter[8]), .O(n23_adj_4940));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(counter[1]), .I1(counter[6]), .I2(counter[10]), 
            .I3(counter[0]), .O(n22_adj_4941));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i12_4_lut (.I0(n23_adj_4940), .I1(counter[2]), .I2(n71340), 
            .I3(counter[9]), .O(n26_adj_4942));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i61977_4_lut (.I0(counter[12]), .I1(n26_adj_4942), .I2(n22_adj_4941), 
            .I3(counter[7]), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i61977_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4943));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4944));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4945));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4946));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4947));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4948));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4949));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4950));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4951));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4952));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4953));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4954));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4955));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4956));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4957));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4958));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4959));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59481_4_lut (.I0(n21), .I1(n19_adj_4959), .I2(n17_adj_4958), 
            .I3(n9_adj_4957), .O(n75316));
    defparam i59481_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59470_4_lut (.I0(n27_adj_4956), .I1(n15_adj_4955), .I2(n13_adj_4954), 
            .I3(n11_adj_4953), .O(n75305));
    defparam i59470_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_4952), 
            .I3(GND_net), .O(n12_adj_4961));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4954), 
            .I3(GND_net), .O(n10_adj_4962));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4961), .I1(n285[17]), .I2(n35_adj_4951), 
            .I3(GND_net), .O(n30_adj_4963));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43942_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(\Ki[1] ), 
            .I3(n37146), .O(n20499[0]));   // verilog/motorControl.v(61[29:40])
    defparam i43942_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i60434_4_lut (.I0(n13_adj_4954), .I1(n11_adj_4953), .I2(n9_adj_4957), 
            .I3(n75338), .O(n76269));
    defparam i60434_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60424_4_lut (.I0(n19_adj_4959), .I1(n17_adj_4958), .I2(n15_adj_4955), 
            .I3(n76269), .O(n76259));
    defparam i60424_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61520_4_lut (.I0(n25_adj_4948), .I1(n23_adj_4947), .I2(n21), 
            .I3(n76259), .O(n77355));
    defparam i61520_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i60891_4_lut (.I0(n31_adj_4950), .I1(n29_adj_4949), .I2(n27_adj_4956), 
            .I3(n77355), .O(n76726));
    defparam i60891_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i43944_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(\Ki[1] ), 
            .I3(n37146), .O(n57998));   // verilog/motorControl.v(61[29:40])
    defparam i43944_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i61658_4_lut (.I0(n37_adj_4), .I1(n35_adj_4951), .I2(n33_adj_4952), 
            .I3(n76726), .O(n77493));
    defparam i61658_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_4946), 
            .I3(GND_net), .O(n16_adj_4965));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61260_3_lut (.I0(n6_adj_4938), .I1(n299), .I2(n21), .I3(GND_net), 
            .O(n77095));   // verilog/motorControl.v(58[23:46])
    defparam i61260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61261_3_lut (.I0(n77095), .I1(n285[11]), .I2(n23_adj_4947), 
            .I3(GND_net), .O(n77096));   // verilog/motorControl.v(58[23:46])
    defparam i61261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_4958), 
            .I3(GND_net), .O(n8_adj_4966));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4965), .I1(n285[22]), .I2(n45_adj_4945), 
            .I3(GND_net), .O(n24_adj_4967));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59436_4_lut (.I0(n43_adj_4946), .I1(n25_adj_4948), .I2(n23_adj_4947), 
            .I3(n75316), .O(n75271));
    defparam i59436_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61069_4_lut (.I0(n24_adj_4967), .I1(n8_adj_4966), .I2(n45_adj_4945), 
            .I3(n75267), .O(n76904));   // verilog/motorControl.v(58[23:46])
    defparam i61069_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59994_3_lut (.I0(n77096), .I1(n285[12]), .I2(n25_adj_4948), 
            .I3(GND_net), .O(n75829));   // verilog/motorControl.v(58[23:46])
    defparam i59994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_4968));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i61258_3_lut (.I0(n4_adj_4968), .I1(n285[13]), .I2(n27_adj_4956), 
            .I3(GND_net), .O(n77093));   // verilog/motorControl.v(58[23:46])
    defparam i61258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61259_3_lut (.I0(n77093), .I1(n285[14]), .I2(n29_adj_4949), 
            .I3(GND_net), .O(n77094));   // verilog/motorControl.v(58[23:46])
    defparam i61259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59462_4_lut (.I0(n33_adj_4952), .I1(n31_adj_4950), .I2(n29_adj_4949), 
            .I3(n75305), .O(n75297));
    defparam i59462_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61646_4_lut (.I0(n30_adj_4963), .I1(n10_adj_4962), .I2(n35_adj_4951), 
            .I3(n75291), .O(n77481));   // verilog/motorControl.v(58[23:46])
    defparam i61646_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59996_3_lut (.I0(n77094), .I1(n285[15]), .I2(n31_adj_4950), 
            .I3(GND_net), .O(n75831));   // verilog/motorControl.v(58[23:46])
    defparam i59996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61758_4_lut (.I0(n75831), .I1(n77481), .I2(n35_adj_4951), 
            .I3(n75297), .O(n77593));   // verilog/motorControl.v(58[23:46])
    defparam i61758_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61759_3_lut (.I0(n77593), .I1(n291), .I2(n37_adj_4), .I3(GND_net), 
            .O(n77594));   // verilog/motorControl.v(58[23:46])
    defparam i61759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61718_3_lut (.I0(n77594), .I1(n285[19]), .I2(n39_adj_4944), 
            .I3(GND_net), .O(n77553));   // verilog/motorControl.v(58[23:46])
    defparam i61718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43808_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(\Ki[1] ), 
            .I3(n37336), .O(n20416[0]));   // verilog/motorControl.v(61[29:40])
    defparam i43808_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i43810_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n340), .I2(\Ki[1] ), 
            .I3(n37336), .O(n57846));   // verilog/motorControl.v(61[29:40])
    defparam i43810_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i59440_4_lut (.I0(n43_adj_4946), .I1(n41_adj_4943), .I2(n39_adj_4944), 
            .I3(n77493), .O(n75275));
    defparam i59440_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61582_4_lut (.I0(n75829), .I1(n76904), .I2(n45_adj_4945), 
            .I3(n75271), .O(n77417));   // verilog/motorControl.v(58[23:46])
    defparam i61582_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i60002_3_lut (.I0(n77553), .I1(n285[20]), .I2(n41_adj_4943), 
            .I3(GND_net), .O(n75837));   // verilog/motorControl.v(58[23:46])
    defparam i60002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61584_4_lut (.I0(n75837), .I1(n77417), .I2(n45_adj_4945), 
            .I3(n75275), .O(n77419));   // verilog/motorControl.v(58[23:46])
    defparam i61584_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Ki[3] ), .I1(n340), .I2(n4_adj_4969), 
            .I3(n20490[1]), .O(n20462[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i44036_3_lut_4_lut (.I0(\Ki[3] ), .I1(n340), .I2(n4_adj_4969), 
            .I3(n20490[1]), .O(n6_adj_4507));   // verilog/motorControl.v(61[29:40])
    defparam i44036_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i44028_3_lut_4_lut (.I0(n62_adj_4491), .I1(n131), .I2(n204), 
            .I3(n20493), .O(n4_adj_4969));   // verilog/motorControl.v(61[29:40])
    defparam i44028_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i61585_3_lut (.I0(n77419), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i61585_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_961 (.I0(n62_adj_4491), .I1(n131), .I2(n204), 
            .I3(n20493), .O(n20465));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_961.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4970));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4971));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4972));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4973));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n239), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4974));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4975));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4976));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4977));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4978));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4979));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4980));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4981));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4982));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4983));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4984));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4985));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4986));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4987));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n247), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4988));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i59553_4_lut (.I0(n21_adj_4988), .I1(n19_adj_4987), .I2(n17_adj_4986), 
            .I3(n9_adj_4985), .O(n75388));
    defparam i59553_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i59541_4_lut (.I0(n27_adj_4983), .I1(n15_adj_4982), .I2(n13_adj_4981), 
            .I3(n11_adj_4980), .O(n75376));
    defparam i59541_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33_adj_4984), 
            .I3(GND_net), .O(n12_adj_4989));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_4981), 
            .I3(GND_net), .O(n10_adj_4990));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_4989), .I1(n233[17]), .I2(n35_adj_4979), 
            .I3(GND_net), .O(n30_adj_4991));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i60498_4_lut (.I0(n13_adj_4981), .I1(n11_adj_4980), .I2(n9_adj_4985), 
            .I3(n75406), .O(n76333));
    defparam i60498_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i60488_4_lut (.I0(n19_adj_4987), .I1(n17_adj_4986), .I2(n15_adj_4982), 
            .I3(n76333), .O(n76323));
    defparam i60488_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i61536_4_lut (.I0(n25_adj_4978), .I1(n23_adj_4977), .I2(n21_adj_4988), 
            .I3(n76323), .O(n77371));
    defparam i61536_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i60925_4_lut (.I0(n31_adj_4976), .I1(n29_adj_4975), .I2(n27_adj_4983), 
            .I3(n77371), .O(n76760));
    defparam i60925_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i61664_4_lut (.I0(n37_adj_4974), .I1(n35_adj_4979), .I2(n33_adj_4984), 
            .I3(n76760), .O(n77499));
    defparam i61664_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43_adj_4973), 
            .I3(GND_net), .O(n16_adj_4992));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61266_3_lut (.I0(n6_adj_4937), .I1(n247), .I2(n21_adj_4988), 
            .I3(GND_net), .O(n77101));   // verilog/motorControl.v(56[14:36])
    defparam i61266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61267_3_lut (.I0(n77101), .I1(n233[11]), .I2(n23_adj_4977), 
            .I3(GND_net), .O(n77102));   // verilog/motorControl.v(56[14:36])
    defparam i61267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43903_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n62), 
            .I3(GND_net), .O(n20370[0]));   // verilog/motorControl.v(61[20:26])
    defparam i43903_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_4986), 
            .I3(GND_net), .O(n8_adj_4993));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4992), .I1(n233[22]), .I2(n45_adj_4972), 
            .I3(GND_net), .O(n24_adj_4994));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59511_4_lut (.I0(n43_adj_4973), .I1(n25_adj_4978), .I2(n23_adj_4977), 
            .I3(n75388), .O(n75346));
    defparam i59511_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61067_4_lut (.I0(n24_adj_4994), .I1(n8_adj_4993), .I2(n45_adj_4972), 
            .I3(n75342), .O(n76902));   // verilog/motorControl.v(56[14:36])
    defparam i61067_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59984_3_lut (.I0(n77102), .I1(n233[12]), .I2(n25_adj_4978), 
            .I3(GND_net), .O(n75819));   // verilog/motorControl.v(56[14:36])
    defparam i59984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4995));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i61264_3_lut (.I0(n4_adj_4995), .I1(n233[13]), .I2(n27_adj_4983), 
            .I3(GND_net), .O(n77099));   // verilog/motorControl.v(56[14:36])
    defparam i61264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61265_3_lut (.I0(n77099), .I1(n233[14]), .I2(n29_adj_4975), 
            .I3(GND_net), .O(n77100));   // verilog/motorControl.v(56[14:36])
    defparam i61265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59535_4_lut (.I0(n33_adj_4984), .I1(n31_adj_4976), .I2(n29_adj_4975), 
            .I3(n75376), .O(n75370));
    defparam i59535_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61614_4_lut (.I0(n30_adj_4991), .I1(n10_adj_4990), .I2(n35_adj_4979), 
            .I3(n75364), .O(n77449));   // verilog/motorControl.v(56[14:36])
    defparam i61614_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i59986_3_lut (.I0(n77100), .I1(n233[15]), .I2(n31_adj_4976), 
            .I3(GND_net), .O(n75821));   // verilog/motorControl.v(56[14:36])
    defparam i59986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61756_4_lut (.I0(n75821), .I1(n77449), .I2(n35_adj_4979), 
            .I3(n75370), .O(n77591));   // verilog/motorControl.v(56[14:36])
    defparam i61756_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut_4_lut_adj_962 (.I0(\Kp[1] ), .I1(n207[22]), .I2(n62), 
            .I3(n70879), .O(n20370[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut_adj_962.LUT_INIT = 16'h7f80;
    SB_LUT4 i61757_3_lut (.I0(n77591), .I1(n239), .I2(n37_adj_4974), .I3(GND_net), 
            .O(n77592));   // verilog/motorControl.v(56[14:36])
    defparam i61757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61720_3_lut (.I0(n77592), .I1(n233[19]), .I2(n39_adj_4971), 
            .I3(GND_net), .O(n77555));   // verilog/motorControl.v(56[14:36])
    defparam i61720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i59515_4_lut (.I0(n43_adj_4973), .I1(n41_adj_4970), .I2(n39_adj_4971), 
            .I3(n77499), .O(n75350));
    defparam i59515_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i61578_4_lut (.I0(n75819), .I1(n76902), .I2(n45_adj_4972), 
            .I3(n75346), .O(n77413));   // verilog/motorControl.v(56[14:36])
    defparam i61578_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i59992_3_lut (.I0(n77555), .I1(n233[20]), .I2(n41_adj_4970), 
            .I3(GND_net), .O(n75827));   // verilog/motorControl.v(56[14:36])
    defparam i59992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i61580_4_lut (.I0(n75827), .I1(n77413), .I2(n45_adj_4972), 
            .I3(n75350), .O(n77415));   // verilog/motorControl.v(56[14:36])
    defparam i61580_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i61581_3_lut (.I0(n77415), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i61581_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n359));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n359), .I2(GND_net), .I3(GND_net), 
            .O(n46[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4655));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4654));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4653));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4996[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4652));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4651));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4650));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4649));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4648));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4647));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4646));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n11880_bdd_4_lut_62943 (.I0(n11880), .I1(n74624), .I2(setpoint[14]), 
            .I3(n4734), .O(n78813));
    defparam n11880_bdd_4_lut_62943.LUT_INIT = 16'he4aa;
    SB_LUT4 n78813_bdd_4_lut (.I0(n78813), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4734), .O(n78816));
    defparam n78813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4645));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    
endmodule
