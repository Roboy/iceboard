// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Jan 28 16:13:57 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    output SCL;   // verilog/TinyFPGA_B.v(21[10:13])
    input SDA /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, CLK_c, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(42[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(88[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(89[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(123[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n4;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n29529, n29519, n29517, n29513, n29511;
    wire [31:0]motor_state_23__N_50;
    wire [23:0]displacement_23__N_26;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n4_adj_4466, n29936, n15010, n7410, n4169, n29802, n7, 
        n30906, n4167, n15009, n15008, n15007, n15006, n15005, 
        n15004, n15003, n15002, n15001, n15000, n14999, n14998, 
        n14997, n14996, n14995, n14994, n14993, n14992, n14991, 
        n14990, n14989, n14988, n14987, n14986, n14985, n14984, 
        n14983, n14982, n14981, n21995, n21980, n14980, n14979, 
        n14978, n14977, n14976;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n15, n15_adj_4467, n3, n4_adj_4468, n5, n6, n7_adj_4469, 
        n8, n9, n10, n11, n12, n13, n14, n15_adj_4470, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n21994, n21993, n7330;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire n21979, tx_active, n21978, n21977, n123, n21992;
    wire [31:0]\FRAME_MATCHER.state_31__N_2380 ;
    
    wire n30136, n14975, n14974, n14973, n14972, n14971, n1554, 
        n21991, n21990, n21976, n30064, n29704, n29702, n21989, 
        n21975, n21974, n21988, n21981, n18503, n21987, n21985, 
        n21986, n21984, n21983, n21982, n22106, n22105, n22104, 
        n22103, n22102, n22101, n22100, n22099, n13620, n13652, 
        n22098, n22097, n30253, n4_adj_4471, n22096, n30134, n10_adj_4472, 
        n3303, n22095;
    wire [31:0]\FRAME_MATCHER.state_31__N_2508 ;
    
    wire n22094, n22093, n22092, n22091, n52, n22090;
    wire [31:0]\FRAME_MATCHER.state_31__N_2540 ;
    
    wire n20610, n22089, n22088, n22087, n22086, n22085, n22084, 
        n107, n15476, n15475, n15474, n15473, n15472, n15471, 
        n15470, n15469, n15468, n15467, n15466, n15465, n15464, 
        n15463, n15462, n15461, n15460, n15459, n15458, n15457, 
        n15456, n15455, n15454, n15453, n15452, n15451, n15450, 
        n15449, n15448, n15447, n15446, n15442, n15441, n15436, 
        n15435, n15434, n15433, n15432, n15431, n15430, n15429, 
        n15428, n15427, n15426, n15425, n15424, n15423, n15422, 
        n15421, n15420, n15419, n15418, n15417, n15416, n15415, 
        n15414, n15413, n15412, n15411, n15410, n15409, n15408, 
        n15407, n14970, n14969, n29290, n63, n29288, n29975, n63_adj_4473, 
        n27693, n30923, n14_adj_4474, n15231, n15230, n15229, n15228, 
        n15227, n15226, n30135, n15225, n15224, n15223, quadA_debounced, 
        quadB_debounced, n10_adj_4475, quadA_debounced_adj_4476, quadB_debounced_adj_4477, 
        n15222, n15221, n15220, n15219, n15218, n15217, n15216, 
        n15215, n15214, n15213, n15212, n15211, n15210, n15209, 
        n15208, n15207, n29911, n15206, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n15205, n13483, n5_adj_4478, n14968, n15204, n15203, n15202, 
        n15201, n15200, n15199, n15198, n4_adj_4479, n3_adj_4480, 
        n15197;
    wire [2:0]r_SM_Main_2__N_3262;
    
    wire n15196, n15195, n15194, n15193, n15192, n15191, n15190, 
        n15189, n15188, n15187, n15186, n15185, n15184, n15183, 
        n15182;
    wire [2:0]r_SM_Main_adj_4574;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_4576;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3333;
    
    wire n15181, n15180, n15179, n15178, n15177, n15176, n15175, 
        n15174, n15173, n15172, n15171, n15170, n15169, n15168, 
        n15167, n15166, n15165, n15164, n15163, n15162, n15161, 
        n15160, n15159, n15158, n2;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15157, n15156, n15155, n15154, n15153, n15152, n15151, 
        n15150;
    wire [1:0]reg_B_adj_4587;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n15149, n15148, n15147, n15146, n15145, n14794, n15144, 
        n15143, n15142, n15141, n15140, n15139, n15138, n15137, 
        n15136, n15135, n15134, n15133, n15132, n15131, n15130, 
        n15129, n15128, n15127, n15126, n15125, n15124, n15123, 
        n15122, n15121, n15120, n15119, n15118, n15117, n15116, 
        n15115, n15114, n15113, n15112, n15111, n14744, n15110, 
        n15109, n15108, n15107, n4_adj_4487, n15106, n15105, n15104, 
        n15103, n15102, n15101, n6_adj_4488, n7_adj_4489, n8_adj_4490, 
        n9_adj_4491, n10_adj_4492, n11_adj_4493, n12_adj_4494, n13_adj_4495, 
        n14_adj_4496, n15_adj_4497, n16_adj_4498, n17_adj_4499, n18_adj_4500, 
        n19_adj_4501, n20_adj_4502, n21_adj_4503, n22_adj_4504, n23_adj_4505, 
        n24_adj_4506, n25_adj_4507, n15100, n14964, n29913, n15099, 
        n15098, n13646, n4_adj_4508, n6_adj_4509, n7_adj_4510, n8_adj_4511, 
        n9_adj_4512, n10_adj_4513, n11_adj_4514, n12_adj_4515, n13_adj_4516, 
        n15_adj_4517, n17_adj_4518, n19_adj_4519, n21_adj_4520, n29935, 
        n23_adj_4521, n25_adj_4522, n27, n29, n30, n31, n33, n35, 
        n29934, n30062, n7_adj_4523, n26830, n26810, n14921, n26721, 
        n15097, n15096, n15095, n15094, n15093, n15092, n15091, 
        n15090, n15089, n15088, n15087, n15086, n15085, n15084, 
        n15083, n15082, n15081, n15080, n15079, n15078, n15077, 
        n15076, n15075, n15074, n15073, n15072, n15071, n15070, 
        n15069, n15068, n15067, n15066, n26676, n15065, n15064, 
        n15063, n15062, n15061, n15060, n15059, n15058, n15057, 
        n15056, n15055, n15054, n15053, n15052, n15051, n15050, 
        n15049, n15048, n15047, n15046, n15045, n15044, n15043, 
        n15042, n14961, n14958, n14957, n14956, n15041, n15040, 
        n15039, n15038, n15037, n15036, n15035, n15034, n14955, 
        n14954, n14953, n14952, n14950, n14949, n14948, n14947, 
        n15033, n15032, n15031, n15030, n15029, n15028, n15027, 
        n15026, n15025, n15024, n15023, n15022, n15021, n15020, 
        n15019, n15018, n15017, n15016, n15015, n15014, n15013, 
        n15012, n15011, n13618, n13615, n30113, n30063, n25972, 
        n30021, n30018, n29867, n14946, n14945, n6_adj_4524, n30907, 
        n29792, n27279, n14941, n6_adj_4525, n28252, n25630, n13657, 
        n4_adj_4526, n13493, n7480, n24720, n10927, n29933, n6_adj_4527, 
        n13481;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced, 
            quadB_debounced}), .n28252(n28252), .reg_B({reg_B}), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .VCC_net(VCC_net), .n15441(n15441), .n14954(n14954), .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_LUT4 i11351_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n10927), .I3(GND_net), .O(n15182));   // verilog/coms.v(127[12] 300[6])
    defparam i11351_3_lut.LUT_INIT = 16'hcaca;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_26 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF h2_25 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i11352_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n10927), .I3(GND_net), .O(n15183));   // verilog/coms.v(127[12] 300[6])
    defparam i11352_3_lut.LUT_INIT = 16'hcaca;
    neopixel nx (.\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .timer({timer}), .VCC_net(VCC_net), .start(start), 
            .\state[0] (state[0]), .\state[1] (state[1]), .n4(n4_adj_4526), 
            .n20610(n20610), .n107(n107), .n26721(n26721), .n27279(n27279), 
            .n1554(n1554), .neopxl_color({neopxl_color}), .n14958(n14958), 
            .n15476(n15476), .n15475(n15475), .n15474(n15474), .n15473(n15473), 
            .n15472(n15472), .n15471(n15471), .n15470(n15470), .n15469(n15469), 
            .n15468(n15468), .n15467(n15467), .n15466(n15466), .n15465(n15465), 
            .n15464(n15464), .n15463(n15463), .n15462(n15462), .n15461(n15461), 
            .n15460(n15460), .n15459(n15459), .n15458(n15458), .n15457(n15457), 
            .n15456(n15456), .n15455(n15455), .n15454(n15454), .n15453(n15453), 
            .n15452(n15452), .n15451(n15451), .n15450(n15450), .n15449(n15449), 
            .n15448(n15448), .n15447(n15447), .n15446(n15446), .n24720(n24720), 
            .LED_c(LED_c), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(44[10] 50[2])
    SB_LUT4 i11353_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n10927), .I3(GND_net), .O(n15184));   // verilog/coms.v(127[12] 300[6])
    defparam i11353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_4472));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4472), .I2(control_mode[2]), 
            .I3(GND_net), .O(n13646));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11354_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n10927), .I3(GND_net), .O(n15185));   // verilog/coms.v(127[12] 300[6])
    defparam i11354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11355_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n10927), .I3(GND_net), .O(n15186));   // verilog/coms.v(127[12] 300[6])
    defparam i11355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n13493), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n13646), 
            .I3(GND_net), .O(n15_adj_4467));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i11356_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n10927), .I3(GND_net), .O(n15187));   // verilog/coms.v(127[12] 300[6])
    defparam i11356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11357_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n10927), .I3(GND_net), .O(n15188));   // verilog/coms.v(127[12] 300[6])
    defparam i11357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4507));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11358_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n10927), .I3(GND_net), .O(n15189));   // verilog/coms.v(127[12] 300[6])
    defparam i11358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11359_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n10927), .I3(GND_net), .O(n15190));   // verilog/coms.v(127[12] 300[6])
    defparam i11359_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dir_30 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i11360_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n10927), .I3(GND_net), .O(n15191));   // verilog/coms.v(127[12] 300[6])
    defparam i11360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11361_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n10927), .I3(GND_net), .O(n15192));   // verilog/coms.v(127[12] 300[6])
    defparam i11361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11362_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n10927), .I3(GND_net), .O(n15193));   // verilog/coms.v(127[12] 300[6])
    defparam i11362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11363_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n10927), .I3(GND_net), .O(n15194));   // verilog/coms.v(127[12] 300[6])
    defparam i11363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11364_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n10927), .I3(GND_net), .O(n15195));   // verilog/coms.v(127[12] 300[6])
    defparam i11364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11365_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n10927), .I3(GND_net), .O(n15196));   // verilog/coms.v(127[12] 300[6])
    defparam i11365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11366_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n10927), .I3(GND_net), .O(n15197));   // verilog/coms.v(127[12] 300[6])
    defparam i11366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11162_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4167), .I3(GND_net), .O(n14993));   // verilog/coms.v(127[12] 300[6])
    defparam i11162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11367_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n10927), .I3(GND_net), .O(n15198));   // verilog/coms.v(127[12] 300[6])
    defparam i11367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11368_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n10927), .I3(GND_net), .O(n15199));   // verilog/coms.v(127[12] 300[6])
    defparam i11368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11369_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n10927), .I3(GND_net), .O(n15200));   // verilog/coms.v(127[12] 300[6])
    defparam i11369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11370_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n10927), .I3(GND_net), .O(n15201));   // verilog/coms.v(127[12] 300[6])
    defparam i11370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11371_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n10927), .I3(GND_net), .O(n15202));   // verilog/coms.v(127[12] 300[6])
    defparam i11371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11372_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n10927), .I3(GND_net), .O(n15203));   // verilog/coms.v(127[12] 300[6])
    defparam i11372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11373_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n10927), .I3(GND_net), .O(n15204));   // verilog/coms.v(127[12] 300[6])
    defparam i11373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11374_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n10927), .I3(GND_net), .O(n15205));   // verilog/coms.v(127[12] 300[6])
    defparam i11374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11375_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n10927), .I3(GND_net), .O(n15206));   // verilog/coms.v(127[12] 300[6])
    defparam i11375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11376_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n10927), .I3(GND_net), .O(n15207));   // verilog/coms.v(127[12] 300[6])
    defparam i11376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11163_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4167), .I3(GND_net), .O(n14994));   // verilog/coms.v(127[12] 300[6])
    defparam i11163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11377_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n10927), .I3(GND_net), .O(n15208));   // verilog/coms.v(127[12] 300[6])
    defparam i11377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11378_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n4169), .I3(GND_net), .O(n15209));   // verilog/coms.v(127[12] 300[6])
    defparam i11378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11379_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n4169), .I3(GND_net), .O(n15210));   // verilog/coms.v(127[12] 300[6])
    defparam i11379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11380_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n4169), .I3(GND_net), .O(n15211));   // verilog/coms.v(127[12] 300[6])
    defparam i11380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11381_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n4169), .I3(GND_net), .O(n15212));   // verilog/coms.v(127[12] 300[6])
    defparam i11381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11382_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n4169), .I3(GND_net), .O(n15213));   // verilog/coms.v(127[12] 300[6])
    defparam i11382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11383_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n4169), .I3(GND_net), .O(n15214));   // verilog/coms.v(127[12] 300[6])
    defparam i11383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11384_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n4169), .I3(GND_net), .O(n15215));   // verilog/coms.v(127[12] 300[6])
    defparam i11384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11385_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n4169), .I3(GND_net), .O(n15216));   // verilog/coms.v(127[12] 300[6])
    defparam i11385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11386_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n4169), .I3(GND_net), .O(n15217));   // verilog/coms.v(127[12] 300[6])
    defparam i11386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11387_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n4169), .I3(GND_net), .O(n15218));   // verilog/coms.v(127[12] 300[6])
    defparam i11387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11388_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n4169), .I3(GND_net), .O(n15219));   // verilog/coms.v(127[12] 300[6])
    defparam i11388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11389_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n4169), .I3(GND_net), .O(n15220));   // verilog/coms.v(127[12] 300[6])
    defparam i11389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11390_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n4169), .I3(GND_net), .O(n15221));   // verilog/coms.v(127[12] 300[6])
    defparam i11390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11391_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n4169), .I3(GND_net), .O(n15222));   // verilog/coms.v(127[12] 300[6])
    defparam i11391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11392_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n4169), .I3(GND_net), .O(n15223));   // verilog/coms.v(127[12] 300[6])
    defparam i11392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11393_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n4169), .I3(GND_net), .O(n15224));   // verilog/coms.v(127[12] 300[6])
    defparam i11393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11394_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n4169), .I3(GND_net), .O(n15225));   // verilog/coms.v(127[12] 300[6])
    defparam i11394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11395_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n4169), .I3(GND_net), .O(n15226));   // verilog/coms.v(127[12] 300[6])
    defparam i11395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4506));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11396_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n4169), .I3(GND_net), .O(n15227));   // verilog/coms.v(127[12] 300[6])
    defparam i11396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11397_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n4169), .I3(GND_net), .O(n15228));   // verilog/coms.v(127[12] 300[6])
    defparam i11397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11398_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n4169), .I3(GND_net), .O(n15229));   // verilog/coms.v(127[12] 300[6])
    defparam i11398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11399_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n4169), .I3(GND_net), .O(n15230));   // verilog/coms.v(127[12] 300[6])
    defparam i11399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11400_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n4169), .I3(GND_net), .O(n15231));   // verilog/coms.v(127[12] 300[6])
    defparam i11400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4505));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4504));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4503));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4502));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4475));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[29]), .I2(pwm_counter[25]), 
            .I3(pwm_counter[26]), .O(n14_adj_4474));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[30]), .I1(n14_adj_4474), .I2(n10_adj_4475), 
            .I3(pwm_counter[24]), .O(n13481));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4501));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4500));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11161_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4167), .I3(GND_net), .O(n14992));   // verilog/coms.v(127[12] 300[6])
    defparam i11161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4499));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_37_i16_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[15]), 
            .I3(encoder0_position[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_38_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11175_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15006));   // verilog/coms.v(127[12] 300[6])
    defparam i11175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3262[2]), 
            .I3(r_SM_Main[0]), .O(n14744));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n14744), 
            .I3(rx_data_ready), .O(n25630));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i25131_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n25972));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i25131_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n2), .I3(n22106), .O(displacement_23__N_26[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4480), .I3(n22105), .O(displacement_23__N_26[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n22105), .I0(encoder1_position[22]), 
            .I1(n3_adj_4480), .CO(n22106));
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n4_adj_4479), .I3(n22104), .O(displacement_23__N_26[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n22104), .I0(encoder1_position[21]), 
            .I1(n4_adj_4479), .CO(n22105));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4478), .I3(n22103), .O(displacement_23__N_26[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n22103), .I0(encoder1_position[20]), 
            .I1(n5_adj_4478), .CO(n22104));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4488), .I3(n22102), .O(displacement_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n22102), .I0(encoder1_position[19]), 
            .I1(n6_adj_4488), .CO(n22103));
    SB_DFF h1_24 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4489), .I3(n22101), .O(displacement_23__N_26[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4469));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4498));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4497));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n22101), .I0(encoder1_position[18]), 
            .I1(n7_adj_4489), .CO(n22102));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4490), .I3(n22100), .O(displacement_23__N_26[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n22100), .I0(encoder1_position[17]), 
            .I1(n8_adj_4490), .CO(n22101));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4491), .I3(n22099), .O(displacement_23__N_26[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n22099), .I0(encoder1_position[16]), 
            .I1(n9_adj_4491), .CO(n22100));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4492), .I3(n22098), .O(displacement_23__N_26[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4496));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4495));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_485_24_lut (.I0(duty[22]), .I1(n30253), .I2(n3), .I3(n21995), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n22098), .I0(encoder1_position[15]), 
            .I1(n10_adj_4492), .CO(n22099));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4493), .I3(n22097), .O(displacement_23__N_26[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_485_23_lut (.I0(duty[21]), .I1(n30253), .I2(n4_adj_4468), 
            .I3(n21994), .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_23 (.CI(n21994), .I0(n30253), .I1(n4_adj_4468), .CO(n21995));
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n22097), .I0(encoder1_position[14]), 
            .I1(n11_adj_4493), .CO(n22098));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4494), .I3(n22096), .O(displacement_23__N_26[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4494));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4468));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n22096), .I0(encoder1_position[13]), 
            .I1(n12_adj_4494), .CO(n22097));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4493));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4495), .I3(n22095), .O(displacement_23__N_26[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n22095), .I0(encoder1_position[12]), 
            .I1(n13_adj_4495), .CO(n22096));
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4496), .I3(n22094), .O(displacement_23__N_26[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4492));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_26[23]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_LUT4 add_485_22_lut (.I0(duty[20]), .I1(n30253), .I2(n5), .I3(n21993), 
            .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4491));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n22094), .I0(encoder1_position[11]), 
            .I1(n14_adj_4496), .CO(n22095));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4490));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_485_22 (.CI(n21993), .I0(n30253), .I1(n5), .CO(n21994));
    SB_LUT4 add_485_21_lut (.I0(duty[19]), .I1(n30253), .I2(n6), .I3(n21992), 
            .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4497), .I3(n22093), .O(displacement_23__N_26[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_485_21 (.CI(n21992), .I0(n30253), .I1(n6), .CO(n21993));
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n22093), .I0(encoder1_position[10]), 
            .I1(n15_adj_4497), .CO(n22094));
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4498), .I3(n22092), .O(displacement_23__N_26[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_485_20_lut (.I0(duty[18]), .I1(n30253), .I2(n7_adj_4469), 
            .I3(n21991), .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4489));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4488));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4478));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_485_20 (.CI(n21991), .I0(n30253), .I1(n7_adj_4469), .CO(n21992));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4479));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11576_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4167), .I3(GND_net), .O(n15407));   // verilog/coms.v(127[12] 300[6])
    defparam i11576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11164_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4487), 
            .I3(n13657), .O(n14995));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11164_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11577_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4167), .I3(GND_net), .O(n15408));   // verilog/coms.v(127[12] 300[6])
    defparam i11577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11578_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4167), .I3(GND_net), .O(n15409));   // verilog/coms.v(127[12] 300[6])
    defparam i11578_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n22092), .I0(encoder1_position[9]), 
            .I1(n16_adj_4498), .CO(n22093));
    SB_LUT4 i11579_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4167), .I3(GND_net), .O(n15410));   // verilog/coms.v(127[12] 300[6])
    defparam i11579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4480));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(201[21:58])
    defparam encoder1_position_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_485_19_lut (.I0(duty[17]), .I1(n30253), .I2(n8), .I3(n21990), 
            .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4499), .I3(n22091), .O(displacement_23__N_26[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11165_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14996));   // verilog/coms.v(127[12] 300[6])
    defparam i11165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11166_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14997));   // verilog/coms.v(127[12] 300[6])
    defparam i11166_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_19 (.CI(n21990), .I0(n30253), .I1(n8), .CO(n21991));
    SB_LUT4 add_485_18_lut (.I0(duty[16]), .I1(n30253), .I2(n9), .I3(n21989), 
            .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11580_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4167), .I3(GND_net), .O(n15411));   // verilog/coms.v(127[12] 300[6])
    defparam i11580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n22091), .I0(encoder1_position[8]), 
            .I1(n17_adj_4499), .CO(n22092));
    SB_LUT4 i11581_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4167), .I3(GND_net), .O(n15412));   // verilog/coms.v(127[12] 300[6])
    defparam i11581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11582_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4167), .I3(GND_net), .O(n15413));   // verilog/coms.v(127[12] 300[6])
    defparam i11582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11583_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4167), .I3(GND_net), .O(n15414));   // verilog/coms.v(127[12] 300[6])
    defparam i11583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11584_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n4167), .I3(GND_net), .O(n15415));   // verilog/coms.v(127[12] 300[6])
    defparam i11584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11585_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4167), .I3(GND_net), .O(n15416));   // verilog/coms.v(127[12] 300[6])
    defparam i11585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4500), .I3(n22090), .O(displacement_23__N_26[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11586_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4167), .I3(GND_net), .O(n15417));   // verilog/coms.v(127[12] 300[6])
    defparam i11586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11587_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4167), .I3(GND_net), .O(n15418));   // verilog/coms.v(127[12] 300[6])
    defparam i11587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11588_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4167), .I3(GND_net), .O(n15419));   // verilog/coms.v(127[12] 300[6])
    defparam i11588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11589_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4167), .I3(GND_net), .O(n15420));   // verilog/coms.v(127[12] 300[6])
    defparam i11589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11590_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4167), .I3(GND_net), .O(n15421));   // verilog/coms.v(127[12] 300[6])
    defparam i11590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11591_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4167), .I3(GND_net), .O(n15422));   // verilog/coms.v(127[12] 300[6])
    defparam i11591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11592_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4167), .I3(GND_net), .O(n15423));   // verilog/coms.v(127[12] 300[6])
    defparam i11592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11593_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4167), .I3(GND_net), .O(n15424));   // verilog/coms.v(127[12] 300[6])
    defparam i11593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11594_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4167), .I3(GND_net), .O(n15425));   // verilog/coms.v(127[12] 300[6])
    defparam i11594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11595_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4167), .I3(GND_net), .O(n15426));   // verilog/coms.v(127[12] 300[6])
    defparam i11595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11596_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n4167), .I3(GND_net), .O(n15427));   // verilog/coms.v(127[12] 300[6])
    defparam i11596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11597_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4167), .I3(GND_net), .O(n15428));   // verilog/coms.v(127[12] 300[6])
    defparam i11597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11598_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4167), .I3(GND_net), .O(n15429));   // verilog/coms.v(127[12] 300[6])
    defparam i11598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11599_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4167), .I3(GND_net), .O(n15430));   // verilog/coms.v(127[12] 300[6])
    defparam i11599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11600_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4167), .I3(GND_net), .O(n15431));   // verilog/coms.v(127[12] 300[6])
    defparam i11600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11601_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4167), .I3(GND_net), .O(n15432));   // verilog/coms.v(127[12] 300[6])
    defparam i11601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11602_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4167), .I3(GND_net), .O(n15433));   // verilog/coms.v(127[12] 300[6])
    defparam i11602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11603_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4167), .I3(GND_net), .O(n15434));   // verilog/coms.v(127[12] 300[6])
    defparam i11603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11604_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4167), .I3(GND_net), .O(n15435));   // verilog/coms.v(127[12] 300[6])
    defparam i11604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11167_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14998));   // verilog/coms.v(127[12] 300[6])
    defparam i11167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11605_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4167), .I3(GND_net), .O(n15436));   // verilog/coms.v(127[12] 300[6])
    defparam i11605_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n22090), .I0(encoder1_position[7]), 
            .I1(n18_adj_4500), .CO(n22091));
    SB_LUT4 i1_4_lut (.I0(n123), .I1(n26676), .I2(n63), .I3(n6_adj_4527), 
            .O(n7_adj_4523));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'haf23;
    SB_LUT4 mux_37_i17_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[16]), 
            .I3(encoder0_position[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i2_4_lut (.I0(n7_adj_4523), .I1(n123), .I2(n13618), .I3(n7480), 
            .O(n6_adj_4524));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'haeaf;
    SB_LUT4 i3_4_lut (.I0(n63_adj_4473), .I1(n6_adj_4524), .I2(n13615), 
            .I3(\FRAME_MATCHER.state_31__N_2508 [1]), .O(n30907));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hdfdd;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_26[22]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n63_adj_4473), .I1(n13618), .I2(n7480), 
            .I3(n52), .O(n6_adj_4525));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'h7555;
    SB_LUT4 i2_4_lut_adj_1608 (.I0(\FRAME_MATCHER.state_31__N_2380 [2]), .I1(n3303), 
            .I2(n6_adj_4527), .I3(n13615), .O(n7));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1608.LUT_INIT = 16'ha0ee;
    SB_LUT4 i4_4_lut_adj_1609 (.I0(n7), .I1(\FRAME_MATCHER.state_31__N_2540 [2]), 
            .I2(n6_adj_4525), .I3(n13620), .O(n30906));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1609.LUT_INIT = 16'hfafe;
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4501), .I3(n22089), .O(displacement_23__N_26[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n22089), .I0(encoder1_position[6]), 
            .I1(n19_adj_4501), .CO(n22090));
    SB_LUT4 i24455_4_lut (.I0(n27279), .I1(n107), .I2(n26721), .I3(state[0]), 
            .O(n29290));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24455_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i18_4_lut (.I0(n29290), .I1(n29288), .I2(state[1]), .I3(n4_adj_4526), 
            .O(n24720));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i11610_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n28252), 
            .I3(GND_net), .O(n15441));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11610_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11611_3_lut (.I0(quadA_debounced_adj_4476), .I1(reg_B_adj_4587[1]), 
            .I2(n27693), .I3(GND_net), .O(n15442));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11611_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11133_3_lut (.I0(n14921), .I1(r_Bit_Index[0]), .I2(n14794), 
            .I3(GND_net), .O(n14964));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11133_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i11130_3_lut (.I0(n26830), .I1(r_Bit_Index_adj_4576[0]), .I2(n26810), 
            .I3(GND_net), .O(n14961));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11130_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i11615_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n1554), .I3(GND_net), .O(n15446));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11616_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n1554), .I3(GND_net), .O(n15447));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11617_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n1554), .I3(GND_net), .O(n15448));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11618_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n1554), .I3(GND_net), .O(n15449));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11619_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n1554), .I3(GND_net), .O(n15450));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11620_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n1554), .I3(GND_net), .O(n15451));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11621_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n1554), .I3(GND_net), .O(n15452));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11622_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n1554), .I3(GND_net), .O(n15453));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11623_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n1554), .I3(GND_net), .O(n15454));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11624_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n1554), .I3(GND_net), .O(n15455));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11625_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n1554), .I3(GND_net), .O(n15456));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11626_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n1554), .I3(GND_net), .O(n15457));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11627_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n1554), .I3(GND_net), .O(n15458));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11628_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n1554), .I3(GND_net), .O(n15459));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11629_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n1554), .I3(GND_net), .O(n15460));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11630_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n1554), .I3(GND_net), .O(n15461));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11630_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_26[21]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_26[20]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_26[19]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_26[18]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_26[17]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_26[16]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_26[15]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_26[14]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_26[13]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_26[12]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_26[11]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_26[10]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_26[9]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_26[8]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_26[7]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_26[6]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_26[5]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_26[4]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_26[3]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_26[2]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_26[1]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(97[10] 110[6])
    SB_LUT4 i11176_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15007));   // verilog/coms.v(127[12] 300[6])
    defparam i11176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11177_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15008));   // verilog/coms.v(127[12] 300[6])
    defparam i11177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11631_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n1554), .I3(GND_net), .O(n15462));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4502), .I3(n22088), .O(displacement_23__N_26[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11632_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n1554), .I3(GND_net), .O(n15463));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11633_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n1554), .I3(GND_net), .O(n15464));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11633_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_18 (.CI(n21989), .I0(n30253), .I1(n9), .CO(n21990));
    SB_LUT4 i11634_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n1554), .I3(GND_net), .O(n15465));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11635_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n1554), .I3(GND_net), .O(n15466));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11635_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n22088), .I0(encoder1_position[5]), 
            .I1(n20_adj_4502), .CO(n22089));
    SB_LUT4 i11636_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n1554), .I3(GND_net), .O(n15467));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_485_17_lut (.I0(duty[15]), .I1(n30253), .I2(n10), .I3(n21988), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11637_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n1554), .I3(GND_net), .O(n15468));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4503), .I3(n22087), .O(displacement_23__N_26[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11638_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n1554), .I3(GND_net), .O(n15469));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11639_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n1554), .I3(GND_net), .O(n15470));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11639_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n22087), .I0(encoder1_position[4]), 
            .I1(n21_adj_4503), .CO(n22088));
    SB_LUT4 i11640_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n1554), .I3(GND_net), .O(n15471));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4504), .I3(n22086), .O(displacement_23__N_26[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11641_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n1554), .I3(GND_net), .O(n15472));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11642_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n1554), .I3(GND_net), .O(n15473));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11642_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n22086), .I0(encoder1_position[3]), 
            .I1(n22_adj_4504), .CO(n22087));
    SB_LUT4 mux_37_i18_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[17]), 
            .I3(encoder0_position[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11643_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n1554), .I3(GND_net), .O(n15474));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11644_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n1554), .I3(GND_net), .O(n15475));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11644_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_17 (.CI(n21988), .I0(n30253), .I1(n10), .CO(n21989));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4505), .I3(n22085), .O(displacement_23__N_26[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n22085), .I0(encoder1_position[2]), 
            .I1(n23_adj_4505), .CO(n22086));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4506), .I3(n22084), .O(displacement_23__N_26[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n22084), .I0(encoder1_position[1]), 
            .I1(n24_adj_4506), .CO(n22085));
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_485_16_lut (.I0(duty[14]), .I1(n30253), .I2(n11), .I3(n21987), 
            .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4507), .I3(VCC_net), .O(displacement_23__N_26[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_485_16 (.CI(n21987), .I0(n30253), .I1(n11), .CO(n21988));
    SB_LUT4 add_485_15_lut (.I0(duty[13]), .I1(n30253), .I2(n12), .I3(n21986), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11168_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14999));   // verilog/coms.v(127[12] 300[6])
    defparam i11168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11169_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15000));   // verilog/coms.v(127[12] 300[6])
    defparam i11169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11170_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15001));   // verilog/coms.v(127[12] 300[6])
    defparam i11170_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4507), .CO(n22084));
    SB_LUT4 mux_37_i24_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[23]), 
            .I3(encoder0_position[23]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_38_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_38_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_485_15 (.CI(n21986), .I0(n30253), .I1(n12), .CO(n21987));
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_485_14_lut (.I0(duty[12]), .I1(n30253), .I2(n13), .I3(n21985), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i11171_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15002));   // verilog/coms.v(127[12] 300[6])
    defparam i11171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11172_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15003));   // verilog/coms.v(127[12] 300[6])
    defparam i11172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11173_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15004));   // verilog/coms.v(127[12] 300[6])
    defparam i11173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11645_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n1554), .I3(GND_net), .O(n15476));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11174_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15005));   // verilog/coms.v(127[12] 300[6])
    defparam i11174_3_lut.LUT_INIT = 16'hcaca;
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO SCL_pad (.PACKAGE_PIN(SCL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam SCL_pad.PIN_TYPE = 6'b011001;
    defparam SCL_pad.PULLUP = 1'b0;
    defparam SCL_pad.NEG_TRIGGER = 1'b0;
    defparam SCL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 mux_38_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_37_i19_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[18]), 
            .I3(encoder0_position[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11126_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n13657), 
            .O(n14957));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11126_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11127_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n1554), .I3(GND_net), .O(n14958));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11137_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4487), 
            .I3(n13652), .O(n14968));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11137_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11138_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n13652), 
            .O(n14969));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11138_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11139_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4466), 
            .I3(n13657), .O(n14970));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11139_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11140_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4466), 
            .I3(n13652), .O(n14971));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11140_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11141_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4167), .I3(GND_net), .O(n14972));   // verilog/coms.v(127[12] 300[6])
    defparam i11141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11142_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4167), .I3(GND_net), .O(n14973));   // verilog/coms.v(127[12] 300[6])
    defparam i11142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11143_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4167), .I3(GND_net), .O(n14974));   // verilog/coms.v(127[12] 300[6])
    defparam i11143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11144_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4167), .I3(GND_net), .O(n14975));   // verilog/coms.v(127[12] 300[6])
    defparam i11144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11145_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4167), .I3(GND_net), .O(n14976));   // verilog/coms.v(127[12] 300[6])
    defparam i11145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11146_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4167), .I3(GND_net), .O(n14977));   // verilog/coms.v(127[12] 300[6])
    defparam i11146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11147_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4167), .I3(GND_net), .O(n14978));   // verilog/coms.v(127[12] 300[6])
    defparam i11147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11148_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4167), .I3(GND_net), .O(n14979));   // verilog/coms.v(127[12] 300[6])
    defparam i11148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11149_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4167), .I3(GND_net), .O(n14980));   // verilog/coms.v(127[12] 300[6])
    defparam i11149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11150_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4167), .I3(GND_net), .O(n14981));   // verilog/coms.v(127[12] 300[6])
    defparam i11150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11151_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4167), .I3(GND_net), .O(n14982));   // verilog/coms.v(127[12] 300[6])
    defparam i11151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11152_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4167), .I3(GND_net), .O(n14983));   // verilog/coms.v(127[12] 300[6])
    defparam i11152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11153_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4167), .I3(GND_net), .O(n14984));   // verilog/coms.v(127[12] 300[6])
    defparam i11153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11154_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4167), .I3(GND_net), .O(n14985));   // verilog/coms.v(127[12] 300[6])
    defparam i11154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11155_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4167), .I3(GND_net), .O(n14986));   // verilog/coms.v(127[12] 300[6])
    defparam i11155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11156_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4167), .I3(GND_net), .O(n14987));   // verilog/coms.v(127[12] 300[6])
    defparam i11156_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_14 (.CI(n21985), .I0(n30253), .I1(n13), .CO(n21986));
    SB_LUT4 mux_38_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_37_i20_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[19]), 
            .I3(encoder0_position[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_4574[1]), .I1(r_SM_Main_adj_4574[0]), 
            .I2(r_SM_Main_adj_4574[2]), .I3(r_SM_Main_2__N_3333[1]), .O(n30923));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 mux_38_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11157_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4167), .I3(GND_net), .O(n14988));   // verilog/coms.v(127[12] 300[6])
    defparam i11157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11158_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4167), .I3(GND_net), .O(n14989));   // verilog/coms.v(127[12] 300[6])
    defparam i11158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11159_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4167), .I3(GND_net), .O(n14990));   // verilog/coms.v(127[12] 300[6])
    defparam i11159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_557_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4509));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11160_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4167), .I3(GND_net), .O(n14991));   // verilog/coms.v(127[12] 300[6])
    defparam i11160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_485_13_lut (.I0(duty[11]), .I1(n30253), .I2(n14), .I3(n21984), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_38_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_557_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4513));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i24421_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n29511));
    defparam i24421_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_485_13 (.CI(n21984), .I0(n30253), .I1(n14), .CO(n21985));
    SB_LUT4 add_485_12_lut (.I0(duty[10]), .I1(n30253), .I2(n15_adj_4470), 
            .I3(n21983), .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_38_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_557_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4515));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_485_12 (.CI(n21983), .I0(n30253), .I1(n15_adj_4470), 
            .CO(n21984));
    SB_LUT4 add_485_11_lut (.I0(duty[9]), .I1(n30253), .I2(n16), .I3(n21982), 
            .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_11 (.CI(n21982), .I0(n30253), .I1(n16), .CO(n21983));
    SB_LUT4 mux_38_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_485_10_lut (.I0(duty[8]), .I1(n30253), .I2(n17), .I3(n21981), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_557_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4511));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24439_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n29529));
    defparam i24439_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_485_10 (.CI(n21981), .I0(n30253), .I1(n17), .CO(n21982));
    SB_LUT4 add_485_9_lut (.I0(duty[7]), .I1(n30253), .I2(n18), .I3(n21980), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_9 (.CI(n21980), .I0(n30253), .I1(n18), .CO(n21981));
    SB_LUT4 add_485_8_lut (.I0(duty[6]), .I1(n30253), .I2(n19), .I3(n21979), 
            .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_8 (.CI(n21979), .I0(n30253), .I1(n19), .CO(n21980));
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_485_7_lut (.I0(duty[5]), .I1(n30253), .I2(n20), .I3(n21978), 
            .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_38_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11178_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15009));   // verilog/coms.v(127[12] 300[6])
    defparam i11178_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_7 (.CI(n21978), .I0(n30253), .I1(n20), .CO(n21979));
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_38_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_485_6_lut (.I0(duty[4]), .I1(n30253), .I2(n21), .I3(n21977), 
            .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_6 (.CI(n21977), .I0(n30253), .I1(n21), .CO(n21978));
    SB_LUT4 add_485_5_lut (.I0(duty[3]), .I1(n30253), .I2(n22), .I3(n21976), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_5 (.CI(n21976), .I0(n30253), .I1(n22), .CO(n21977));
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4470));   // verilog/TinyFPGA_B.v(107[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_485_4_lut (.I0(duty[2]), .I1(n30253), .I2(n23), .I3(n21975), 
            .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_37_i21_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[20]), 
            .I3(encoder0_position[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i22_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[21]), 
            .I3(encoder0_position[21]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i23_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[22]), 
            .I3(encoder0_position[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_38_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_557_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4512));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4514));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4518));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_485_4 (.CI(n21975), .I0(n30253), .I1(n23), .CO(n21976));
    SB_LUT4 LessThan_557_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4517));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4516));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_485_3_lut (.I0(duty[1]), .I1(n30253), .I2(n24), .I3(n21974), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_485_3 (.CI(n21974), .I0(n30253), .I1(n24), .CO(n21975));
    SB_LUT4 mux_38_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_557_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4510));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4520));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4521));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4519));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_557_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4522));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_485_2_lut (.I0(duty[0]), .I1(n30253), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_485_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_557_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11179_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15010));   // verilog/coms.v(127[12] 300[6])
    defparam i11179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1610 (.I0(n13481), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n13483));
    defparam i1_2_lut_adj_1610.LUT_INIT = 16'heeee;
    SB_LUT4 i24427_4_lut (.I0(n27), .I1(n15_adj_4517), .I2(n13_adj_4516), 
            .I3(n11_adj_4514), .O(n29517));
    defparam i24427_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24710_4_lut (.I0(n9_adj_4512), .I1(n7_adj_4510), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n29802));
    defparam i24710_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i11180_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15011));   // verilog/coms.v(127[12] 300[6])
    defparam i11180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24821_4_lut (.I0(n15_adj_4517), .I1(n13_adj_4516), .I2(n11_adj_4514), 
            .I3(n29802), .O(n29913));
    defparam i24821_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i11181_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15012));   // verilog/coms.v(127[12] 300[6])
    defparam i11181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11182_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15013));   // verilog/coms.v(127[12] 300[6])
    defparam i11182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11183_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15014));   // verilog/coms.v(127[12] 300[6])
    defparam i11183_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_485_2 (.CI(VCC_net), .I0(n30253), .I1(n25), .CO(n21974));
    SB_LUT4 i11184_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15015));   // verilog/coms.v(127[12] 300[6])
    defparam i11184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11185_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15016));   // verilog/coms.v(127[12] 300[6])
    defparam i11185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11186_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15017));   // verilog/coms.v(127[12] 300[6])
    defparam i11186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24819_4_lut (.I0(n21_adj_4520), .I1(n19_adj_4519), .I2(n17_adj_4518), 
            .I3(n29913), .O(n29911));
    defparam i24819_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24429_4_lut (.I0(n27), .I1(n25_adj_4522), .I2(n23_adj_4521), 
            .I3(n29911), .O(n29519));
    defparam i24429_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_557_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4508));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i24841_3_lut (.I0(n4_adj_4508), .I1(pwm_setpoint[13]), .I2(n27), 
            .I3(GND_net), .O(n29933));   // verilog/pwm.v(21[8:24])
    defparam i24841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11187_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15018));   // verilog/coms.v(127[12] 300[6])
    defparam i11187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_557_i30_3_lut (.I0(n12_adj_4515), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam LessThan_557_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24842_3_lut (.I0(n29933), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n29934));   // verilog/pwm.v(21[8:24])
    defparam i24842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24423_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n29517), 
            .O(n29513));
    defparam i24423_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24972_4_lut (.I0(n30), .I1(n10_adj_4513), .I2(n35), .I3(n29511), 
            .O(n30064));   // verilog/pwm.v(21[8:24])
    defparam i24972_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24612_3_lut (.I0(n29934), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n29704));   // verilog/pwm.v(21[8:24])
    defparam i24612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24843_3_lut (.I0(n6_adj_4509), .I1(pwm_setpoint[10]), .I2(n21_adj_4520), 
            .I3(GND_net), .O(n29935));   // verilog/pwm.v(21[8:24])
    defparam i24843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24844_3_lut (.I0(n29935), .I1(pwm_setpoint[11]), .I2(n23_adj_4521), 
            .I3(GND_net), .O(n29936));   // verilog/pwm.v(21[8:24])
    defparam i24844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24700_4_lut (.I0(n23_adj_4521), .I1(n21_adj_4520), .I2(n19_adj_4519), 
            .I3(n29529), .O(n29792));
    defparam i24700_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24775_3_lut (.I0(n8_adj_4511), .I1(pwm_setpoint[9]), .I2(n19_adj_4519), 
            .I3(GND_net), .O(n29867));   // verilog/pwm.v(21[8:24])
    defparam i24775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24610_3_lut (.I0(n29936), .I1(pwm_setpoint[12]), .I2(n25_adj_4522), 
            .I3(GND_net), .O(n29702));   // verilog/pwm.v(21[8:24])
    defparam i24610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24883_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n29519), 
            .O(n29975));
    defparam i24883_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25021_4_lut (.I0(n29704), .I1(n30064), .I2(n35), .I3(n29513), 
            .O(n30113));   // verilog/pwm.v(21[8:24])
    defparam i25021_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24926_4_lut (.I0(n29702), .I1(n29867), .I2(n25_adj_4522), 
            .I3(n29792), .O(n30018));   // verilog/pwm.v(21[8:24])
    defparam i24926_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i25043_4_lut (.I0(n30018), .I1(n30113), .I2(n35), .I3(n29975), 
            .O(n30135));   // verilog/pwm.v(21[8:24])
    defparam i25043_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i11188_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15019));   // verilog/coms.v(127[12] 300[6])
    defparam i11188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25044_3_lut (.I0(n30135), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n30136));   // verilog/pwm.v(21[8:24])
    defparam i25044_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25042_3_lut (.I0(n30136), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n30134));   // verilog/pwm.v(21[8:24])
    defparam i25042_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11189_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15020));   // verilog/coms.v(127[12] 300[6])
    defparam i11189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11190_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15021));   // verilog/coms.v(127[12] 300[6])
    defparam i11190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11191_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15022));   // verilog/coms.v(127[12] 300[6])
    defparam i11191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11192_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15023));   // verilog/coms.v(127[12] 300[6])
    defparam i11192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11193_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15024));   // verilog/coms.v(127[12] 300[6])
    defparam i11193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11194_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15025));   // verilog/coms.v(127[12] 300[6])
    defparam i11194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11195_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n15026));   // verilog/coms.v(127[12] 300[6])
    defparam i11195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11196_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n7330), 
            .I3(GND_net), .O(n15027));   // verilog/coms.v(127[12] 300[6])
    defparam i11196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11197_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n7330), 
            .I3(GND_net), .O(n15028));   // verilog/coms.v(127[12] 300[6])
    defparam i11197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11198_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n7330), 
            .I3(GND_net), .O(n15029));   // verilog/coms.v(127[12] 300[6])
    defparam i11198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11199_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n7330), 
            .I3(GND_net), .O(n15030));   // verilog/coms.v(127[12] 300[6])
    defparam i11199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11200_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n7330), 
            .I3(GND_net), .O(n15031));   // verilog/coms.v(127[12] 300[6])
    defparam i11200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11201_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n7330), 
            .I3(GND_net), .O(n15032));   // verilog/coms.v(127[12] 300[6])
    defparam i11201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11202_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n7330), 
            .I3(GND_net), .O(n15033));   // verilog/coms.v(127[12] 300[6])
    defparam i11202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11203_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n7330), 
            .I3(GND_net), .O(n15034));   // verilog/coms.v(127[12] 300[6])
    defparam i11203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11204_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n7330), 
            .I3(GND_net), .O(n15035));   // verilog/coms.v(127[12] 300[6])
    defparam i11204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11205_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n7330), 
            .I3(GND_net), .O(n15036));   // verilog/coms.v(127[12] 300[6])
    defparam i11205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11206_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n7330), 
            .I3(GND_net), .O(n15037));   // verilog/coms.v(127[12] 300[6])
    defparam i11206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11207_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n7330), 
            .I3(GND_net), .O(n15038));   // verilog/coms.v(127[12] 300[6])
    defparam i11207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11208_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n7330), 
            .I3(GND_net), .O(n15039));   // verilog/coms.v(127[12] 300[6])
    defparam i11208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11209_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n7330), 
            .I3(GND_net), .O(n15040));   // verilog/coms.v(127[12] 300[6])
    defparam i11209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11210_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n7330), 
            .I3(GND_net), .O(n15041));   // verilog/coms.v(127[12] 300[6])
    defparam i11210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11211_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n7330), 
            .I3(GND_net), .O(n15042));   // verilog/coms.v(127[12] 300[6])
    defparam i11211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11212_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n7330), 
            .I3(GND_net), .O(n15043));   // verilog/coms.v(127[12] 300[6])
    defparam i11212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11213_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n7330), 
            .I3(GND_net), .O(n15044));   // verilog/coms.v(127[12] 300[6])
    defparam i11213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11214_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n7330), 
            .I3(GND_net), .O(n15045));   // verilog/coms.v(127[12] 300[6])
    defparam i11214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24970_3_lut (.I0(n30134), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n30062));   // verilog/pwm.v(21[8:24])
    defparam i24970_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11215_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n7330), 
            .I3(GND_net), .O(n15046));   // verilog/coms.v(127[12] 300[6])
    defparam i11215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11216_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n7330), 
            .I3(GND_net), .O(n15047));   // verilog/coms.v(127[12] 300[6])
    defparam i11216_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_26[0]));   // verilog/TinyFPGA_B.v(200[10] 202[6])
    SB_LUT4 i11217_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n7330), 
            .I3(GND_net), .O(n15048));   // verilog/coms.v(127[12] 300[6])
    defparam i11217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11218_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n7330), 
            .I3(GND_net), .O(n15049));   // verilog/coms.v(127[12] 300[6])
    defparam i11218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11219_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n7330), 
            .I3(GND_net), .O(n15050));   // verilog/coms.v(127[12] 300[6])
    defparam i11219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11220_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n7330), 
            .I3(GND_net), .O(n15051));   // verilog/coms.v(127[12] 300[6])
    defparam i11220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24512_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n20610), 
            .I2(start), .I3(state[0]), .O(n29288));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24512_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_LUT4 i11221_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n7330), 
            .I3(GND_net), .O(n15052));   // verilog/coms.v(127[12] 300[6])
    defparam i11221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11222_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n7330), 
            .I3(GND_net), .O(n15053));   // verilog/coms.v(127[12] 300[6])
    defparam i11222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11223_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n7330), 
            .I3(GND_net), .O(n15054));   // verilog/coms.v(127[12] 300[6])
    defparam i11223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11224_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n7330), 
            .I3(GND_net), .O(n15055));   // verilog/coms.v(127[12] 300[6])
    defparam i11224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11225_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n7330), 
            .I3(GND_net), .O(n15056));   // verilog/coms.v(127[12] 300[6])
    defparam i11225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11226_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n10927), .I3(GND_net), .O(n15057));   // verilog/coms.v(127[12] 300[6])
    defparam i11226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11227_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n10927), .I3(GND_net), .O(n15058));   // verilog/coms.v(127[12] 300[6])
    defparam i11227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11228_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n10927), .I3(GND_net), .O(n15059));   // verilog/coms.v(127[12] 300[6])
    defparam i11228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11229_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n10927), .I3(GND_net), .O(n15060));   // verilog/coms.v(127[12] 300[6])
    defparam i11229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11230_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n10927), .I3(GND_net), .O(n15061));   // verilog/coms.v(127[12] 300[6])
    defparam i11230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11231_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n10927), .I3(GND_net), .O(n15062));   // verilog/coms.v(127[12] 300[6])
    defparam i11231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11232_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n10927), .I3(GND_net), .O(n15063));   // verilog/coms.v(127[12] 300[6])
    defparam i11232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11233_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n10927), .I3(GND_net), .O(n15064));   // verilog/coms.v(127[12] 300[6])
    defparam i11233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11234_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n10927), .I3(GND_net), .O(n15065));   // verilog/coms.v(127[12] 300[6])
    defparam i11234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11110_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4167), .I3(GND_net), .O(n14941));   // verilog/coms.v(127[12] 300[6])
    defparam i11110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11235_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n10927), .I3(GND_net), .O(n15066));   // verilog/coms.v(127[12] 300[6])
    defparam i11235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11236_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n10927), .I3(GND_net), .O(n15067));   // verilog/coms.v(127[12] 300[6])
    defparam i11236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11237_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n10927), .I3(GND_net), .O(n15068));   // verilog/coms.v(127[12] 300[6])
    defparam i11237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11238_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n10927), .I3(GND_net), .O(n15069));   // verilog/coms.v(127[12] 300[6])
    defparam i11238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11239_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n10927), .I3(GND_net), .O(n15070));   // verilog/coms.v(127[12] 300[6])
    defparam i11239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11240_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n10927), .I3(GND_net), .O(n15071));   // verilog/coms.v(127[12] 300[6])
    defparam i11240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11241_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n10927), .I3(GND_net), .O(n15072));   // verilog/coms.v(127[12] 300[6])
    defparam i11241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24971_3_lut (.I0(n30062), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n30063));   // verilog/pwm.v(21[8:24])
    defparam i24971_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11242_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n10927), .I3(GND_net), .O(n15073));   // verilog/coms.v(127[12] 300[6])
    defparam i11242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11243_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n10927), .I3(GND_net), .O(n15074));   // verilog/coms.v(127[12] 300[6])
    defparam i11243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11244_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n10927), .I3(GND_net), .O(n15075));   // verilog/coms.v(127[12] 300[6])
    defparam i11244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11245_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n10927), .I3(GND_net), .O(n15076));   // verilog/coms.v(127[12] 300[6])
    defparam i11245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11246_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n10927), .I3(GND_net), .O(n15077));   // verilog/coms.v(127[12] 300[6])
    defparam i11246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11247_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n10927), .I3(GND_net), .O(n15078));   // verilog/coms.v(127[12] 300[6])
    defparam i11247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11248_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n10927), .I3(GND_net), .O(n15079));   // verilog/coms.v(127[12] 300[6])
    defparam i11248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11249_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n10927), .I3(GND_net), .O(n15080));   // verilog/coms.v(127[12] 300[6])
    defparam i11249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11250_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n10927), .I3(GND_net), .O(n15081));   // verilog/coms.v(127[12] 300[6])
    defparam i11250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11251_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n10927), .I3(GND_net), .O(n15082));   // verilog/coms.v(127[12] 300[6])
    defparam i11251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11252_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n10927), .I3(GND_net), .O(n15083));   // verilog/coms.v(127[12] 300[6])
    defparam i11252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11253_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n10927), .I3(GND_net), .O(n15084));   // verilog/coms.v(127[12] 300[6])
    defparam i11253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11254_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n10927), .I3(GND_net), .O(n15085));   // verilog/coms.v(127[12] 300[6])
    defparam i11254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11255_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n10927), .I3(GND_net), .O(n15086));   // verilog/coms.v(127[12] 300[6])
    defparam i11255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11256_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n10927), .I3(GND_net), .O(n15087));   // verilog/coms.v(127[12] 300[6])
    defparam i11256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11257_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n10927), .I3(GND_net), .O(n15088));   // verilog/coms.v(127[12] 300[6])
    defparam i11257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11258_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n10927), .I3(GND_net), .O(n15089));   // verilog/coms.v(127[12] 300[6])
    defparam i11258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11259_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n10927), .I3(GND_net), .O(n15090));   // verilog/coms.v(127[12] 300[6])
    defparam i11259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11260_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n10927), .I3(GND_net), .O(n15091));   // verilog/coms.v(127[12] 300[6])
    defparam i11260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11261_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n10927), .I3(GND_net), .O(n15092));   // verilog/coms.v(127[12] 300[6])
    defparam i11261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11262_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n10927), .I3(GND_net), .O(n15093));   // verilog/coms.v(127[12] 300[6])
    defparam i11262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11263_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n10927), .I3(GND_net), .O(n15094));   // verilog/coms.v(127[12] 300[6])
    defparam i11263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11264_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n10927), .I3(GND_net), .O(n15095));   // verilog/coms.v(127[12] 300[6])
    defparam i11264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11114_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n18503), 
            .I3(n13657), .O(n14945));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11114_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i11115_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n18503), 
            .I3(n13652), .O(n14946));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11115_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_37_i1_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[0]), 
            .I3(encoder0_position[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11116_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n14947));   // verilog/coms.v(127[12] 300[6])
    defparam i11116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11117_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n7330), 
            .I3(GND_net), .O(n14948));   // verilog/coms.v(127[12] 300[6])
    defparam i11117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11118_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n7330), 
            .I3(GND_net), .O(n14949));   // verilog/coms.v(127[12] 300[6])
    defparam i11118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11265_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n10927), .I3(GND_net), .O(n15096));   // verilog/coms.v(127[12] 300[6])
    defparam i11265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11266_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n10927), .I3(GND_net), .O(n15097));   // verilog/coms.v(127[12] 300[6])
    defparam i11266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i2_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[1]), 
            .I3(encoder0_position[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11267_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n10927), .I3(GND_net), .O(n15098));   // verilog/coms.v(127[12] 300[6])
    defparam i11267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11268_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n10927), .I3(GND_net), .O(n15099));   // verilog/coms.v(127[12] 300[6])
    defparam i11268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11269_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n10927), .I3(GND_net), .O(n15100));   // verilog/coms.v(127[12] 300[6])
    defparam i11269_3_lut.LUT_INIT = 16'hcaca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4476, 
            quadB_debounced_adj_4477}), .n27693(n27693), .reg_B({reg_B_adj_4587}), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .VCC_net(VCC_net), .n15442(n15442), .n14956(n14956)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    SB_LUT4 i11270_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n10927), .I3(GND_net), .O(n15101));   // verilog/coms.v(127[12] 300[6])
    defparam i11270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11271_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n10927), .I3(GND_net), .O(n15102));   // verilog/coms.v(127[12] 300[6])
    defparam i11271_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i11119_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n4169), .I3(GND_net), .O(n14950));   // verilog/coms.v(127[12] 300[6])
    defparam i11119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11121_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4167), .I3(GND_net), .O(n14952));   // verilog/coms.v(127[12] 300[6])
    defparam i11121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11122_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n4167), .I3(GND_net), .O(n14953));   // verilog/coms.v(127[12] 300[6])
    defparam i11122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11123_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n28252), 
            .I3(GND_net), .O(n14954));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24929_3_lut (.I0(n30063), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n30021));   // verilog/pwm.v(21[8:24])
    defparam i24929_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i11124_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_4574[1]), .I2(n7410), 
            .I3(n4_adj_4471), .O(n14955));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i11124_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i11125_3_lut (.I0(quadB_debounced_adj_4477), .I1(reg_B_adj_4587[0]), 
            .I2(n27693), .I3(GND_net), .O(n14956));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i11125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_37_i3_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[2]), 
            .I3(encoder0_position[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11272_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n10927), .I3(GND_net), .O(n15103));   // verilog/coms.v(127[12] 300[6])
    defparam i11272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11273_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n10927), .I3(GND_net), .O(n15104));   // verilog/coms.v(127[12] 300[6])
    defparam i11273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11274_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n10927), .I3(GND_net), .O(n15105));   // verilog/coms.v(127[12] 300[6])
    defparam i11274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11275_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n10927), .I3(GND_net), .O(n15106));   // verilog/coms.v(127[12] 300[6])
    defparam i11275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11276_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n10927), .I3(GND_net), .O(n15107));   // verilog/coms.v(127[12] 300[6])
    defparam i11276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11277_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n10927), .I3(GND_net), .O(n15108));   // verilog/coms.v(127[12] 300[6])
    defparam i11277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i4_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[3]), 
            .I3(encoder0_position[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11278_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n10927), .I3(GND_net), .O(n15109));   // verilog/coms.v(127[12] 300[6])
    defparam i11278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11279_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n10927), .I3(GND_net), .O(n15110));   // verilog/coms.v(127[12] 300[6])
    defparam i11279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11280_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n10927), .I3(GND_net), .O(n15111));   // verilog/coms.v(127[12] 300[6])
    defparam i11280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11281_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n10927), .I3(GND_net), .O(n15112));   // verilog/coms.v(127[12] 300[6])
    defparam i11281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11282_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n10927), .I3(GND_net), .O(n15113));   // verilog/coms.v(127[12] 300[6])
    defparam i11282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i5_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[4]), 
            .I3(encoder0_position[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11283_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n10927), .I3(GND_net), .O(n15114));   // verilog/coms.v(127[12] 300[6])
    defparam i11283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11284_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n10927), .I3(GND_net), .O(n15115));   // verilog/coms.v(127[12] 300[6])
    defparam i11284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11285_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n10927), .I3(GND_net), .O(n15116));   // verilog/coms.v(127[12] 300[6])
    defparam i11285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11286_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n10927), .I3(GND_net), .O(n15117));   // verilog/coms.v(127[12] 300[6])
    defparam i11286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11287_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n10927), .I3(GND_net), .O(n15118));   // verilog/coms.v(127[12] 300[6])
    defparam i11287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11288_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n10927), .I3(GND_net), .O(n15119));   // verilog/coms.v(127[12] 300[6])
    defparam i11288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11289_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n10927), .I3(GND_net), .O(n15120));   // verilog/coms.v(127[12] 300[6])
    defparam i11289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i6_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[5]), 
            .I3(encoder0_position[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_37_i7_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[6]), 
            .I3(encoder0_position[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11290_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n10927), .I3(GND_net), .O(n15121));   // verilog/coms.v(127[12] 300[6])
    defparam i11290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11291_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n10927), .I3(GND_net), .O(n15122));   // verilog/coms.v(127[12] 300[6])
    defparam i11291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11292_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n10927), .I3(GND_net), .O(n15123));   // verilog/coms.v(127[12] 300[6])
    defparam i11292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11293_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n10927), .I3(GND_net), .O(n15124));   // verilog/coms.v(127[12] 300[6])
    defparam i11293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11294_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n10927), .I3(GND_net), .O(n15125));   // verilog/coms.v(127[12] 300[6])
    defparam i11294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11295_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n10927), .I3(GND_net), .O(n15126));   // verilog/coms.v(127[12] 300[6])
    defparam i11295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11296_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n10927), .I3(GND_net), .O(n15127));   // verilog/coms.v(127[12] 300[6])
    defparam i11296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11297_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n10927), .I3(GND_net), .O(n15128));   // verilog/coms.v(127[12] 300[6])
    defparam i11297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11298_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n10927), .I3(GND_net), .O(n15129));   // verilog/coms.v(127[12] 300[6])
    defparam i11298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11299_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n10927), .I3(GND_net), .O(n15130));   // verilog/coms.v(127[12] 300[6])
    defparam i11299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11300_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n10927), .I3(GND_net), .O(n15131));   // verilog/coms.v(127[12] 300[6])
    defparam i11300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11301_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n10927), .I3(GND_net), .O(n15132));   // verilog/coms.v(127[12] 300[6])
    defparam i11301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11302_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n10927), .I3(GND_net), .O(n15133));   // verilog/coms.v(127[12] 300[6])
    defparam i11302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11303_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n10927), .I3(GND_net), .O(n15134));   // verilog/coms.v(127[12] 300[6])
    defparam i11303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11304_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n10927), .I3(GND_net), .O(n15135));   // verilog/coms.v(127[12] 300[6])
    defparam i11304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11305_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n10927), .I3(GND_net), .O(n15136));   // verilog/coms.v(127[12] 300[6])
    defparam i11305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i8_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[7]), 
            .I3(encoder0_position[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11306_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n10927), 
            .I3(GND_net), .O(n15137));   // verilog/coms.v(127[12] 300[6])
    defparam i11306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11307_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n10927), 
            .I3(GND_net), .O(n15138));   // verilog/coms.v(127[12] 300[6])
    defparam i11307_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 i11308_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n10927), 
            .I3(GND_net), .O(n15139));   // verilog/coms.v(127[12] 300[6])
    defparam i11308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11309_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n10927), 
            .I3(GND_net), .O(n15140));   // verilog/coms.v(127[12] 300[6])
    defparam i11309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11310_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n10927), 
            .I3(GND_net), .O(n15141));   // verilog/coms.v(127[12] 300[6])
    defparam i11310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11311_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n10927), 
            .I3(GND_net), .O(n15142));   // verilog/coms.v(127[12] 300[6])
    defparam i11311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11312_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n10927), 
            .I3(GND_net), .O(n15143));   // verilog/coms.v(127[12] 300[6])
    defparam i11312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11313_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n10927), 
            .I3(GND_net), .O(n15144));   // verilog/coms.v(127[12] 300[6])
    defparam i11313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11314_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n10927), 
            .I3(GND_net), .O(n15145));   // verilog/coms.v(127[12] 300[6])
    defparam i11314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11315_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n10927), 
            .I3(GND_net), .O(n15146));   // verilog/coms.v(127[12] 300[6])
    defparam i11315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11316_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n10927), 
            .I3(GND_net), .O(n15147));   // verilog/coms.v(127[12] 300[6])
    defparam i11316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11317_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n10927), 
            .I3(GND_net), .O(n15148));   // verilog/coms.v(127[12] 300[6])
    defparam i11317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11318_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n10927), 
            .I3(GND_net), .O(n15149));   // verilog/coms.v(127[12] 300[6])
    defparam i11318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11319_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n10927), 
            .I3(GND_net), .O(n15150));   // verilog/coms.v(127[12] 300[6])
    defparam i11319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11320_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n10927), 
            .I3(GND_net), .O(n15151));   // verilog/coms.v(127[12] 300[6])
    defparam i11320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11321_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n10927), 
            .I3(GND_net), .O(n15152));   // verilog/coms.v(127[12] 300[6])
    defparam i11321_3_lut.LUT_INIT = 16'hcaca;
    motorControl control (.\Ki[1] (Ki[1]), .GND_net(GND_net), .\Ki[8] (Ki[8]), 
            .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .PWMLimit({PWMLimit}), .\Ki[3] (Ki[3]), 
            .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Kp[5] (Kp[5]), .\Kp[1] (Kp[1]), 
            .IntegralLimit({IntegralLimit}), .duty({duty}), .\Kp[9] (Kp[9]), 
            .\Kp[6] (Kp[6]), .\Kp[4] (Kp[4]), .\Kp[3] (Kp[3]), .\Kp[2] (Kp[2]), 
            .\Kp[0] (Kp[0]), .\Kp[10] (Kp[10]), .\Kp[8] (Kp[8]), .\Kp[7] (Kp[7]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Kp[15] (Kp[15]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .clk32MHz(clk32MHz), 
            .n30253(n30253), .VCC_net(VCC_net), .setpoint({setpoint}), 
            .motor_state({motor_state}), .n25(n25)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_LUT4 i11322_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n10927), 
            .I3(GND_net), .O(n15153));   // verilog/coms.v(127[12] 300[6])
    defparam i11322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11323_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n10927), 
            .I3(GND_net), .O(n15154));   // verilog/coms.v(127[12] 300[6])
    defparam i11323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i9_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[8]), 
            .I3(encoder0_position[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11324_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n10927), 
            .I3(GND_net), .O(n15155));   // verilog/coms.v(127[12] 300[6])
    defparam i11324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11325_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n10927), 
            .I3(GND_net), .O(n15156));   // verilog/coms.v(127[12] 300[6])
    defparam i11325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i10_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[9]), 
            .I3(encoder0_position[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_38_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_37_i11_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[10]), 
            .I3(encoder0_position[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11326_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n10927), 
            .I3(GND_net), .O(n15157));   // verilog/coms.v(127[12] 300[6])
    defparam i11326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i12_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[11]), 
            .I3(encoder0_position[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11327_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n10927), 
            .I3(GND_net), .O(n15158));   // verilog/coms.v(127[12] 300[6])
    defparam i11327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i13_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[12]), 
            .I3(encoder0_position[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11328_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n10927), 
            .I3(GND_net), .O(n15159));   // verilog/coms.v(127[12] 300[6])
    defparam i11328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11329_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n10927), 
            .I3(GND_net), .O(n15160));   // verilog/coms.v(127[12] 300[6])
    defparam i11329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11330_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n10927), .I3(GND_net), .O(n15161));   // verilog/coms.v(127[12] 300[6])
    defparam i11330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_38_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4467), .I3(n15), .O(motor_state_23__N_50[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_38_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i11331_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n10927), .I3(GND_net), .O(n15162));   // verilog/coms.v(127[12] 300[6])
    defparam i11331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11332_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n10927), .I3(GND_net), .O(n15163));   // verilog/coms.v(127[12] 300[6])
    defparam i11332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11333_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n10927), .I3(GND_net), .O(n15164));   // verilog/coms.v(127[12] 300[6])
    defparam i11333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i14_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[13]), 
            .I3(encoder0_position[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11334_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n10927), .I3(GND_net), .O(n15165));   // verilog/coms.v(127[12] 300[6])
    defparam i11334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11335_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n10927), .I3(GND_net), .O(n15166));   // verilog/coms.v(127[12] 300[6])
    defparam i11335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_37_i15_3_lut_4_lut (.I0(n13493), .I1(control_mode[1]), .I2(motor_state_23__N_50[14]), 
            .I3(encoder0_position[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_37_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i11336_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n10927), .I3(GND_net), .O(n15167));   // verilog/coms.v(127[12] 300[6])
    defparam i11336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11337_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n10927), .I3(GND_net), .O(n15168));   // verilog/coms.v(127[12] 300[6])
    defparam i11337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11338_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n10927), .I3(GND_net), .O(n15169));   // verilog/coms.v(127[12] 300[6])
    defparam i11338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11339_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n10927), .I3(GND_net), .O(n15170));   // verilog/coms.v(127[12] 300[6])
    defparam i11339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_4472), .I3(control_mode[2]), .O(n13493));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11340_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n10927), .I3(GND_net), .O(n15171));   // verilog/coms.v(127[12] 300[6])
    defparam i11340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11341_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n10927), .I3(GND_net), .O(n15172));   // verilog/coms.v(127[12] 300[6])
    defparam i11341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11342_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n10927), .I3(GND_net), .O(n15173));   // verilog/coms.v(127[12] 300[6])
    defparam i11342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11343_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n10927), .I3(GND_net), .O(n15174));   // verilog/coms.v(127[12] 300[6])
    defparam i11343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11344_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n10927), .I3(GND_net), .O(n15175));   // verilog/coms.v(127[12] 300[6])
    defparam i11344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11345_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n10927), .I3(GND_net), .O(n15176));   // verilog/coms.v(127[12] 300[6])
    defparam i11345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11346_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n10927), .I3(GND_net), .O(n15177));   // verilog/coms.v(127[12] 300[6])
    defparam i11346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11347_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n10927), .I3(GND_net), .O(n15178));   // verilog/coms.v(127[12] 300[6])
    defparam i11347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11348_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n10927), .I3(GND_net), .O(n15179));   // verilog/coms.v(127[12] 300[6])
    defparam i11348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11349_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n10927), .I3(GND_net), .O(n15180));   // verilog/coms.v(127[12] 300[6])
    defparam i11349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11350_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n10927), .I3(GND_net), .O(n15181));   // verilog/coms.v(127[12] 300[6])
    defparam i11350_3_lut.LUT_INIT = 16'hcaca;
    coms neopxl_color_23__I_0 (.\data_out_frame[19] ({\data_out_frame[19] }), 
         .n15009(n15009), .\data_in[1] ({\data_in[1] }), .clk32MHz(clk32MHz), 
         .GND_net(GND_net), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .setpoint({setpoint}), .n15008(n15008), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n15007(n15007), .n4167(n4167), .n10927(n10927), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .n4169(n4169), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .rx_data({rx_data}), 
         .n15006(n15006), .\data_in_frame[1] ({\data_in_frame[1] }), .n15005(n15005), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n15004(n15004), .n15003(n15003), 
         .n15002(n15002), .\data_in[0] ({\data_in[0] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .n15001(n15001), .n15000(n15000), .n14999(n14999), .rx_data_ready(rx_data_ready), 
         .n14998(n14998), .n14997(n14997), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n14996(n14996), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .n123(n123), .n63(n63), 
         .n13620(n13620), .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .n3303(n3303), .\FRAME_MATCHER.state_31__N_2508[1] (\FRAME_MATCHER.state_31__N_2508 [1]), 
         .n52(n52), .n7480(n7480), .\FRAME_MATCHER.state_31__N_2380[2] (\FRAME_MATCHER.state_31__N_2380 [2]), 
         .\FRAME_MATCHER.state_31__N_2540[2] (\FRAME_MATCHER.state_31__N_2540 [2]), 
         .\data_in[3] ({\data_in[3] }), .\data_in[2] ({\data_in[2] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .n63_adj_3(n63_adj_4473), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .n13615(n13615), .n26676(n26676), 
         .n13618(n13618), .n6(n6_adj_4527), .n14994(n14994), .IntegralLimit({IntegralLimit}), 
         .n14993(n14993), .tx_active(tx_active), .n14992(n14992), .DE_c(DE_c), 
         .LED_c(LED_c), .n14991(n14991), .n14990(n14990), .n14989(n14989), 
         .n14988(n14988), .n14987(n14987), .n14986(n14986), .n14985(n14985), 
         .n14984(n14984), .n14983(n14983), .n14982(n14982), .n14981(n14981), 
         .n14980(n14980), .n14979(n14979), .n14978(n14978), .n14977(n14977), 
         .n14976(n14976), .n14975(n14975), .n14974(n14974), .n14973(n14973), 
         .n14972(n14972), .n7330(n7330), .n30906(n30906), .n30907(n30907), 
         .n15436(n15436), .PWMLimit({PWMLimit}), .n15435(n15435), .n15434(n15434), 
         .n15433(n15433), .n15432(n15432), .n15431(n15431), .n15430(n15430), 
         .n15429(n15429), .n15428(n15428), .n15427(n15427), .n15426(n15426), 
         .n15425(n15425), .n15424(n15424), .n15423(n15423), .n15422(n15422), 
         .n15421(n15421), .n15420(n15420), .n15419(n15419), .n15418(n15418), 
         .n15417(n15417), .n15416(n15416), .n15415(n15415), .n15414(n15414), 
         .n15413(n15413), .control_mode({control_mode}), .n15412(n15412), 
         .n15411(n15411), .n15410(n15410), .n15409(n15409), .n15408(n15408), 
         .n15407(n15407), .n15231(n15231), .neopxl_color({neopxl_color}), 
         .n15230(n15230), .n15229(n15229), .n15228(n15228), .n15227(n15227), 
         .n15226(n15226), .n15225(n15225), .n15224(n15224), .n15223(n15223), 
         .n15222(n15222), .n15221(n15221), .n15220(n15220), .n15219(n15219), 
         .n15218(n15218), .n15217(n15217), .n15216(n15216), .n15215(n15215), 
         .n15214(n15214), .n15213(n15213), .n15212(n15212), .n15211(n15211), 
         .n15210(n15210), .n15209(n15209), .n15208(n15208), .n15207(n15207), 
         .n15206(n15206), .n15205(n15205), .n15204(n15204), .n15203(n15203), 
         .n15202(n15202), .n15201(n15201), .n15200(n15200), .n15199(n15199), 
         .n15198(n15198), .n15197(n15197), .n15196(n15196), .n15195(n15195), 
         .n15194(n15194), .n15193(n15193), .n15192(n15192), .n15191(n15191), 
         .n15190(n15190), .n15189(n15189), .n15188(n15188), .n15187(n15187), 
         .n15186(n15186), .n15185(n15185), .n15184(n15184), .n15183(n15183), 
         .n15182(n15182), .n15181(n15181), .n15180(n15180), .n15179(n15179), 
         .n15178(n15178), .n15177(n15177), .n15176(n15176), .n15175(n15175), 
         .n15174(n15174), .n15173(n15173), .n15172(n15172), .n15171(n15171), 
         .n15170(n15170), .n15169(n15169), .n15168(n15168), .n15167(n15167), 
         .n15166(n15166), .n15165(n15165), .n15164(n15164), .n15163(n15163), 
         .n15162(n15162), .n15161(n15161), .n15160(n15160), .n15159(n15159), 
         .n15158(n15158), .n15157(n15157), .n15156(n15156), .n15155(n15155), 
         .n15154(n15154), .n15153(n15153), .n15152(n15152), .n15151(n15151), 
         .n15150(n15150), .n15149(n15149), .n15148(n15148), .n15147(n15147), 
         .n15146(n15146), .n15145(n15145), .n15144(n15144), .n15143(n15143), 
         .n15142(n15142), .n15141(n15141), .n15140(n15140), .n15139(n15139), 
         .n15138(n15138), .n15137(n15137), .n15136(n15136), .n15135(n15135), 
         .n15134(n15134), .n15133(n15133), .n15132(n15132), .n15131(n15131), 
         .n15130(n15130), .n15129(n15129), .n15128(n15128), .n15127(n15127), 
         .n15126(n15126), .n15125(n15125), .n15124(n15124), .n15123(n15123), 
         .n15122(n15122), .n15121(n15121), .n15120(n15120), .n15119(n15119), 
         .n15118(n15118), .n15117(n15117), .n15116(n15116), .n15115(n15115), 
         .n15114(n15114), .n15113(n15113), .n15112(n15112), .n15111(n15111), 
         .n15110(n15110), .n15109(n15109), .n15108(n15108), .n15107(n15107), 
         .n15106(n15106), .n15105(n15105), .n15104(n15104), .n15103(n15103), 
         .n14953(n14953), .n14952(n14952), .n14950(n14950), .n15102(n15102), 
         .n15101(n15101), .n15100(n15100), .n15099(n15099), .n15098(n15098), 
         .n15097(n15097), .n15096(n15096), .n14949(n14949), .\Ki[0] (Ki[0]), 
         .n14948(n14948), .\Kp[0] (Kp[0]), .n14947(n14947), .n15095(n15095), 
         .n15094(n15094), .n15093(n15093), .n15092(n15092), .n15091(n15091), 
         .n15090(n15090), .n15089(n15089), .n15088(n15088), .n15087(n15087), 
         .n15086(n15086), .n15085(n15085), .n15084(n15084), .n15083(n15083), 
         .n15082(n15082), .n15081(n15081), .n15080(n15080), .n15079(n15079), 
         .n15078(n15078), .n15077(n15077), .n15076(n15076), .n15075(n15075), 
         .n15074(n15074), .n15073(n15073), .n15072(n15072), .n15071(n15071), 
         .n15070(n15070), .n15069(n15069), .n15068(n15068), .n15067(n15067), 
         .n15066(n15066), .n14941(n14941), .n15065(n15065), .n15064(n15064), 
         .n15063(n15063), .n15062(n15062), .n15061(n15061), .n15060(n15060), 
         .n15059(n15059), .n15058(n15058), .n15057(n15057), .n15056(n15056), 
         .\Ki[15] (Ki[15]), .n15055(n15055), .\Ki[14] (Ki[14]), .n15054(n15054), 
         .\Ki[13] (Ki[13]), .n15053(n15053), .\Ki[12] (Ki[12]), .n15052(n15052), 
         .\Ki[11] (Ki[11]), .n15051(n15051), .\Ki[10] (Ki[10]), .n15050(n15050), 
         .\Ki[9] (Ki[9]), .n15049(n15049), .\Ki[8] (Ki[8]), .n15048(n15048), 
         .\Ki[7] (Ki[7]), .n15047(n15047), .\Ki[6] (Ki[6]), .n15046(n15046), 
         .\Ki[5] (Ki[5]), .n15045(n15045), .\Ki[4] (Ki[4]), .n15044(n15044), 
         .\Ki[3] (Ki[3]), .n15043(n15043), .\Ki[2] (Ki[2]), .n15042(n15042), 
         .\Ki[1] (Ki[1]), .n15041(n15041), .\Kp[15] (Kp[15]), .n15040(n15040), 
         .\Kp[14] (Kp[14]), .n15039(n15039), .\Kp[13] (Kp[13]), .n15038(n15038), 
         .\Kp[12] (Kp[12]), .n15037(n15037), .\Kp[11] (Kp[11]), .n15036(n15036), 
         .\Kp[10] (Kp[10]), .n15035(n15035), .\Kp[9] (Kp[9]), .n15034(n15034), 
         .\Kp[8] (Kp[8]), .n15033(n15033), .\Kp[7] (Kp[7]), .n15032(n15032), 
         .\Kp[6] (Kp[6]), .n15031(n15031), .\Kp[5] (Kp[5]), .n15030(n15030), 
         .\Kp[4] (Kp[4]), .n15029(n15029), .\Kp[3] (Kp[3]), .n15028(n15028), 
         .\Kp[2] (Kp[2]), .n15027(n15027), .\Kp[1] (Kp[1]), .n15026(n15026), 
         .n15025(n15025), .n15024(n15024), .n15023(n15023), .n15022(n15022), 
         .n15021(n15021), .n15020(n15020), .n15019(n15019), .n15018(n15018), 
         .n15017(n15017), .n15016(n15016), .n15015(n15015), .n15014(n15014), 
         .n15013(n15013), .n15012(n15012), .n15011(n15011), .n15010(n15010), 
         .n26810(n26810), .n26830(n26830), .\r_Bit_Index[0] (r_Bit_Index_adj_4576[0]), 
         .r_SM_Main({r_SM_Main_adj_4574}), .tx_o(tx_o), .\r_SM_Main_2__N_3333[1] (r_SM_Main_2__N_3333[1]), 
         .VCC_net(VCC_net), .n14961(n14961), .n4(n4_adj_4471), .n14955(n14955), 
         .n30923(n30923), .n7410(n7410), .tx_enable(tx_enable), .n14794(n14794), 
         .n14921(n14921), .r_SM_Main_adj_11({r_SM_Main}), .r_Rx_Data(r_Rx_Data), 
         .RX_N_2(RX_N_2), .n14995(n14995), .\r_SM_Main_2__N_3262[2] (r_SM_Main_2__N_3262[2]), 
         .\r_Bit_Index[0]_adj_7 (r_Bit_Index[0]), .n13657(n13657), .n4_adj_8(n4_adj_4487), 
         .n4_adj_9(n4), .n13652(n13652), .n4_adj_10(n4_adj_4466), .n25972(n25972), 
         .n14971(n14971), .n14970(n14970), .n14969(n14969), .n14968(n14968), 
         .n14957(n14957), .n14964(n14964), .n25630(n25630), .n18503(n18503), 
         .n14946(n14946), .n14945(n14945)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    pwm PWM (.n30021(n30021), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n13483(n13483), .pwm_counter({pwm_counter}), .GND_net(GND_net), 
        .n13481(n13481)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(90[6] 95[3])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, clk32MHz, 
            data_o, n28252, reg_B, ENCODER0_B_c_0, VCC_net, n15441, 
            n14954, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n28252;
    output [1:0]reg_B;
    input ENCODER0_B_c_0;
    input VCC_net;
    input n15441;
    input n14954;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n22056, n2470, n22057;
    wire [23:0]n2474;
    
    wire n22055, n22054, n22053, count_enable, B_delayed, A_delayed, 
        n22052, n22051, n22050, n22049, n22048, n22047, n22046, 
        n22045, n22044, n22043, n22042, n22041, n22040, n22039, 
        n22038, count_direction, n22037, n22060, n22059, n22058;
    
    SB_CARRY add_554_21 (.CI(n22056), .I0(encoder0_position[19]), .I1(n2470), 
            .CO(n22057));
    SB_LUT4 add_554_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2470), 
            .I3(n22055), .O(n2474[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_20 (.CI(n22055), .I0(encoder0_position[18]), .I1(n2470), 
            .CO(n22056));
    SB_LUT4 add_554_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2470), 
            .I3(n22054), .O(n2474[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_19 (.CI(n22054), .I0(encoder0_position[17]), .I1(n2470), 
            .CO(n22055));
    SB_LUT4 add_554_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2470), 
            .I3(n22053), .O(n2474[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_554_18 (.CI(n22053), .I0(encoder0_position[16]), .I1(n2470), 
            .CO(n22054));
    SB_LUT4 add_554_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2470), 
            .I3(n22052), .O(n2474[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_17 (.CI(n22052), .I0(encoder0_position[15]), .I1(n2470), 
            .CO(n22053));
    SB_LUT4 add_554_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2470), 
            .I3(n22051), .O(n2474[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_16 (.CI(n22051), .I0(encoder0_position[14]), .I1(n2470), 
            .CO(n22052));
    SB_LUT4 add_554_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2470), 
            .I3(n22050), .O(n2474[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_15 (.CI(n22050), .I0(encoder0_position[13]), .I1(n2470), 
            .CO(n22051));
    SB_LUT4 add_554_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2470), 
            .I3(n22049), .O(n2474[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_14 (.CI(n22049), .I0(encoder0_position[12]), .I1(n2470), 
            .CO(n22050));
    SB_LUT4 add_554_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2470), 
            .I3(n22048), .O(n2474[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_13 (.CI(n22048), .I0(encoder0_position[11]), .I1(n2470), 
            .CO(n22049));
    SB_LUT4 add_554_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2470), 
            .I3(n22047), .O(n2474[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_12 (.CI(n22047), .I0(encoder0_position[10]), .I1(n2470), 
            .CO(n22048));
    SB_LUT4 add_554_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2470), 
            .I3(n22046), .O(n2474[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_11 (.CI(n22046), .I0(encoder0_position[9]), .I1(n2470), 
            .CO(n22047));
    SB_LUT4 add_554_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2470), 
            .I3(n22045), .O(n2474[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_10 (.CI(n22045), .I0(encoder0_position[8]), .I1(n2470), 
            .CO(n22046));
    SB_LUT4 add_554_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2470), 
            .I3(n22044), .O(n2474[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_9 (.CI(n22044), .I0(encoder0_position[7]), .I1(n2470), 
            .CO(n22045));
    SB_LUT4 add_554_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2470), 
            .I3(n22043), .O(n2474[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_8 (.CI(n22043), .I0(encoder0_position[6]), .I1(n2470), 
            .CO(n22044));
    SB_LUT4 add_554_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2470), 
            .I3(n22042), .O(n2474[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_7 (.CI(n22042), .I0(encoder0_position[5]), .I1(n2470), 
            .CO(n22043));
    SB_LUT4 add_554_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2470), 
            .I3(n22041), .O(n2474[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_6 (.CI(n22041), .I0(encoder0_position[4]), .I1(n2470), 
            .CO(n22042));
    SB_LUT4 add_554_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2470), 
            .I3(n22040), .O(n2474[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_5 (.CI(n22040), .I0(encoder0_position[3]), .I1(n2470), 
            .CO(n22041));
    SB_LUT4 add_554_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2470), 
            .I3(n22039), .O(n2474[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_4 (.CI(n22039), .I0(encoder0_position[2]), .I1(n2470), 
            .CO(n22040));
    SB_LUT4 add_554_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2470), 
            .I3(n22038), .O(n2474[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_3 (.CI(n22038), .I0(encoder0_position[1]), .I1(n2470), 
            .CO(n22039));
    SB_LUT4 add_554_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n22037), .O(n2474[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_2 (.CI(n22037), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n22038));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_554_1 (.CI(GND_net), .I0(n2470), .I1(n2470), .CO(n22037));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2474[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 i846_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2470));   // quad.v(37[5] 40[8])
    defparam i846_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_554_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2470), 
            .I3(n22060), .O(n2474[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_554_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2470), 
            .I3(n22059), .O(n2474[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_24 (.CI(n22059), .I0(encoder0_position[22]), .I1(n2470), 
            .CO(n22060));
    SB_LUT4 add_554_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2470), 
            .I3(n22058), .O(n2474[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_23 (.CI(n22058), .I0(encoder0_position[21]), .I1(n2470), 
            .CO(n22059));
    SB_LUT4 add_554_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2470), 
            .I3(n22057), .O(n2474[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_554_22 (.CI(n22057), .I0(encoder0_position[20]), .I1(n2470), 
            .CO(n22058));
    SB_LUT4 add_554_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2470), 
            .I3(n22056), .O(n2474[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_554_21_lut.LUT_INIT = 16'hC33C;
    \grp_debouncer(2,100)_U0  debounce (.n28252(n28252), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .VCC_net(VCC_net), .n15441(n15441), .data_o({data_o}), .n14954(n14954), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n28252, reg_B, GND_net, clk32MHz, 
            ENCODER0_B_c_0, VCC_net, n15441, data_o, n14954, ENCODER0_A_c_1);
    output n28252;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input ENCODER0_B_c_0;
    input VCC_net;
    input n15441;
    output [1:0]data_o;
    input n14954;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3576;
    wire [6:0]n33;
    
    wire n22445, n22444, n22443, n22442, n22441, n22440;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n28252));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n28252), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1133__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1133_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22445), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1133_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22444), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_7 (.CI(n22444), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22445));
    SB_LUT4 cnt_reg_1133_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22443), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_6 (.CI(n22443), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22444));
    SB_LUT4 cnt_reg_1133_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22442), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_5 (.CI(n22442), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22443));
    SB_LUT4 cnt_reg_1133_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22441), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_4 (.CI(n22441), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22442));
    SB_LUT4 cnt_reg_1133_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22440), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_3 (.CI(n22440), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22441));
    SB_LUT4 cnt_reg_1133_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1133_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1133_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22440));
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n15441));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n14954));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1133__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1133__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1133__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1133__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1133__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1133__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.t0 , GND_net, \neo_pixel_transmitter.done , 
            clk32MHz, timer, VCC_net, start, \state[0] , \state[1] , 
            n4, n20610, n107, n26721, n27279, n1554, neopxl_color, 
            n14958, n15476, n15475, n15474, n15473, n15472, n15471, 
            n15470, n15469, n15468, n15467, n15466, n15465, n15464, 
            n15463, n15462, n15461, n15460, n15459, n15458, n15457, 
            n15456, n15455, n15454, n15453, n15452, n15451, n15450, 
            n15449, n15448, n15447, n15446, n24720, LED_c, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output [31:0]timer;
    input VCC_net;
    output start;
    output \state[0] ;
    output \state[1] ;
    output n4;
    output n20610;
    output n107;
    output n26721;
    output n27279;
    output n1554;
    input [23:0]neopxl_color;
    input n14958;
    input n15476;
    input n15475;
    input n15474;
    input n15473;
    input n15472;
    input n15471;
    input n15470;
    input n15469;
    input n15468;
    input n15467;
    input n15466;
    input n15465;
    input n15464;
    input n15463;
    input n15462;
    input n15461;
    input n15460;
    input n15459;
    input n15458;
    input n15457;
    input n15456;
    input n15455;
    input n15454;
    input n15453;
    input n15452;
    input n15451;
    input n15450;
    input n15449;
    input n15448;
    input n15447;
    input n15446;
    input n24720;
    input LED_c;
    output NEOPXL_c;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n56;
    
    wire n1897, n1798, n1829, n22267, \neo_pixel_transmitter.done_N_456 , 
        n25967;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n1409, n19021, n1405, n1403, n1406, n16, n1402, n1404, 
        n1400, n1407, n17, n22345, n22346, n1408, n1401, n1433, 
        n22268;
    wire [31:0]n133;
    
    wire n22344;
    wire [31:0]n255;
    
    wire n14736, n14862, n1334, n30257, n3004, n2989, n2990, n3007, 
        n40, n3006, n2984, n2988, n2986, n44, n3008, n3003, 
        n2994, n3002, n42, n2999, n3000, n2992, n2997, n43, 
        n2996, n2985, n2995, n2987, n41, n3001, n2993, n38, 
        n2998, n2991, n46, n50, n3005, n3009, n37, n3017, n22343, 
        n21915, n1898, n1799, n22266, n22006, n2199, n2225, n22007, 
        n2299, n2200, n22005, n21916, n21907, n2390, n2291, n2324, 
        n23155, n2391, n2292, n23154, n2392, n2293, n23153, n2393, 
        n2294, n23152, n2394, n2295, n23151, n2395, n2296, n23150, 
        n2396, n2297, n23149, n2397, n2298, n23148, n2398, n23147, 
        n2399, n2300, n23146, n2400, n2301, n23145, n2401, n2302, 
        n23144, n2402, n2303, n23143, n2403, n2304, n23142, n2404, 
        n2305, n23141, n2405, n2306, n23140, n2406, n2307, n23139, 
        n2407, n2308, n23138, n2408, n2309, n30252, n23137, n2409, 
        n3116, n30256, n1304, n1305, n10_adj_4312, n1303, n1309, 
        n12_adj_4313, n1306, n1308, n1302, n16_adj_4314, n1307, 
        n1301, n1998, n2004, n18, n2003, n1999, n1996, n2007, 
        n28, n1997, n2005, n2000, n2002, n26, n2001, n2008, 
        n1994, n1995, n27, n2006, n2009, n25, n2027, n22342, 
        n1235, n30255, n22341, n21908, n3102, n3090, n3103, n3085, 
        n42_adj_4315, n3089, n3094, n3101, n3098, n46_adj_4316, 
        n3099, n3091, n3106, n3100, n44_adj_4317, n3097, n3088, 
        n3104, n3092, n45, n3105, n3083, n3093, n3096, n43_adj_4318, 
        n3108, n3109, n40_adj_4319, n3107, n3087, n3086, n48, 
        n52, n3095, n3084, n39, n1928, n30254, n1899, n1800, 
        n22265, n22340, n21914, n3209, n18991, n35, n11_adj_4321, 
        n29, n51, n48_adj_4322, n37_adj_4323, n23, n53, n39_adj_4324, 
        n46_adj_4325, n27_adj_4326, n57, n63, n43_adj_4327, n47, 
        n25_adj_4328, n33, n47_adj_4329, n61, n45_adj_4330, n59, 
        n17_adj_4331, n15_adj_4332, n55, n44_adj_4333, n31, n41_adj_4334, 
        n49, n43_adj_4335, n54, n45_adj_4336, n13_adj_4337, n19_adj_4338, 
        n21, n49_adj_4339, n23352, n23676, n1506, n1503, n1500, 
        n1501, n18_adj_4340, n1504, n1502, n1499, n20, n1505, 
        n1509, n15_adj_4341, n1508, n1507, n1532, n2201, n22004, 
        n2908, n2909, n29_adj_4343, n2900, n2895, n2901, n2906, 
        n39_adj_4344, n2891, n2896, n2889, n38_adj_4345, n2897, 
        n2899, n2887, n2892, n43_adj_4346, n2905, n2903, n2888, 
        n2907, n42_adj_4347, n2898, n2886, n2893, n2904, n41_adj_4348, 
        n2890, n2902, n45_adj_4349, n2894, n2885, n47_adj_4350, 
        n2918, n30259, n30260, n2103, n2097, n18_adj_4351, n2109, 
        n18999, n2093, n2108, n2100, n30, n2098, n2094, n2099, 
        n28_adj_4352, n2105, n2096, n2095, n2102, n29_adj_4353, 
        n2101, n2107, n2104, n2106, n27_adj_4354, n2126, n1900, 
        n1801, n22264, n21906, n1901, n1802, n22263, n21913, n22339, 
        n2202, n22003, n1902, n1803, n22262, n30258, n2203, n22002, 
        n2204, n22001, n1903, n1804, n22261, n1904, n1805, n22260, 
        n22338, n2205, n22000, n1905, n1806, n22259, n22337, n21935, 
        n1906, n1807, n22258, n2206, n21999, n1907, n1808, n22257, 
        n21934, n22336, n2207, n21998, n1908, n1809, n30250, n22256, 
        n1205, n1206, n1204, n1207, n14_adj_4355, n1203, n1209, 
        n9_adj_4356, n1202, n1208, n2208, n21997, n22335, n2209, 
        n30251, n21996, n22334, n21933, n1909, n21912, n1895, 
        n22255, n21932, n22333, n1896, n22254, n21931, n22253, 
        n26_adj_4358, n19_adj_4359, n16_adj_4360, n24, n28_adj_4361, 
        n21905, n22252, n22332, n22251, n22331, n22250, n22249, 
        n22248, n22330, n22247, n22246, n21911, n21930, n22245, 
        n22244, n27_adj_4362, n22161;
    wire [31:0]one_wire_N_399;
    
    wire n22, n22160, n22243, n21929, n23_adj_4363, n22159, n28_adj_4364, 
        n22158, n21928, n22329, n26_adj_4365, n22157, n22242, n22_adj_4366, 
        n30_adj_4367, n34, n32, n33_adj_4368, n31_adj_4369, n22241, 
        n2193, n2194, n28_adj_4370, n32_adj_4371, n2192, n2196, 
        n30_adj_4372, n2195, n31_adj_4373, n2197, n2198, n29_adj_4374, 
        n22328, n22650, n22649, n22648, n46_adj_4375, n44_adj_4376, 
        n45_adj_4377, n43_adj_4378, n42_adj_4379, n41_adj_4380, n52_adj_4381, 
        n47_adj_4382, n11306, n28371, n20565, n33_adj_4383, n20572, 
        n6_adj_4384, n22647, n22646, n21927, n22645, n22644, n22643, 
        n22642, n29293, n13644, n1, n29274, n22641, n26806, n22640, 
        n22639, n21_adj_4386, n22156, n22327, n22326, n22638, n22637, 
        n22325, n22636, n22635, n22634, n22240, n22633, n22324, 
        n22239, n22323, n22155, n22322, n22321, n22238, n22632, 
        n22631, n22630, n1037, n30270, n2_adj_4387;
    wire [31:0]n971;
    
    wire n1007, n1006, n906, n1005, n14818, n905, n26696, n8_adj_4388, 
        n12170, n1009, n1008, n22629, n22154, n28385, n22320, 
        n22319, n22237, n22628, n22627, n6_adj_4389, n22236, n22626, 
        n22625, n22624, n26662, n11764, n807, n838, n4_adj_4390, 
        n29_adj_4391, n22153, n60, n22318, n22623, n22317, n22235, 
        n22152, n22316, n22622, n22621, n22620, n22619, n22618, 
        n22617, n22616, n22615, n22614, n22613, n22234, n22612, 
        n30_adj_4392, n22151, n22233, n22315, n608, n22314, n22232, 
        n708, n18738, n26710, n26798, n22611, n22610, n22609, 
        n22608, n22607, n22231, n22606, n22605, n23680, n24_adj_4393, 
        n22150, n22230, n22313, n22229, n2423, n30269, n27_adj_4394, 
        n33_adj_4395, n32_adj_4396, n31_adj_4397, n35_adj_4398, n37_adj_4399, 
        n2522, n30268, n22312, n22228, n25_adj_4400, n22149, n22311, 
        n22227, n22148, n22310, n22226, n22309, n22225, n22308, 
        n22147, n22604, n22603, n22307, n22602, n2491, n2504, 
        n24_adj_4401, n36, n2496, n2505, n2500, n2499, n34_adj_4402, 
        n37_adj_4403, n2497, n2509, n22_adj_4404, n2490, n2494, 
        n38_adj_4405, n2501, n2502, n2506, n2492, n36_adj_4406, 
        n2495, n2498, n2493, n37_adj_4407, n2507, n2508, n2503, 
        n2489, n35_adj_4408, n2621, n30266, n28317, n30568, n28389, 
        n22224, n22223, n22601, n22306, n22222, n21926, n22600, 
        n22599, n22598, n30478, n30481, n22597, n22596, n22221, 
        n22595, n22594, n22593, n22220, n30424, n28518, n30418, 
        n28521, n30406, n30409, n22146, n22592, n1598, n22305, 
        n30388, n29915, n30382, n30385, n22219, n22145, n22218, 
        n1599, n22304, n22144, n1600, n22303, n22591, n22590, 
        n22589, n22588, n22587, n22586, n22585, n22584, n22583, 
        n22582, n22217, n9_adj_4413, n7_adj_4414, n8_adj_4415, n22581, 
        n27201, n22580, n26727, n33_adj_4417, n22579, n22216, n22578, 
        n2591, n2608, n2601, n2605, n36_adj_4418, n2606, n2609, 
        n25_adj_4419, n2593, n2596, n2600, n2590, n34_adj_4420, 
        n2594, n2589, n40_adj_4421, n2602, n2588, n2604, n2607, 
        n38_adj_4422, n2598, n2603, n39_adj_4423, n2592, n2597, 
        n2595, n2599, n37_adj_4424, n1608, n1606, n1604, n1603, 
        n20_adj_4425, n1602, n1609, n13_adj_4426, n18_adj_4427, n1605, 
        n22_adj_4428, n1601, n1607, n1631, n22577, n22576, n2720, 
        n30265, n22215, n22575, n22574, n22302, color_bit;
    wire [3:0]state_3__N_248;
    
    wire n20573, n22143, n30263, n30262, n22573, n2786, n2819, 
        n22572, n2787, n22571, n21925, n2788, n22570, n2789, n22569, 
        n22301, n22214, n2790, n22568, n2791, n22567, n22300, 
        n22213, n30261, n22142, n2792, n22566, n22299, n22212, 
        n2793, n22565, n2794, n22564, n2795, n22563, n2796, n22562, 
        n21924, n2797, n22561, n22211, n2798, n22560, n2693, n2704, 
        n28_adj_4435, n2799, n22559, n22141, n22298, n2699, n2706, 
        n2694, n2691, n38_adj_4437, n2800, n22558, n22210, n2709, 
        n19005, n2701, n2696, n2697, n36_adj_4438, n2801, n22557, 
        n2700, n2705, n42_adj_4439, n2702, n2690, n2689, n2708, 
        n40_adj_4440, n22297, n2687, n2703, n2695, n41_adj_4441, 
        n2688, n2698, n2692, n2707, n39_adj_4442, n22296, n2802, 
        n22556, n21923, n2803, n22555, n30264, n20611, n21910, 
        n22140, n7_adj_4445, n20561, n2804, n22554, n22139, n2805, 
        n22553, n2806, n22552, n2807, n22551, n2808, n22550, n2809, 
        n22549, n22209, n22548, n22547, n22138, n22137, n22208, 
        n22546, n22545;
    wire [4:0]color_bit_N_442;
    
    wire n22544, n22_adj_4446, n22543, n22542, n22541, n22540, n22539, 
        n22538, n22295, n22537, n22136, n22536, n22535, n22534, 
        n22533, n22532, n22531, n22530, n24_adj_4447, n22529, n22528, 
        n22527, n22526, n22135, n1697, n22294, n22525, n21922, 
        n22524, n1698, n22293, n22523, n22522, n22521, n22520, 
        n22519, n22518, n22517, n22516, n22134, n22515, n40_adj_4448, 
        n1699, n22292, n22133, n22514, n22132, n38_adj_4449, n22513, 
        n22512, n21921, n39_adj_4450, n37_adj_4451, n22511, n22510, 
        n4_adj_4452, n22131, n34_adj_4453, n22509, n1700, n22291, 
        n22508, n22507, n42_adj_4454, n46_adj_4455, n33_adj_4456, 
        n22_adj_4457, n22506, n22505, n22504, n22503, n22502, n22501, 
        n22500, n22499, n1701, n22290, n22498, n22497, n22496, 
        n22495, n22494, n22493, n22492, n22491, n22490, n22489, 
        n22488, n22487, n22486, n22485, n22484, n1797, n23_adj_4458, 
        n1796, n21_adj_4459, n22483, n22482, n22481, n22480, n22479, 
        n22478, n22477, n22476, n22475, n22474, n22473, n22472, 
        n22471, n22470, n22469, n22468, n22467, n22466, n22465, 
        n22464, n22463, n22462, n22461, n22460, n22459, n22458, 
        n1103, n22457, n1104, n22456, n1105, n22455, n1106, n22454, 
        n1107, n22453, n1108, n22452, n1109, n1702, n22289, n21909, 
        n1703, n22288, n1704, n22287, n22013, n21920, n1705, n22286, 
        n1706, n22285, n1730, n30272, n28257, n1707, n22284, n21919, 
        n1708, n30267, n22283, \neo_pixel_transmitter.done_N_462 , n26842, 
        n22012, n21918, n1136, n22401, n22400, n22399, n22398, 
        n22397, n22396, n1709, n17_adj_4460, n21_adj_4461, n22011, 
        n20_adj_4462, n24_adj_4463, n30271, n22395, n22010, n11_adj_4464, 
        n21917, n22282, n22281, n22280, n22009, n22279, n22008, 
        n22278, n22277, n22276, n22275, n22274, n22273, n22272, 
        n19015, n22271, n12_adj_4465, n29601, n29332, n26838, n22270, 
        n22363, n22362, n22361, n22360, n22359, n22358, n22357, 
        n22356, n22355, n22354, n22269, n22353, n22352, n22351, 
        n22350, n22349, n22348, n22347;
    
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n22267), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n25967), .D(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i15193_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n19021));
    defparam i15193_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(n1405), .I1(n19021), .I2(n1403), .I3(n1406), 
            .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1126_add_4_15 (.CI(n22345), .I0(GND_net), .I1(timer[13]), 
            .CO(n22346));
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n1408), .I2(n16), .I3(n1401), .O(n1433));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1272_14 (.CI(n22267), .I0(n1798), .I1(n1829), .CO(n22268));
    SB_LUT4 timer_1126_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n22344), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n14736), 
            .D(n255[15]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i25167_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30257));
    defparam i25167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40), .I2(n2991), .I3(GND_net), 
            .O(n46));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37), .I1(n50), .I2(n46), .I3(n38), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1126_add_4_14 (.CI(n22344), .I0(GND_net), .I1(timer[12]), 
            .CO(n22345));
    SB_LUT4 timer_1126_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n22343), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n21915), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n22266), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n22006), .I0(n2199), .I1(n2225), .CO(n22007));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n22005), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n21915), .I0(bit_ctr[11]), .I1(GND_net), .CO(n21916));
    SB_CARRY mod_5_add_1540_12 (.CI(n22005), .I0(n2200), .I1(n2225), .CO(n22006));
    SB_CARRY mod_5_add_1272_13 (.CI(n22266), .I0(n1799), .I1(n1829), .CO(n22267));
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n21907), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n23155), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n23154), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n23154), .I0(n2292), .I1(n2324), .CO(n23155));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n23153), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n23153), .I0(n2293), .I1(n2324), .CO(n23154));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n23152), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n23152), .I0(n2294), .I1(n2324), .CO(n23153));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n23151), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n23151), .I0(n2295), .I1(n2324), .CO(n23152));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n23150), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n23150), .I0(n2296), .I1(n2324), .CO(n23151));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n23149), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n23149), .I0(n2297), .I1(n2324), .CO(n23150));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n23148), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n23148), .I0(n2298), .I1(n2324), .CO(n23149));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n23147), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n23147), .I0(n2299), .I1(n2324), .CO(n23148));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n23146), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n23146), .I0(n2300), .I1(n2324), .CO(n23147));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n23145), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n23145), .I0(n2301), .I1(n2324), .CO(n23146));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n23144), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n23144), .I0(n2302), .I1(n2324), .CO(n23145));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n23143), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n23143), .I0(n2303), .I1(n2324), .CO(n23144));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n23142), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n23142), .I0(n2304), .I1(n2324), .CO(n23143));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n23141), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n23141), .I0(n2305), .I1(n2324), .CO(n23142));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n23140), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n23140), .I0(n2306), .I1(n2324), .CO(n23141));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n23139), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n23139), .I0(n2307), .I1(n2324), .CO(n23140));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n23138), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n23138), .I0(n2308), .I1(n2324), .CO(n23139));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n30252), 
            .I3(n23137), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n23137), .I0(n2309), .I1(n30252), .CO(n23138));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n30252), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n30252), 
            .CO(n23137));
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n14736), 
            .D(n255[14]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n14736), 
            .D(n255[13]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n14736), 
            .D(n255[12]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n14736), 
            .D(n255[11]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n14736), 
            .D(n255[10]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n14736), 
            .D(n255[9]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n14736), 
            .D(n255[8]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n14736), 
            .D(n255[7]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n14736), 
            .D(n255[6]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n14736), 
            .D(n255[5]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n14736), 
            .D(n255[4]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n14736), 
            .D(n255[3]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n14736), 
            .D(n255[2]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1126_add_4_13 (.CI(n22343), .I0(GND_net), .I1(timer[11]), 
            .CO(n22344));
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n14736), 
            .D(n255[1]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25166_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30256));
    defparam i25166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4312));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4313));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1478 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4312), 
            .O(n16_adj_4314));
    defparam i7_4_lut_adj_1478.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16_adj_4314), .I2(n12_adj_4313), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1479 (.I0(bit_ctr[15]), .I1(n18), .I2(n2006), 
            .I3(n2009), .O(n25));
    defparam i9_4_lut_adj_1479.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1480 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n2027));
    defparam i15_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1126_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n22342), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25165_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30255));
    defparam i25165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1126_add_4_12 (.CI(n22342), .I0(GND_net), .I1(timer[10]), 
            .CO(n22343));
    SB_LUT4 timer_1126_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n22341), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_5 (.CI(n21907), .I0(bit_ctr[3]), .I1(GND_net), .CO(n21908));
    SB_LUT4 i15_4_lut_adj_1481 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_4315));
    defparam i15_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_4316));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1482 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_4317));
    defparam i17_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1483 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45));
    defparam i18_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1484 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_4318));
    defparam i16_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), .I3(GND_net), 
            .O(n40_adj_4319));
    defparam i13_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i21_4_lut (.I0(n3107), .I1(n42_adj_4315), .I2(n3087), .I3(n3086), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1485 (.I0(n43_adj_4318), .I1(n45), .I2(n44_adj_4317), 
            .I3(n46_adj_4316), .O(n52));
    defparam i25_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1486 (.I0(n3095), .I1(n3084), .I2(GND_net), 
            .I3(GND_net), .O(n39));
    defparam i12_2_lut_adj_1486.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut (.I0(n39), .I1(n52), .I2(n48), .I3(n40_adj_4319), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25164_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30254));
    defparam i25164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1126_add_4_11 (.CI(n22341), .I0(GND_net), .I1(timer[9]), 
            .CO(n22342));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n22265), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1126_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n22340), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n21914), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15163_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n18991));
    defparam i15163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n11_adj_4321), .I2(n29), .I3(n51), 
            .O(n48_adj_4322));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1487 (.I0(n37_adj_4323), .I1(n23), .I2(n53), 
            .I3(n39_adj_4324), .O(n46_adj_4325));
    defparam i18_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1488 (.I0(n27_adj_4326), .I1(n57), .I2(n63), 
            .I3(n43_adj_4327), .O(n47));
    defparam i19_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1489 (.I0(n25_adj_4328), .I1(n33), .I2(n47_adj_4329), 
            .I3(n61), .O(n45_adj_4330));
    defparam i17_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1490 (.I0(n59), .I1(n17_adj_4331), .I2(n15_adj_4332), 
            .I3(n55), .O(n44_adj_4333));
    defparam i16_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1491 (.I0(n31), .I1(n41_adj_4334), .I2(n49), 
            .I3(n18991), .O(n43_adj_4335));
    defparam i15_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1492 (.I0(n45_adj_4330), .I1(n47), .I2(n46_adj_4325), 
            .I3(n48_adj_4322), .O(n54));
    defparam i26_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1493 (.I0(n45_adj_4336), .I1(n13_adj_4337), .I2(n19_adj_4338), 
            .I3(n21), .O(n49_adj_4339));
    defparam i21_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4339), .I1(n54), .I2(n43_adj_4335), 
            .I3(n44_adj_4333), .O(n23352));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(bit_ctr[3]), .I1(n23352), .I2(GND_net), 
            .I3(GND_net), .O(n23676));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1495 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4340));
    defparam i7_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1496 (.I0(n1504), .I1(n18_adj_4340), .I2(n1502), 
            .I3(n1499), .O(n20));
    defparam i9_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), .I3(GND_net), 
            .O(n15_adj_4341));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1497 (.I0(n15_adj_4341), .I1(n20), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n22004), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_3_lut_adj_1498 (.I0(bit_ctr[6]), .I1(n2908), .I2(n2909), 
            .I3(GND_net), .O(n29_adj_4343));
    defparam i4_3_lut_adj_1498.LUT_INIT = 16'hecec;
    SB_LUT4 i14_4_lut_adj_1499 (.I0(n2900), .I1(n2895), .I2(n2901), .I3(n2906), 
            .O(n39_adj_4344));
    defparam i14_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1500 (.I0(n2891), .I1(n2896), .I2(n2889), .I3(GND_net), 
            .O(n38_adj_4345));
    defparam i13_3_lut_adj_1500.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1501 (.I0(n2897), .I1(n2899), .I2(n2887), .I3(n2892), 
            .O(n43_adj_4346));
    defparam i18_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1502 (.I0(n2905), .I1(n2903), .I2(n2888), .I3(n2907), 
            .O(n42_adj_4347));
    defparam i17_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1503 (.I0(n2898), .I1(n2886), .I2(n2893), .I3(n2904), 
            .O(n41_adj_4348));
    defparam i16_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1504 (.I0(n39_adj_4344), .I1(n29_adj_4343), .I2(n2890), 
            .I3(n2902), .O(n45_adj_4349));
    defparam i20_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43_adj_4346), .I1(n2894), .I2(n38_adj_4345), 
            .I3(n2885), .O(n47_adj_4350));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1505 (.I0(n47_adj_4350), .I1(n45_adj_4349), .I2(n41_adj_4348), 
            .I3(n42_adj_4347), .O(n2918));
    defparam i24_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i25169_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30259));
    defparam i25169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25170_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30260));
    defparam i25170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1506 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4351));
    defparam i1_2_lut_adj_1506.LUT_INIT = 16'heeee;
    SB_LUT4 i15171_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n18999));
    defparam i15171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4351), 
            .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1507 (.I0(n2098), .I1(n18999), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4352));
    defparam i11_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1508 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4353));
    defparam i12_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1509 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4354));
    defparam i10_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1510 (.I0(n27_adj_4354), .I1(n29_adj_4353), .I2(n28_adj_4352), 
            .I3(n30), .O(n2126));
    defparam i16_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n14736), 
            .D(n255[18]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_12 (.CI(n21914), .I0(bit_ctr[10]), .I1(GND_net), .CO(n21915));
    SB_CARRY mod_5_add_1272_12 (.CI(n22265), .I0(n1800), .I1(n1829), .CO(n22266));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n22264), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n21906), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_10 (.CI(n22340), .I0(GND_net), .I1(timer[8]), 
            .CO(n22341));
    SB_CARRY mod_5_add_1272_11 (.CI(n22264), .I0(n1801), .I1(n1829), .CO(n22265));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n22263), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n22004), .I0(n2201), .I1(n2225), .CO(n22005));
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n14736), 
            .D(n255[17]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n14736), 
            .D(n255[25]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n21913), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n14736), 
            .D(n255[24]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_11 (.CI(n21913), .I0(bit_ctr[9]), .I1(GND_net), .CO(n21914));
    SB_LUT4 timer_1126_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n22339), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n21906), .I0(bit_ctr[2]), .I1(GND_net), .CO(n21907));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n22003), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n22263), .I0(n1802), .I1(n1829), .CO(n22264));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n22262), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n22003), .I0(n2202), .I1(n2225), .CO(n22004));
    SB_LUT4 i25168_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30258));
    defparam i25168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n22002), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n22002), .I0(n2203), .I1(n2225), .CO(n22003));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n22001), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n22262), .I0(n1803), .I1(n1829), .CO(n22263));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n22261), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1126_add_4_9 (.CI(n22339), .I0(GND_net), .I1(timer[7]), 
            .CO(n22340));
    SB_CARRY mod_5_add_1272_8 (.CI(n22261), .I0(n1804), .I1(n1829), .CO(n22262));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n22260), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1126_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n22338), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n22001), .I0(n2204), .I1(n2225), .CO(n22002));
    SB_CARRY timer_1126_add_4_8 (.CI(n22338), .I0(GND_net), .I1(timer[6]), 
            .CO(n22339));
    SB_CARRY mod_5_add_1272_7 (.CI(n22260), .I0(n1805), .I1(n1829), .CO(n22261));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n22000), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n22259), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1126_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n22337), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n21935), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n14736), 
            .D(n255[16]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1272_6 (.CI(n22259), .I0(n1806), .I1(n1829), .CO(n22260));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n22258), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n22000), .I0(n2205), .I1(n2225), .CO(n22001));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n21999), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n22258), .I0(n1807), .I1(n1829), .CO(n22259));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n22257), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1126_add_4_7 (.CI(n22337), .I0(GND_net), .I1(timer[5]), 
            .CO(n22338));
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n21934), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1126_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n22336), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n21999), .I0(n2206), .I1(n2225), .CO(n22000));
    SB_CARRY timer_1126_add_4_6 (.CI(n22336), .I0(GND_net), .I1(timer[4]), 
            .CO(n22337));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n21998), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n22257), .I0(n1808), .I1(n1829), .CO(n22258));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n30250), 
            .I3(n22256), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_5 (.CI(n21998), .I0(n2207), .I1(n2225), .CO(n21999));
    SB_LUT4 i6_4_lut_adj_1511 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4355));
    defparam i6_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n9_adj_4356));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1512 (.I0(n9_adj_4356), .I1(n14_adj_4355), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n21997), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n21997), .I0(n2208), .I1(n2225), .CO(n21998));
    SB_LUT4 timer_1126_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n22335), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n22256), .I0(n1809), .I1(n30250), .CO(n22257));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n30251), 
            .I3(n21996), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1126_add_4_5 (.CI(n22335), .I0(GND_net), .I1(timer[3]), 
            .CO(n22336));
    SB_CARRY add_21_32 (.CI(n21934), .I0(bit_ctr[30]), .I1(GND_net), .CO(n21935));
    SB_LUT4 timer_1126_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n22334), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n21996), .I0(n2209), .I1(n30251), .CO(n21997));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n21933), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n30251), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n30250), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_31 (.CI(n21933), .I0(bit_ctr[29]), .I1(GND_net), .CO(n21934));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n21912), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n30251), 
            .CO(n21996));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n30250), 
            .CO(n22256));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n22255), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1126_add_4_4 (.CI(n22334), .I0(GND_net), .I1(timer[2]), 
            .CO(n22335));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n21932), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n21932), .I0(bit_ctr[28]), .I1(GND_net), .CO(n21933));
    SB_LUT4 timer_1126_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n22333), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n22254), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1126_add_4_3 (.CI(n22333), .I0(GND_net), .I1(timer[1]), 
            .CO(n22334));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n21931), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n22254), .I0(n1896), .I1(n1928), .CO(n22255));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n22253), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1126_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_10 (.CI(n21912), .I0(bit_ctr[8]), .I1(GND_net), .CO(n21913));
    SB_LUT4 i11_4_lut_adj_1513 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4358));
    defparam i11_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1514 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4359));
    defparam i4_3_lut_adj_1514.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4360));
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'heeee;
    SB_CARRY add_21_29 (.CI(n21931), .I0(bit_ctr[27]), .I1(GND_net), .CO(n21932));
    SB_LUT4 i9_4_lut_adj_1516 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24));
    defparam i9_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1517 (.I0(n19_adj_4359), .I1(n26_adj_4358), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4361));
    defparam i13_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1518 (.I0(n1896), .I1(n28_adj_4361), .I2(n24), 
            .I3(n16_adj_4360), .O(n1928));
    defparam i14_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n21905), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n22253), .I0(n1897), .I1(n1928), .CO(n22254));
    SB_LUT4 i25161_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30251));
    defparam i25161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n22252), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1126_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n22333));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n22332), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n22252), .I0(n1898), .I1(n1928), .CO(n22253));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n22251), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25160_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30250));
    defparam i25160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n22331), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n22251), .I0(n1899), .I1(n1928), .CO(n22252));
    SB_CARRY mod_5_add_870_9 (.CI(n22331), .I0(n1203), .I1(n1235), .CO(n22332));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n22250), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n22250), .I0(n1900), .I1(n1928), .CO(n22251));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n22249), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n22249), .I0(n1901), .I1(n1928), .CO(n22250));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n22248), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n22330), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n22248), .I0(n1902), .I1(n1928), .CO(n22249));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n22247), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n22247), .I0(n1903), .I1(n1928), .CO(n22248));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n22246), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n21911), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n22246), .I0(n1904), .I1(n1928), .CO(n22247));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n21930), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n22245), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n22245), .I0(n1905), .I1(n1928), .CO(n22246));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n22244), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_399[16]), .I1(timer[31]), 
            .I2(n56[31]), .I3(n22161), .O(n27_adj_4362)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_399[24]), .I1(timer[30]), 
            .I2(n56[30]), .I3(n22160), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1339_6 (.CI(n22244), .I0(n1906), .I1(n1928), .CO(n22245));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n22243), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_28 (.CI(n21930), .I0(bit_ctr[26]), .I1(GND_net), .CO(n21931));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n21929), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n21929), .I0(bit_ctr[25]), .I1(GND_net), .CO(n21930));
    SB_CARRY sub_14_add_2_32 (.CI(n22160), .I0(timer[30]), .I1(n56[30]), 
            .CO(n22161));
    SB_CARRY mod_5_add_870_8 (.CI(n22330), .I0(n1204), .I1(n1235), .CO(n22331));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_399[22]), .I1(timer[29]), 
            .I2(n56[29]), .I3(n22159), .O(n23_adj_4363)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n22159), .I0(timer[29]), .I1(n56[29]), 
            .CO(n22160));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_399[18]), .I1(timer[28]), 
            .I2(n56[28]), .I3(n22158), .O(n28_adj_4364)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1339_5 (.CI(n22243), .I0(n1907), .I1(n1928), .CO(n22244));
    SB_LUT4 i25162_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30252));
    defparam i25162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n21928), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_30 (.CI(n22158), .I0(timer[28]), .I1(n56[28]), 
            .CO(n22159));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n22329), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_399[25]), .I1(timer[27]), 
            .I2(n56[27]), .I3(n22157), .O(n26_adj_4365)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n22242), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4366));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1519 (.I0(bit_ctr[12]), .I1(n22_adj_4366), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4367));
    defparam i11_4_lut_adj_1519.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1520 (.I0(n2294), .I1(n30_adj_4367), .I2(n2306), 
            .I3(n2297), .O(n34));
    defparam i15_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1521 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32));
    defparam i13_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1522 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4368));
    defparam i14_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1523 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4369));
    defparam i12_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1524 (.I0(n31_adj_4369), .I1(n33_adj_4368), .I2(n32), 
            .I3(n34), .O(n2324));
    defparam i18_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1339_4 (.CI(n22242), .I0(n1908), .I1(n1928), .CO(n22243));
    SB_CARRY mod_5_add_870_7 (.CI(n22329), .I0(n1205), .I1(n1235), .CO(n22330));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n30254), 
            .I3(n22241), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10_4_lut_adj_1525 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4370));
    defparam i10_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1526 (.I0(n2203), .I1(n28_adj_4370), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4371));
    defparam i14_4_lut_adj_1526.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1527 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4372));
    defparam i12_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1528 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4373));
    defparam i13_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1529 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4374));
    defparam i11_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1530 (.I0(n29_adj_4374), .I1(n31_adj_4373), .I2(n30_adj_4372), 
            .I3(n32_adj_4371), .O(n2225));
    defparam i17_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n22328), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n22650), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n22649), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n22649), .I0(n3084), .I1(n3116), .CO(n22650));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n22648), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n22648), .I0(n3085), .I1(n3116), .CO(n22649));
    SB_LUT4 i19_4_lut_adj_1531 (.I0(bit_ctr[23]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46_adj_4375));   // verilog/neopixel.v(38[12:22])
    defparam i19_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1532 (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[25]), 
            .I3(bit_ctr[10]), .O(n44_adj_4376));   // verilog/neopixel.v(38[12:22])
    defparam i17_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1533 (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45_adj_4377));   // verilog/neopixel.v(38[12:22])
    defparam i18_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1534 (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43_adj_4378));   // verilog/neopixel.v(38[12:22])
    defparam i16_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1535 (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42_adj_4379));   // verilog/neopixel.v(38[12:22])
    defparam i15_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_3_lut (.I0(bit_ctr[26]), .I1(bit_ctr[13]), .I2(bit_ctr[22]), 
            .I3(GND_net), .O(n41_adj_4380));   // verilog/neopixel.v(38[12:22])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i25_4_lut_adj_1536 (.I0(n43_adj_4378), .I1(n45_adj_4377), .I2(n44_adj_4376), 
            .I3(n46_adj_4375), .O(n52_adj_4381));   // verilog/neopixel.v(38[12:22])
    defparam i25_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1537 (.I0(bit_ctr[30]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[8]), .O(n47_adj_4382));   // verilog/neopixel.v(38[12:22])
    defparam i20_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1538 (.I0(n47_adj_4382), .I1(n52_adj_4381), .I2(n41_adj_4380), 
            .I3(n42_adj_4379), .O(n11306));   // verilog/neopixel.v(38[12:22])
    defparam i26_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i16759_4_lut (.I0(start), .I1(n28371), .I2(\state[0] ), .I3(n20565), 
            .O(n33_adj_4383));   // verilog/neopixel.v(16[20:25])
    defparam i16759_4_lut.LUT_INIT = 16'h4540;
    SB_LUT4 i1_2_lut_adj_1539 (.I0(\neo_pixel_transmitter.done ), .I1(n33_adj_4383), 
            .I2(GND_net), .I3(GND_net), .O(n20572));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1539.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(start), .I1(n20565), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n6_adj_4384));   // verilog/neopixel.v(16[20:25])
    defparam i2_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i11031_4_lut (.I0(n14736), .I1(\neo_pixel_transmitter.done ), 
            .I2(n6_adj_4384), .I3(n28371), .O(n14862));   // verilog/neopixel.v(35[12] 117[6])
    defparam i11031_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n22647), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_26 (.CI(n21928), .I0(bit_ctr[24]), .I1(GND_net), .CO(n21929));
    SB_CARRY sub_14_add_2_29 (.CI(n22157), .I0(timer[27]), .I1(n56[27]), 
            .CO(n22158));
    SB_CARRY mod_5_add_2143_26 (.CI(n22647), .I0(n3086), .I1(n3116), .CO(n22648));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n22646), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n22646), .I0(n3087), .I1(n3116), .CO(n22647));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n21927), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n22645), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n22645), .I0(n3088), .I1(n3116), .CO(n22646));
    SB_CARRY mod_5_add_1339_3 (.CI(n22241), .I0(n1909), .I1(n30254), .CO(n22242));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n22644), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_2143_23 (.CI(n22644), .I0(n3089), .I1(n3116), .CO(n22645));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n22643), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n22643), .I0(n3090), .I1(n3116), .CO(n22644));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n22642), .O(n47_adj_4329)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n22642), .I0(n3091), .I1(n3116), .CO(n22643));
    SB_LUT4 i24467_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n20610), 
            .I3(GND_net), .O(n29293));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24467_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_DFF timer_1126__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i1_2_lut_3_lut (.I0(n13644), .I1(one_wire_N_399[9]), .I2(n1), 
            .I3(GND_net), .O(n107));   // verilog/neopixel.v(53[15:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i16763_4_lut (.I0(n20572), .I1(n29274), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n14736));   // verilog/neopixel.v(16[20:25])
    defparam i16763_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n22641), .O(n45_adj_4336)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut (.I0(n13644), .I1(one_wire_N_399[9]), .I2(n26721), 
            .I3(n1), .O(n26806));   // verilog/neopixel.v(53[15:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_20 (.CI(n22641), .I0(n3092), .I1(n3116), .CO(n22642));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n22640), .O(n43_adj_4327)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n22328), .I0(n1206), .I1(n1235), .CO(n22329));
    SB_CARRY mod_5_add_2143_19 (.CI(n22640), .I0(n3093), .I1(n3116), .CO(n22641));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n22639), .O(n41_adj_4334)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n22639), .I0(n3094), .I1(n3116), .CO(n22640));
    SB_LUT4 sub_14_add_2_28_lut (.I0(one_wire_N_399[17]), .I1(timer[26]), 
            .I2(n56[26]), .I3(n22156), .O(n21_adj_4386)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n22327), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n30254), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_5 (.CI(n22327), .I0(n1207), .I1(n1235), .CO(n22328));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n22326), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n22638), .O(n39_adj_4324)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n22638), .I0(n3095), .I1(n3116), .CO(n22639));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n22637), .O(n37_adj_4323)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n22326), .I0(n1208), .I1(n1235), .CO(n22327));
    SB_CARRY mod_5_add_2143_16 (.CI(n22637), .I0(n3096), .I1(n3116), .CO(n22638));
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n30254), 
            .CO(n22241));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n30255), 
            .I3(n22325), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n22636), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_28 (.CI(n22156), .I0(timer[26]), .I1(n56[26]), 
            .CO(n22157));
    SB_CARRY mod_5_add_2143_15 (.CI(n22636), .I0(n3097), .I1(n3116), .CO(n22637));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n22635), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_3 (.CI(n22325), .I0(n1209), .I1(n30255), .CO(n22326));
    SB_CARRY mod_5_add_2143_14 (.CI(n22635), .I0(n3098), .I1(n3116), .CO(n22636));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n22634), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n22634), .I0(n3099), .I1(n3116), .CO(n22635));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n22240), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n30255), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n22633), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n22633), .I0(n3100), .I1(n3116), .CO(n22634));
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n30255), 
            .CO(n22325));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n22324), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n22239), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n22323), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n22323), .I0(n1302), .I1(n1334), .CO(n22324));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n56[25]), 
            .I3(n22155), .O(one_wire_N_399[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n22322), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n22239), .I0(n1995), .I1(n2027), .CO(n22240));
    SB_CARRY mod_5_add_937_9 (.CI(n22322), .I0(n1303), .I1(n1334), .CO(n22323));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n22321), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n22321), .I0(n1304), .I1(n1334), .CO(n22322));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n22238), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n22238), .I0(n1996), .I1(n2027), .CO(n22239));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n22632), .O(n27_adj_4326)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n22632), .I0(n3101), .I1(n3116), .CO(n22633));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n22631), .O(n25_adj_4328)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n22631), .I0(n3102), .I1(n3116), .CO(n22632));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n22630), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25180_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30270));
    defparam i25180_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25125_2_lut (.I0(n2_adj_4387), .I1(n971[28]), .I2(GND_net), 
            .I3(GND_net), .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i25125_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25123_2_lut (.I0(n2_adj_4387), .I1(n971[29]), .I2(GND_net), 
            .I3(GND_net), .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i25123_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2_adj_4387), 
            .I3(GND_net), .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut_adj_1541 (.I0(n14818), .I1(n905), .I2(n26696), .I3(GND_net), 
            .O(n8_adj_4388));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1541.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n8_adj_4388), .I2(n906), .I3(n12170), 
            .O(n2_adj_4387));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h040c;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2_adj_4387), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n12170), .I1(n971[27]), .I2(n2_adj_4387), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY mod_5_add_2143_9 (.CI(n22630), .I0(n3103), .I1(n3116), .CO(n22631));
    SB_CARRY sub_14_add_2_27 (.CI(n22155), .I0(timer[25]), .I1(n56[25]), 
            .CO(n22156));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n22629), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n56[24]), 
            .I3(n22154), .O(one_wire_N_399[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23295_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n28385));
    defparam i23295_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n22320), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n22320), .I0(n1305), .I1(n1334), .CO(n22321));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n22319), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_26 (.CI(n22154), .I0(timer[24]), .I1(n56[24]), 
            .CO(n22155));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n22237), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n22629), .I0(n3104), .I1(n3116), .CO(n22630));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n22628), .O(n19_adj_4338)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n22628), .I0(n3105), .I1(n3116), .CO(n22629));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n22627), .O(n17_adj_4331)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6_adj_4389));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_937_6 (.CI(n22319), .I0(n1306), .I1(n1334), .CO(n22320));
    SB_CARRY mod_5_add_1406_15 (.CI(n22237), .I0(n1997), .I1(n2027), .CO(n22238));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n22236), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n22627), .I0(n3106), .I1(n3116), .CO(n22628));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n22626), .O(n15_adj_4332)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n22626), .I0(n3107), .I1(n3116), .CO(n22627));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n22625), .O(n13_adj_4337)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n22625), .I0(n3108), .I1(n3116), .CO(n22626));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n30256), 
            .I3(n22624), .O(n11_adj_4321)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n22624), .I0(n3109), .I1(n30256), .CO(n22625));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n30256), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_4_lut (.I0(n2_adj_4387), .I1(n6_adj_4389), .I2(n1005), 
            .I3(n28385), .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i3_4_lut_4_lut (.I0(n26662), .I1(n11764), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i25146_2_lut (.I0(n2_adj_4387), .I1(n971[31]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4390));   // verilog/neopixel.v(22[26:36])
    defparam i25146_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25045_3_lut_4_lut (.I0(n11764), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n26662), .O(n26696));   // verilog/neopixel.v(22[26:36])
    defparam i25045_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i1_2_lut_adj_1542 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n12170));
    defparam i1_2_lut_adj_1542.LUT_INIT = 16'h9999;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_399[14]), .I1(timer[23]), 
            .I2(n56[23]), .I3(n22153), .O(n29_adj_4391)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n30256), 
            .CO(n22624));
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY sub_14_add_2_25 (.CI(n22153), .I0(timer[23]), .I1(n56[23]), 
            .CO(n22154));
    SB_CARRY add_21_9 (.CI(n21911), .I0(bit_ctr[7]), .I1(GND_net), .CO(n21912));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n22318), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n22318), .I0(n1307), .I1(n1334), .CO(n22319));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n22623), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n22236), .I0(n1998), .I1(n2027), .CO(n22237));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n22317), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n22235), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n56[22]), 
            .I3(n22152), .O(one_wire_N_399[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n22317), .I0(n1308), .I1(n1334), .CO(n22318));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n30257), 
            .I3(n22316), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n22316), .I0(n1309), .I1(n30257), .CO(n22317));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n30257), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_13 (.CI(n22235), .I0(n1999), .I1(n2027), .CO(n22236));
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n30257), 
            .CO(n22316));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n22622), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n22622), .I0(n2985), .I1(n3017), .CO(n22623));
    SB_CARRY sub_14_add_2_24 (.CI(n22152), .I0(timer[22]), .I1(n56[22]), 
            .CO(n22153));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n22621), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n22621), .I0(n2986), .I1(n3017), .CO(n22622));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n22620), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n22620), .I0(n2987), .I1(n3017), .CO(n22621));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n22619), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n22619), .I0(n2988), .I1(n3017), .CO(n22620));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n22618), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n22618), .I0(n2989), .I1(n3017), .CO(n22619));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n22617), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n22617), .I0(n2990), .I1(n3017), .CO(n22618));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n22616), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n22616), .I0(n2991), .I1(n3017), .CO(n22617));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n22615), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n22615), .I0(n2992), .I1(n3017), .CO(n22616));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n22614), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n22614), .I0(n2993), .I1(n3017), .CO(n22615));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n22613), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n22234), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n22613), .I0(n2994), .I1(n3017), .CO(n22614));
    SB_CARRY mod_5_add_1406_12 (.CI(n22234), .I0(n2000), .I1(n2027), .CO(n22235));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n22612), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_399[15]), .I1(timer[21]), 
            .I2(n56[21]), .I3(n22151), .O(n30_adj_4392)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n22233), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n22315), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15133_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i15133_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n22314), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n22233), .I0(n2001), .I1(n2027), .CO(n22234));
    SB_CARRY sub_14_add_2_23 (.CI(n22151), .I0(timer[21]), .I1(n56[21]), 
            .CO(n22152));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n22232), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n22232), .I0(n2002), .I1(n2027), .CO(n22233));
    SB_CARRY mod_5_add_2076_17 (.CI(n22612), .I0(n2995), .I1(n3017), .CO(n22613));
    SB_LUT4 i2_4_lut_adj_1543 (.I0(n708), .I1(n18738), .I2(n26710), .I3(n608), 
            .O(n26798));
    defparam i2_4_lut_adj_1543.LUT_INIT = 16'hfefa;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n22611), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n22611), .I0(n2996), .I1(n3017), .CO(n22612));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n22610), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n22610), .I0(n2997), .I1(n3017), .CO(n22611));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n22609), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n22609), .I0(n2998), .I1(n3017), .CO(n22610));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n22608), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n22608), .I0(n2999), .I1(n3017), .CO(n22609));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n22607), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1544 (.I0(bit_ctr[28]), .I1(n26798), .I2(GND_net), 
            .I3(GND_net), .O(n11764));
    defparam i1_2_lut_adj_1544.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n22231), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n22607), .I0(n3000), .I1(n3017), .CO(n22608));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n22606), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n22606), .I0(n3001), .I1(n3017), .CO(n22607));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n22605), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24228_3_lut (.I0(n23680), .I1(bit_ctr[28]), .I2(n26798), 
            .I3(GND_net), .O(n26662));
    defparam i24228_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i23222_3_lut (.I0(n26798), .I1(n708), .I2(n26710), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i23222_3_lut.LUT_INIT = 16'h8282;
    SB_CARRY mod_5_add_2076_10 (.CI(n22605), .I0(n3002), .I1(n3017), .CO(n22606));
    SB_CARRY mod_5_add_1004_11 (.CI(n22314), .I0(n1401), .I1(n1433), .CO(n22315));
    SB_CARRY mod_5_add_1406_9 (.CI(n22231), .I0(n2003), .I1(n2027), .CO(n22232));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_399[12]), .I1(timer[20]), 
            .I2(n56[20]), .I3(n22150), .O(n24_adj_4393)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n22230), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n22230), .I0(n2004), .I1(n2027), .CO(n22231));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n22313), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n21927), .I0(bit_ctr[23]), .I1(GND_net), .CO(n21928));
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n22229), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25179_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30269));
    defparam i25179_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), .I3(GND_net), 
            .O(n27_adj_4394));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1406_7 (.CI(n22229), .I0(n2005), .I1(n2027), .CO(n22230));
    SB_CARRY mod_5_add_1004_10 (.CI(n22313), .I0(n1402), .I1(n1433), .CO(n22314));
    SB_LUT4 i13_4_lut_adj_1545 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4395));
    defparam i13_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1546 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4396));
    defparam i12_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1547 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4397));
    defparam i11_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1548 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4398));
    defparam i15_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1549 (.I0(n33_adj_4395), .I1(n27_adj_4394), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4399));
    defparam i17_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1550 (.I0(n37_adj_4399), .I1(n35_adj_4398), .I2(n31_adj_4397), 
            .I3(n32_adj_4396), .O(n2423));
    defparam i19_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i25178_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30268));
    defparam i25178_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n22312), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n22228), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n22150), .I0(timer[20]), .I1(n56[20]), 
            .CO(n22151));
    SB_CARRY mod_5_add_1406_6 (.CI(n22228), .I0(n2006), .I1(n2027), .CO(n22229));
    SB_LUT4 sub_14_add_2_21_lut (.I0(one_wire_N_399[13]), .I1(timer[19]), 
            .I2(n56[19]), .I3(n22149), .O(n25_adj_4400)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1004_9 (.CI(n22312), .I0(n1403), .I1(n1433), .CO(n22313));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n22311), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n22227), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_21 (.CI(n22149), .I0(timer[19]), .I1(n56[19]), 
            .CO(n22150));
    SB_CARRY mod_5_add_1004_8 (.CI(n22311), .I0(n1404), .I1(n1433), .CO(n22312));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n56[18]), 
            .I3(n22148), .O(one_wire_N_399[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n22227), .I0(n2007), .I1(n2027), .CO(n22228));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n22310), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n22226), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n22310), .I0(n1405), .I1(n1433), .CO(n22311));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n22309), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n22226), .I0(n2008), .I1(n2027), .CO(n22227));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n30258), 
            .I3(n22225), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_20 (.CI(n22148), .I0(timer[18]), .I1(n56[18]), 
            .CO(n22149));
    SB_CARRY mod_5_add_1004_6 (.CI(n22309), .I0(n1406), .I1(n1433), .CO(n22310));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n22308), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n56[17]), 
            .I3(n22147), .O(one_wire_N_399[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_5 (.CI(n22308), .I0(n1407), .I1(n1433), .CO(n22309));
    SB_CARRY mod_5_add_1406_3 (.CI(n22225), .I0(n2009), .I1(n30258), .CO(n22226));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n30258), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n30258), 
            .CO(n22225));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n22604), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n22604), .I0(n3003), .I1(n3017), .CO(n22605));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n22603), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n22307), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n22603), .I0(n3004), .I1(n3017), .CO(n22604));
    SB_CARRY mod_5_add_1004_4 (.CI(n22307), .I0(n1408), .I1(n1433), .CO(n22308));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n22602), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut_adj_1551 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4401));
    defparam i3_2_lut_adj_1551.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut_adj_1552 (.I0(n21_adj_4386), .I1(n23_adj_4363), .I2(n22), 
            .I3(n24_adj_4393), .O(n36));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1553 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4402));
    defparam i13_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1554 (.I0(n25_adj_4400), .I1(n27_adj_4362), .I2(n26_adj_4365), 
            .I3(n28_adj_4364), .O(n37_adj_4403));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1555 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4404));
    defparam i1_3_lut_adj_1555.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1556 (.I0(n2490), .I1(n34_adj_4402), .I2(n24_adj_4401), 
            .I3(n2494), .O(n38_adj_4405));
    defparam i17_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1557 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4406));
    defparam i15_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1558 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4404), 
            .O(n37_adj_4407));
    defparam i16_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1559 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4408));
    defparam i14_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1560 (.I0(n35_adj_4408), .I1(n37_adj_4407), .I2(n36_adj_4406), 
            .I3(n38_adj_4405), .O(n2522));
    defparam i20_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i25176_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30266));
    defparam i25176_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16770_4_lut (.I0(n26721), .I1(n27279), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n28317));   // verilog/neopixel.v(16[20:25])
    defparam i16770_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(start), .I2(n107), .I3(n28317), 
            .O(n1554));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n30568));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30568_bdd_4_lut (.I0(n30568), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n28389));
    defparam n30568_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n22224), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n22602), .I0(n3005), .I1(n3017), .CO(n22603));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n22223), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n22601), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n22147), .I0(timer[17]), .I1(n56[17]), 
            .CO(n22148));
    SB_CARRY mod_5_add_1473_18 (.CI(n22223), .I0(n2094), .I1(n2126), .CO(n22224));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n30260), 
            .I3(n22306), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n22222), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n22222), .I0(n2095), .I1(n2126), .CO(n22223));
    SB_CARRY mod_5_add_1004_3 (.CI(n22306), .I0(n1409), .I1(n30260), .CO(n22307));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n21926), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_6 (.CI(n22601), .I0(n3006), .I1(n3017), .CO(n22602));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n22600), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n22600), .I0(n3007), .I1(n3017), .CO(n22601));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n22599), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n22599), .I0(n3008), .I1(n3017), .CO(n22600));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n30259), 
            .I3(n22598), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n22598), .I0(n3009), .I1(n30259), .CO(n22599));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n30259), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25425 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n30478));
    defparam bit_ctr_0__bdd_4_lut_25425.LUT_INIT = 16'he4aa;
    SB_LUT4 n30478_bdd_4_lut (.I0(n30478), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n30481));
    defparam n30478_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n30259), 
            .CO(n22598));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n22597), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n22596), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n22221), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n22596), .I0(n2886), .I1(n2918), .CO(n22597));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n22595), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n22595), .I0(n2887), .I1(n2918), .CO(n22596));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n22594), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n22594), .I0(n2888), .I1(n2918), .CO(n22595));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n22593), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n22593), .I0(n2889), .I1(n2918), .CO(n22594));
    SB_CARRY mod_5_add_1473_16 (.CI(n22221), .I0(n2096), .I1(n2126), .CO(n22222));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n22220), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25351 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n30424));
    defparam bit_ctr_0__bdd_4_lut_25351.LUT_INIT = 16'he4aa;
    SB_LUT4 n30424_bdd_4_lut (.I0(n30424), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n28518));
    defparam n30424_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25306 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n30418));
    defparam bit_ctr_0__bdd_4_lut_25306.LUT_INIT = 16'he4aa;
    SB_LUT4 n30418_bdd_4_lut (.I0(n30418), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n28521));
    defparam n30418_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25301 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n30406));
    defparam bit_ctr_0__bdd_4_lut_25301.LUT_INIT = 16'he4aa;
    SB_LUT4 n30406_bdd_4_lut (.I0(n30406), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n30409));
    defparam n30406_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY mod_5_add_1473_15 (.CI(n22220), .I0(n2097), .I1(n2126), .CO(n22221));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n30260), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n56[16]), 
            .I3(n22146), .O(one_wire_N_399[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n30260), 
            .CO(n22306));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n22592), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_18 (.CI(n22146), .I0(timer[16]), .I1(n56[16]), 
            .CO(n22147));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n22305), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 bit_ctr_0__bdd_4_lut_25291 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n30388));
    defparam bit_ctr_0__bdd_4_lut_25291.LUT_INIT = 16'he4aa;
    SB_LUT4 n30388_bdd_4_lut (.I0(n30388), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n29915));
    defparam n30388_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n28518), .I2(n28521), 
            .I3(n23676), .O(n30382));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30382_bdd_4_lut (.I0(n30382), .I1(n29915), .I2(n28389), .I3(n23676), 
            .O(n30385));
    defparam n30382_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n22219), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n56[15]), 
            .I3(n22145), .O(one_wire_N_399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_22 (.CI(n22592), .I0(n2890), .I1(n2918), .CO(n22593));
    SB_CARRY mod_5_add_1473_14 (.CI(n22219), .I0(n2098), .I1(n2126), .CO(n22220));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n22218), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_17 (.CI(n22145), .I0(timer[15]), .I1(n56[15]), 
            .CO(n22146));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n22304), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n22304), .I0(n1500), .I1(n1532), .CO(n22305));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n56[14]), 
            .I3(n22144), .O(one_wire_N_399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n22303), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n22218), .I0(n2099), .I1(n2126), .CO(n22219));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n22591), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n22591), .I0(n2891), .I1(n2918), .CO(n22592));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n22590), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n22590), .I0(n2892), .I1(n2918), .CO(n22591));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n22589), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n22589), .I0(n2893), .I1(n2918), .CO(n22590));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n22588), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n22588), .I0(n2894), .I1(n2918), .CO(n22589));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n22587), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n22587), .I0(n2895), .I1(n2918), .CO(n22588));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n22586), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n22586), .I0(n2896), .I1(n2918), .CO(n22587));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n22585), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n22585), .I0(n2897), .I1(n2918), .CO(n22586));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n22584), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19_4_lut_adj_1561 (.I0(n37_adj_4403), .I1(n29_adj_4391), .I2(n36), 
            .I3(n30_adj_4392), .O(n13644));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_14 (.CI(n22584), .I0(n2898), .I1(n2918), .CO(n22585));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n22583), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n22583), .I0(n2899), .I1(n2918), .CO(n22584));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n22582), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n22217), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n22303), .I0(n1501), .I1(n1532), .CO(n22304));
    SB_LUT4 i5_3_lut (.I0(n9_adj_4413), .I1(n7_adj_4414), .I2(n8_adj_4415), 
            .I3(GND_net), .O(n1));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1473_12 (.CI(n22217), .I0(n2100), .I1(n2126), .CO(n22218));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_12 (.CI(n22582), .I0(n2900), .I1(n2918), .CO(n22583));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n22581), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_adj_1562 (.I0(one_wire_N_399[2]), .I1(one_wire_N_399[4]), 
            .I2(one_wire_N_399[3]), .I3(GND_net), .O(n27279));   // verilog/neopixel.v(6[16:24])
    defparam i2_3_lut_adj_1562.LUT_INIT = 16'h8080;
    SB_CARRY mod_5_add_2009_11 (.CI(n22581), .I0(n2901), .I1(n2918), .CO(n22582));
    SB_LUT4 i21643_3_lut (.I0(one_wire_N_399[4]), .I1(n27201), .I2(one_wire_N_399[3]), 
            .I3(GND_net), .O(n26721));
    defparam i21643_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n22580), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i23283_2_lut (.I0(n107), .I1(n26721), .I2(GND_net), .I3(GND_net), 
            .O(n28371));
    defparam i23283_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1563 (.I0(n27279), .I1(n107), .I2(GND_net), .I3(GND_net), 
            .O(n20565));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut_adj_1563.LUT_INIT = 16'heeee;
    SB_LUT4 i21649_2_lut (.I0(\state[1] ), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n26727));
    defparam i21649_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_2009_10 (.CI(n22580), .I0(n2902), .I1(n2918), .CO(n22581));
    SB_LUT4 i1_4_lut_adj_1564 (.I0(n20565), .I1(n28371), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n33_adj_4417));
    defparam i1_4_lut_adj_1564.LUT_INIT = 16'h3553;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n22579), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n22579), .I0(n2903), .I1(n2918), .CO(n22580));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n22216), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25148_2_lut (.I0(n33_adj_4417), .I1(n26727), .I2(GND_net), 
            .I3(GND_net), .O(n25967));
    defparam i25148_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n22578), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1565 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4418));
    defparam i14_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1566 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4419));
    defparam i3_3_lut_adj_1566.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1567 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4420));
    defparam i12_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1568 (.I0(n25_adj_4419), .I1(n36_adj_4418), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4421));
    defparam i18_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1569 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4422));
    defparam i16_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4420), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4423));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1570 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4424));
    defparam i15_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_8 (.CI(n22578), .I0(n2904), .I1(n2918), .CO(n22579));
    SB_LUT4 i21_4_lut_adj_1571 (.I0(n37_adj_4424), .I1(n39_adj_4423), .I2(n38_adj_4422), 
            .I3(n40_adj_4421), .O(n2621));
    defparam i21_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1572 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4425));
    defparam i8_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1573 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4426));
    defparam i1_3_lut_adj_1573.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4427));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1574 (.I0(n13_adj_4426), .I1(n20_adj_4425), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4428));
    defparam i10_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1575 (.I0(n1601), .I1(n22_adj_4428), .I2(n18_adj_4427), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n22577), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n22577), .I0(n2905), .I1(n2918), .CO(n22578));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n22576), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25175_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30265));
    defparam i25175_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n14736), 
            .D(n255[0]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_6 (.CI(n22576), .I0(n2906), .I1(n2918), .CO(n22577));
    SB_CARRY mod_5_add_1473_11 (.CI(n22216), .I0(n2101), .I1(n2126), .CO(n22217));
    SB_CARRY sub_14_add_2_16 (.CI(n22144), .I0(timer[14]), .I1(n56[14]), 
            .CO(n22145));
    SB_LUT4 i16817_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_456 ));   // verilog/neopixel.v(16[20:25])
    defparam i16817_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n22215), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n22575), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n22575), .I0(n2907), .I1(n2918), .CO(n22576));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n22574), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n22574), .I0(n2908), .I1(n2918), .CO(n22575));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n22302), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut_adj_1576 (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(color_bit), 
            .I3(n11306), .O(state_3__N_248[0]));
    defparam i2_3_lut_4_lut_adj_1576.LUT_INIT = 16'h0070;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n11306), 
            .I3(GND_net), .O(n20573));
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'hf8f8;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1071_10 (.CI(n22302), .I0(n1502), .I1(n1532), .CO(n22303));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n56[13]), 
            .I3(n22143), .O(one_wire_N_399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n22215), .I0(n2102), .I1(n2126), .CO(n22216));
    SB_LUT4 i25173_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30263));
    defparam i25173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n30262), 
            .I3(n22573), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_15 (.CI(n22143), .I0(timer[13]), .I1(n56[13]), 
            .CO(n22144));
    SB_CARRY mod_5_add_2009_3 (.CI(n22573), .I0(n2909), .I1(n30262), .CO(n22574));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n30262), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n30262), 
            .CO(n22573));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n22572), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_24 (.CI(n21926), .I0(bit_ctr[22]), .I1(GND_net), .CO(n21927));
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n22571), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n21925), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_25 (.CI(n22571), .I0(n2787), .I1(n2819), .CO(n22572));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n22570), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n22570), .I0(n2788), .I1(n2819), .CO(n22571));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n22569), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n22301), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n22214), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n22569), .I0(n2789), .I1(n2819), .CO(n22570));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n22568), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n22568), .I0(n2790), .I1(n2819), .CO(n22569));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n22567), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n22214), .I0(n2103), .I1(n2126), .CO(n22215));
    SB_CARRY mod_5_add_1071_9 (.CI(n22301), .I0(n1503), .I1(n1532), .CO(n22302));
    SB_CARRY mod_5_add_1942_21 (.CI(n22567), .I0(n2791), .I1(n2819), .CO(n22568));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n22300), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n22213), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25171_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30261));
    defparam i25171_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_23 (.CI(n21925), .I0(bit_ctr[21]), .I1(GND_net), .CO(n21926));
    SB_CARRY mod_5_add_1473_8 (.CI(n22213), .I0(n2104), .I1(n2126), .CO(n22214));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n56[12]), 
            .I3(n22142), .O(one_wire_N_399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n22566), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n22300), .I0(n1504), .I1(n1532), .CO(n22301));
    SB_CARRY mod_5_add_1942_20 (.CI(n22566), .I0(n2792), .I1(n2819), .CO(n22567));
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n22299), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n22299), .I0(n1505), .I1(n1532), .CO(n22300));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n22212), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n22565), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n22565), .I0(n2793), .I1(n2819), .CO(n22566));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n22564), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_18 (.CI(n22564), .I0(n2794), .I1(n2819), .CO(n22565));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n22563), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n22563), .I0(n2795), .I1(n2819), .CO(n22564));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n22562), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_14 (.CI(n22142), .I0(timer[12]), .I1(n56[12]), 
            .CO(n22143));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n21924), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n22212), .I0(n2105), .I1(n2126), .CO(n22213));
    SB_CARRY mod_5_add_1942_16 (.CI(n22562), .I0(n2796), .I1(n2819), .CO(n22563));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n22561), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n22561), .I0(n2797), .I1(n2819), .CO(n22562));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n22211), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n22560), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n22211), .I0(n2106), .I1(n2126), .CO(n22212));
    SB_CARRY add_21_22 (.CI(n21924), .I0(bit_ctr[20]), .I1(GND_net), .CO(n21925));
    SB_CARRY mod_5_add_1942_14 (.CI(n22560), .I0(n2798), .I1(n2819), .CO(n22561));
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4435));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n22559), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n56[11]), 
            .I3(n22141), .O(one_wire_N_399[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n22298), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1578 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4437));
    defparam i15_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_13 (.CI(n22559), .I0(n2799), .I1(n2819), .CO(n22560));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n22558), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n22210), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15177_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n19005));
    defparam i15177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1579 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n19005), 
            .O(n36_adj_4438));
    defparam i13_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_12 (.CI(n22558), .I0(n2800), .I1(n2819), .CO(n22559));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n22557), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_13 (.CI(n22141), .I0(timer[11]), .I1(n56[11]), 
            .CO(n22142));
    SB_LUT4 i19_4_lut_adj_1580 (.I0(n2700), .I1(n38_adj_4437), .I2(n28_adj_4435), 
            .I3(n2705), .O(n42_adj_4439));
    defparam i19_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1581 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4440));
    defparam i17_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1071_6 (.CI(n22298), .I0(n1506), .I1(n1532), .CO(n22299));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n22297), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1582 (.I0(n2687), .I1(n36_adj_4438), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4441));
    defparam i18_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_11 (.CI(n22557), .I0(n2801), .I1(n2819), .CO(n22558));
    SB_CARRY mod_5_add_1071_5 (.CI(n22297), .I0(n1507), .I1(n1532), .CO(n22298));
    SB_LUT4 i16_4_lut_adj_1583 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4442));
    defparam i16_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n22296), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n22556), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i22_4_lut_adj_1584 (.I0(n39_adj_4442), .I1(n41_adj_4441), .I2(n40_adj_4440), 
            .I3(n42_adj_4439), .O(n2720));
    defparam i22_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_10 (.CI(n22556), .I0(n2802), .I1(n2819), .CO(n22557));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n21923), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n22555), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25174_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30264));
    defparam i25174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1585 (.I0(\neo_pixel_transmitter.done ), .I1(n20610), 
            .I2(GND_net), .I3(GND_net), .O(n20611));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'h4444;
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n21910), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n13644), .I1(one_wire_N_399[11]), .I2(one_wire_N_399[9]), 
            .I3(one_wire_N_399[10]), .O(n20610));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'heeea;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n56[10]), 
            .I3(n22140), .O(one_wire_N_399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n7_adj_4445), 
            .D(state_3__N_248[0]), .S(n20561));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_12 (.CI(n22140), .I0(timer[10]), .I1(n56[10]), 
            .CO(n22141));
    SB_CARRY mod_5_add_1942_9 (.CI(n22555), .I0(n2803), .I1(n2819), .CO(n22556));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n22554), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n22554), .I0(n2804), .I1(n2819), .CO(n22555));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n56[9]), 
            .I3(n22139), .O(one_wire_N_399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n22553), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n22553), .I0(n2805), .I1(n2819), .CO(n22554));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n22552), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n22552), .I0(n2806), .I1(n2819), .CO(n22553));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n22551), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n22551), .I0(n2807), .I1(n2819), .CO(n22552));
    SB_LUT4 i23_4_lut (.I0(n29293), .I1(n33_adj_4383), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n20561));   // verilog/neopixel.v(16[20:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n22550), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n22550), .I0(n2808), .I1(n2819), .CO(n22551));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n30264), 
            .I3(n22549), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_5 (.CI(n22210), .I0(n2107), .I1(n2126), .CO(n22211));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n22209), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_3 (.CI(n22549), .I0(n2809), .I1(n30264), .CO(n22550));
    SB_CARRY mod_5_add_1473_4 (.CI(n22209), .I0(n2108), .I1(n2126), .CO(n22210));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n30264), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_11 (.CI(n22139), .I0(timer[9]), .I1(n56[9]), 
            .CO(n22140));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n30264), 
            .CO(n22549));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n22548), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n22547), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_399[11]), .I1(timer[8]), 
            .I2(n56[8]), .I3(n22138), .O(n7_adj_4414)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_24 (.CI(n22547), .I0(n2688), .I1(n2720), .CO(n22548));
    SB_CARRY sub_14_add_2_10 (.CI(n22138), .I0(timer[8]), .I1(n56[8]), 
            .CO(n22139));
    SB_LUT4 sub_14_add_2_9_lut (.I0(one_wire_N_399[5]), .I1(timer[7]), .I2(n56[7]), 
            .I3(n22137), .O(n8_adj_4415)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n30261), 
            .I3(n22208), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n22546), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n22546), .I0(n2689), .I1(n2720), .CO(n22547));
    SB_LUT4 i15_4_lut_adj_1587 (.I0(n20572), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n20611), .O(n7_adj_4445));
    defparam i15_4_lut_adj_1587.LUT_INIT = 16'hfaca;
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n22545), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i2239_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n23352), 
            .I3(GND_net), .O(color_bit_N_442[4]));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2239_3_lut.LUT_INIT = 16'h6a6a;
    SB_CARRY mod_5_add_1875_22 (.CI(n22545), .I0(n2690), .I1(n2720), .CO(n22546));
    SB_CARRY mod_5_add_1473_3 (.CI(n22208), .I0(n2109), .I1(n30261), .CO(n22209));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n22544), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n22544), .I0(n2691), .I1(n2720), .CO(n22545));
    SB_LUT4 i1541971_i1_3_lut (.I0(n30481), .I1(n30409), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n22_adj_4446));
    defparam i1541971_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 color_bit_I_0_i31_4_lut (.I0(n30385), .I1(n22_adj_4446), .I2(color_bit_N_442[4]), 
            .I3(n23676), .O(color_bit));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n22543), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_9 (.CI(n22137), .I0(timer[7]), .I1(n56[7]), 
            .CO(n22138));
    SB_CARRY mod_5_add_1071_4 (.CI(n22296), .I0(n1508), .I1(n1532), .CO(n22297));
    SB_CARRY mod_5_add_1875_20 (.CI(n22543), .I0(n2692), .I1(n2720), .CO(n22544));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n22542), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_3 (.CI(n21905), .I0(bit_ctr[1]), .I1(GND_net), .CO(n21906));
    SB_CARRY mod_5_add_1875_19 (.CI(n22542), .I0(n2693), .I1(n2720), .CO(n22543));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n22541), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n22541), .I0(n2694), .I1(n2720), .CO(n22542));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n22540), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n22540), .I0(n2695), .I1(n2720), .CO(n22541));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n22539), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n22539), .I0(n2696), .I1(n2720), .CO(n22540));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n22538), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n30263), 
            .I3(n22295), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_15 (.CI(n22538), .I0(n2697), .I1(n2720), .CO(n22539));
    SB_CARRY mod_5_add_1071_3 (.CI(n22295), .I0(n1509), .I1(n30263), .CO(n22296));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n22537), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n22537), .I0(n2698), .I1(n2720), .CO(n22538));
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n30261), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_399[10]), .I1(timer[6]), 
            .I2(n56[6]), .I3(n22136), .O(n9_adj_4413)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n22536), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n14736), 
            .D(n255[23]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1875_13 (.CI(n22536), .I0(n2699), .I1(n2720), .CO(n22537));
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n14736), 
            .D(n255[22]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n22535), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n21910), .I0(bit_ctr[6]), .I1(GND_net), .CO(n21911));
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n14736), 
            .D(n255[21]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1875_12 (.CI(n22535), .I0(n2700), .I1(n2720), .CO(n22536));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n22534), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n22534), .I0(n2701), .I1(n2720), .CO(n22535));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n22533), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n22533), .I0(n2702), .I1(n2720), .CO(n22534));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n22532), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n22532), .I0(n2703), .I1(n2720), .CO(n22533));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n22531), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n22531), .I0(n2704), .I1(n2720), .CO(n22532));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n22530), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1588 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4447));
    defparam i10_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_7 (.CI(n22530), .I0(n2705), .I1(n2720), .CO(n22531));
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n14736), 
            .D(n255[20]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n22529), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n22529), .I0(n2706), .I1(n2720), .CO(n22530));
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n30261), 
            .CO(n22208));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n22528), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_8 (.CI(n22136), .I0(timer[6]), .I1(n56[6]), 
            .CO(n22137));
    SB_CARRY mod_5_add_1875_5 (.CI(n22528), .I0(n2707), .I1(n2720), .CO(n22529));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n30263), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n30263), 
            .CO(n22295));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n22527), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n22527), .I0(n2708), .I1(n2720), .CO(n22528));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n30265), 
            .I3(n22526), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n22526), .I0(n2709), .I1(n30265), .CO(n22527));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n56[5]), 
            .I3(n22135), .O(one_wire_N_399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_21 (.CI(n21923), .I0(bit_ctr[19]), .I1(GND_net), .CO(n21924));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n22294), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n30265), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n30265), 
            .CO(n22526));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n22525), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n21922), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n22524), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n22293), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n22524), .I0(n2589), .I1(n2621), .CO(n22525));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n22523), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n22523), .I0(n2590), .I1(n2621), .CO(n22524));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n22522), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n22522), .I0(n2591), .I1(n2621), .CO(n22523));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n22521), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n22521), .I0(n2592), .I1(n2621), .CO(n22522));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n22520), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n22520), .I0(n2593), .I1(n2621), .CO(n22521));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n22519), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n21922), .I0(bit_ctr[18]), .I1(GND_net), .CO(n21923));
    SB_CARRY mod_5_add_1808_18 (.CI(n22519), .I0(n2594), .I1(n2621), .CO(n22520));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n22518), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n22518), .I0(n2595), .I1(n2621), .CO(n22519));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n22517), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n22517), .I0(n2596), .I1(n2621), .CO(n22518));
    SB_CARRY sub_14_add_2_7 (.CI(n22135), .I0(timer[5]), .I1(n56[5]), 
            .CO(n22136));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n22516), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n56[4]), 
            .I3(n22134), .O(one_wire_N_399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n22134), .I0(timer[4]), .I1(n56[4]), 
            .CO(n22135));
    SB_CARRY mod_5_add_1138_13 (.CI(n22293), .I0(n1599), .I1(n1631), .CO(n22294));
    SB_CARRY mod_5_add_1808_15 (.CI(n22516), .I0(n2597), .I1(n2621), .CO(n22517));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n22515), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1589 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4448));
    defparam i16_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n22292), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n56[3]), 
            .I3(n22133), .O(one_wire_N_399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_14 (.CI(n22515), .I0(n2598), .I1(n2621), .CO(n22516));
    SB_CARRY sub_14_add_2_5 (.CI(n22133), .I0(timer[3]), .I1(n56[3]), 
            .CO(n22134));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n22514), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n56[2]), 
            .I3(n22132), .O(one_wire_N_399[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_13 (.CI(n22514), .I0(n2599), .I1(n2621), .CO(n22515));
    SB_LUT4 i14_4_lut_adj_1590 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4449));
    defparam i14_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n22513), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n22513), .I0(n2600), .I1(n2621), .CO(n22514));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n22512), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n21921), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n22512), .I0(n2601), .I1(n2621), .CO(n22513));
    SB_LUT4 i15_4_lut_adj_1591 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4450));
    defparam i15_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1592 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4451));
    defparam i13_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n22511), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_4 (.CI(n22132), .I0(timer[2]), .I1(n56[2]), 
            .CO(n22133));
    SB_CARRY mod_5_add_1808_10 (.CI(n22511), .I0(n2602), .I1(n2621), .CO(n22512));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n22510), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n22292), .I0(n1600), .I1(n1631), .CO(n22293));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_399[2]), .I1(timer[1]), .I2(n56[1]), 
            .I3(n22131), .O(n4_adj_4452)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_9 (.CI(n22510), .I0(n2603), .I1(n2621), .CO(n22511));
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4453));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n22509), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n22291), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n22131), .I0(timer[1]), .I1(n56[1]), 
            .CO(n22132));
    SB_LUT4 sub_14_add_2_2_lut (.I0(n4_adj_4452), .I1(timer[0]), .I2(n56[0]), 
            .I3(VCC_net), .O(n27201)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_8 (.CI(n22509), .I0(n2604), .I1(n2621), .CO(n22510));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n22508), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n22508), .I0(n2605), .I1(n2621), .CO(n22509));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n22507), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18_4_lut_adj_1593 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4454));
    defparam i18_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1594 (.I0(n37_adj_4451), .I1(n39_adj_4450), .I2(n38_adj_4449), 
            .I3(n40_adj_4448), .O(n46_adj_4455));
    defparam i22_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4456));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1595 (.I0(n33_adj_4456), .I1(n46_adj_4455), .I2(n42_adj_4454), 
            .I3(n34_adj_4453), .O(n2819));
    defparam i23_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i25172_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30262));
    defparam i25172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1596 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4457));
    defparam i8_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n14958));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1808_6 (.CI(n22507), .I0(n2606), .I1(n2621), .CO(n22508));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n22506), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n14736), 
            .D(n255[19]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1808_5 (.CI(n22506), .I0(n2607), .I1(n2621), .CO(n22507));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n22505), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n22505), .I0(n2608), .I1(n2621), .CO(n22506));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n56[0]), 
            .CO(n22131));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n30266), 
            .I3(n22504), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n22504), .I0(n2609), .I1(n30266), .CO(n22505));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n30266), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n30266), 
            .CO(n22504));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n22503), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n22502), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n22502), .I0(n2490), .I1(n2522), .CO(n22503));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n22501), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n22501), .I0(n2491), .I1(n2522), .CO(n22502));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n22500), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n22500), .I0(n2492), .I1(n2522), .CO(n22501));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n22499), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n15476));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1138_11 (.CI(n22291), .I0(n1601), .I1(n1631), .CO(n22292));
    SB_CARRY mod_5_add_1741_19 (.CI(n22499), .I0(n2493), .I1(n2522), .CO(n22500));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n22290), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n22498), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n22498), .I0(n2494), .I1(n2522), .CO(n22499));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n22497), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n22497), .I0(n2495), .I1(n2522), .CO(n22498));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n22496), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n22496), .I0(n2496), .I1(n2522), .CO(n22497));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n22495), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n22495), .I0(n2497), .I1(n2522), .CO(n22496));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n22494), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n22494), .I0(n2498), .I1(n2522), .CO(n22495));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n22493), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n22493), .I0(n2499), .I1(n2522), .CO(n22494));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n22492), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n22492), .I0(n2500), .I1(n2522), .CO(n22493));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n22491), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n22491), .I0(n2501), .I1(n2522), .CO(n22492));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n22490), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n22490), .I0(n2502), .I1(n2522), .CO(n22491));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n22489), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n22489), .I0(n2503), .I1(n2522), .CO(n22490));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n22488), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n22488), .I0(n2504), .I1(n2522), .CO(n22489));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n22487), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n22487), .I0(n2505), .I1(n2522), .CO(n22488));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n22486), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n22486), .I0(n2506), .I1(n2522), .CO(n22487));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n22485), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n22485), .I0(n2507), .I1(n2522), .CO(n22486));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n22484), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n22484), .I0(n2508), .I1(n2522), .CO(n22485));
    SB_LUT4 i9_4_lut_adj_1597 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4458));
    defparam i9_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1598 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4459));
    defparam i7_3_lut_adj_1598.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n30268), 
            .I3(n22483), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i13_4_lut_adj_1599 (.I0(n21_adj_4459), .I1(n23_adj_4458), .I2(n22_adj_4457), 
            .I3(n24_adj_4447), .O(n1829));
    defparam i13_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_3 (.CI(n22483), .I0(n2509), .I1(n30268), .CO(n22484));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n30268), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n30268), 
            .CO(n22483));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n22482), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n22481), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n22481), .I0(n2391), .I1(n2423), .CO(n22482));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n22480), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n22480), .I0(n2392), .I1(n2423), .CO(n22481));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n22479), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n22479), .I0(n2393), .I1(n2423), .CO(n22480));
    SB_CARRY add_21_19 (.CI(n21921), .I0(bit_ctr[17]), .I1(GND_net), .CO(n21922));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n22478), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n22478), .I0(n2394), .I1(n2423), .CO(n22479));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n22477), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n22477), .I0(n2395), .I1(n2423), .CO(n22478));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n22476), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n22476), .I0(n2396), .I1(n2423), .CO(n22477));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n22475), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n22475), .I0(n2397), .I1(n2423), .CO(n22476));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n22474), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n22474), .I0(n2398), .I1(n2423), .CO(n22475));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n22473), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n22473), .I0(n2399), .I1(n2423), .CO(n22474));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n22472), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n22472), .I0(n2400), .I1(n2423), .CO(n22473));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n22471), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n22471), .I0(n2401), .I1(n2423), .CO(n22472));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n22470), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n22470), .I0(n2402), .I1(n2423), .CO(n22471));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n22469), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n22469), .I0(n2403), .I1(n2423), .CO(n22470));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n22468), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n22468), .I0(n2404), .I1(n2423), .CO(n22469));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n22467), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n22467), .I0(n2405), .I1(n2423), .CO(n22468));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n22466), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n22466), .I0(n2406), .I1(n2423), .CO(n22467));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n22465), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n22465), .I0(n2407), .I1(n2423), .CO(n22466));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n22464), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n22464), .I0(n2408), .I1(n2423), .CO(n22465));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n30269), 
            .I3(n22463), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n22463), .I0(n2409), .I1(n30269), .CO(n22464));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n30269), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n30269), 
            .CO(n22463));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n22462), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n22461), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n22461), .I0(n906), .I1(VCC_net), .CO(n22462));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n26696), .I2(VCC_net), 
            .I3(n22460), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n22460), .I0(n26696), .I1(VCC_net), 
            .CO(n22461));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n14818), .I2(VCC_net), 
            .I3(n22459), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n22459), .I0(n14818), .I1(VCC_net), 
            .CO(n22460));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n12170), .I2(GND_net), 
            .I3(n22458), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n22458), .I0(n12170), .I1(GND_net), 
            .CO(n22459));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n22458));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4390), .I1(n4_adj_4390), .I2(n1037), 
            .I3(n22457), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n22456), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n22456), .I0(n1005), .I1(n1037), .CO(n22457));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n22455), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n22455), .I0(n1006), .I1(n1037), .CO(n22456));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n22454), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n22454), .I0(n1007), .I1(n1037), .CO(n22455));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n22453), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n22453), .I0(n1008), .I1(n1037), .CO(n22454));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n30270), 
            .I3(n22452), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n22452), .I0(n1009), .I1(n30270), .CO(n22453));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n30270), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n30270), 
            .CO(n22452));
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n15475));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n15474));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n15473));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n15472));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n15471));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1138_10 (.CI(n22290), .I0(n1602), .I1(n1631), .CO(n22291));
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n15470));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n15469));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n15468));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n18738), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n15467));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n18738), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n23680));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n15466));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n15465));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n15464));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n15463));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n15462));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n15461));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n15460));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n15459));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n15458));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n15457));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n15456));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n15455));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n15454));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n15453));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n15452));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n15451));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n22289), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n15450));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n15449));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n15448));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n15447));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n15446));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1138_9 (.CI(n22289), .I0(n1603), .I1(n1631), .CO(n22290));
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n24720));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n21909), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n22288), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n22288), .I0(n1604), .I1(n1631), .CO(n22289));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n22287), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n22013), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n21920), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_7 (.CI(n21909), .I0(bit_ctr[5]), .I1(GND_net), .CO(n21910));
    SB_CARRY mod_5_add_1138_7 (.CI(n22287), .I0(n1605), .I1(n1631), .CO(n22288));
    SB_CARRY add_21_18 (.CI(n21920), .I0(bit_ctr[16]), .I1(GND_net), .CO(n21921));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n22286), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n22286), .I0(n1606), .I1(n1631), .CO(n22287));
    SB_LUT4 i14913_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n18738));
    defparam i14913_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n22285), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21632_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n18738), .I2(n608), 
            .I3(bit_ctr[29]), .O(n26710));
    defparam i21632_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_CARRY mod_5_add_1138_5 (.CI(n22285), .I0(n1607), .I1(n1631), .CO(n22286));
    SB_LUT4 i24631_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n26798), .I2(bit_ctr[27]), 
            .I3(n838), .O(n14818));
    defparam i24631_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 i3324_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n26798), .I2(bit_ctr[27]), 
            .I3(n26662), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3324_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_LUT4 i25182_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30272));
    defparam i25182_1_lut.LUT_INIT = 16'h5555;
    SB_DFF timer_1126__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i24462_2_lut_4_lut (.I0(LED_c), .I1(bit_ctr[3]), .I2(bit_ctr[4]), 
            .I3(n11306), .O(n29274));   // verilog/neopixel.v(16[20:25])
    defparam i24462_2_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n20610), 
            .I3(\neo_pixel_transmitter.done ), .O(n28257));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n22284), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n21905));
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n21919), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n21908), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_4 (.CI(n22284), .I0(n1608), .I1(n1631), .CO(n22285));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n30267), 
            .I3(n22283), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n14736), 
            .D(n255[31]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n14736), 
            .D(n255[30]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n14736), 
            .D(n255[29]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n26842), .D(\neo_pixel_transmitter.done_N_462 ), 
            .R(n28257));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n22012), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_3 (.CI(n22283), .I0(n1609), .I1(n30267), .CO(n22284));
    SB_CARRY mod_5_add_1540_19 (.CI(n22012), .I0(n2193), .I1(n2225), .CO(n22013));
    SB_CARRY add_21_17 (.CI(n21919), .I0(bit_ctr[15]), .I1(GND_net), .CO(n21920));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n21918), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n14736), 
            .D(n255[28]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n22401), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n22400), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n22400), .I0(n1104), .I1(n1136), .CO(n22401));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n22399), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n22399), .I0(n1105), .I1(n1136), .CO(n22400));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n22398), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n22398), .I0(n1106), .I1(n1136), .CO(n22399));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n22397), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n22397), .I0(n1107), .I1(n1136), .CO(n22398));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n22396), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n30267), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i4_3_lut_adj_1600 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4460));
    defparam i4_3_lut_adj_1600.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1601 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4461));
    defparam i8_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n22011), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_3_lut_adj_1602 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4462));
    defparam i7_3_lut_adj_1602.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1603 (.I0(n21_adj_4461), .I1(n17_adj_4460), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4463));
    defparam i11_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1604 (.I0(n1700), .I1(n24_adj_4463), .I2(n20_adj_4462), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_4 (.CI(n22396), .I0(n1108), .I1(n1136), .CO(n22397));
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n30267), 
            .CO(n22283));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n30271), 
            .I3(n22395), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n22395), .I0(n1109), .I1(n30271), .CO(n22396));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n30271), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n30271), 
            .CO(n22395));
    SB_CARRY mod_5_add_1540_18 (.CI(n22011), .I0(n2194), .I1(n2225), .CO(n22012));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n22010), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25_4_lut_adj_1605 (.I0(n20572), .I1(n20573), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n11_adj_4464));   // verilog/neopixel.v(16[20:25])
    defparam i25_4_lut_adj_1605.LUT_INIT = 16'hcafa;
    SB_DFF timer_1126__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1126__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n11_adj_4464));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_16 (.CI(n21918), .I0(bit_ctr[14]), .I1(GND_net), .CO(n21919));
    SB_CARRY mod_5_add_1540_17 (.CI(n22010), .I0(n2195), .I1(n2225), .CO(n22011));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n21917), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n21917), .I0(bit_ctr[13]), .I1(GND_net), .CO(n21918));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n22282), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n22281), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n22281), .I0(n1698), .I1(n1730), .CO(n22282));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n22280), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n21916), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n22009), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n22280), .I0(n1699), .I1(n1730), .CO(n22281));
    SB_CARRY mod_5_add_1540_16 (.CI(n22009), .I0(n2196), .I1(n2225), .CO(n22010));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n22279), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n22279), .I0(n1700), .I1(n1730), .CO(n22280));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n22008), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n22278), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n22278), .I0(n1701), .I1(n1730), .CO(n22279));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n22277), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n21908), .I0(bit_ctr[4]), .I1(GND_net), .CO(n21909));
    SB_CARRY mod_5_add_1205_10 (.CI(n22277), .I0(n1702), .I1(n1730), .CO(n22278));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n22276), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n22008), .I0(n2197), .I1(n2225), .CO(n22009));
    SB_CARRY add_21_14 (.CI(n21916), .I0(bit_ctr[12]), .I1(GND_net), .CO(n21917));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n22007), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n22276), .I0(n1703), .I1(n1730), .CO(n22277));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n22275), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n22275), .I0(n1704), .I1(n1730), .CO(n22276));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n22274), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n22274), .I0(n1705), .I1(n1730), .CO(n22275));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n22273), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n22273), .I0(n1706), .I1(n1730), .CO(n22274));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n22272), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25181_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30271));
    defparam i25181_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_5 (.CI(n22272), .I0(n1707), .I1(n1730), .CO(n22273));
    SB_LUT4 i15187_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n19015));
    defparam i15187_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n22271), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n19015), .I3(n1108), 
            .O(n12_adj_4465));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_14 (.CI(n22007), .I0(n2198), .I1(n2225), .CO(n22008));
    SB_LUT4 i6_4_lut_adj_1606 (.I0(n1107), .I1(n12_adj_4465), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i24725_4_lut (.I0(n20565), .I1(n26806), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n29601));
    defparam i24725_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i24242_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n29332));
    defparam i24242_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53_4_lut (.I0(n26806), .I1(n20610), .I2(\state[1] ), .I3(start), 
            .O(n26838));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n26838), .I1(n26727), .I2(n29332), .I3(n29601), 
            .O(n26842));
    defparam i52_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i59_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_462 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i59_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_4 (.CI(n22271), .I0(n1708), .I1(n1730), .CO(n22272));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n30272), 
            .I3(n22270), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n22270), .I0(n1709), .I1(n30272), .CO(n22271));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n30272), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n30272), 
            .CO(n22270));
    SB_LUT4 timer_1126_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n22363), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1126_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n22362), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25177_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30267));
    defparam i25177_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1126_add_4_32 (.CI(n22362), .I0(GND_net), .I1(timer[30]), 
            .CO(n22363));
    SB_LUT4 timer_1126_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n22361), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_31 (.CI(n22361), .I0(GND_net), .I1(timer[29]), 
            .CO(n22362));
    SB_LUT4 timer_1126_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n22360), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_30 (.CI(n22360), .I0(GND_net), .I1(timer[28]), 
            .CO(n22361));
    SB_LUT4 timer_1126_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n22359), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_29 (.CI(n22359), .I0(GND_net), .I1(timer[27]), 
            .CO(n22360));
    SB_LUT4 timer_1126_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n22358), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_28 (.CI(n22358), .I0(GND_net), .I1(timer[26]), 
            .CO(n22359));
    SB_LUT4 timer_1126_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n22357), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_27 (.CI(n22357), .I0(GND_net), .I1(timer[25]), 
            .CO(n22358));
    SB_LUT4 timer_1126_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n22356), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_26 (.CI(n22356), .I0(GND_net), .I1(timer[24]), 
            .CO(n22357));
    SB_LUT4 timer_1126_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n22355), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_25 (.CI(n22355), .I0(GND_net), .I1(timer[23]), 
            .CO(n22356));
    SB_LUT4 timer_1126_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n22354), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_24 (.CI(n22354), .I0(GND_net), .I1(timer[22]), 
            .CO(n22355));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n22269), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n14736), 
            .D(n255[27]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n22268), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1126_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n22353), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_23 (.CI(n22353), .I0(GND_net), .I1(timer[21]), 
            .CO(n22354));
    SB_LUT4 timer_1126_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n22352), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n22006), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n14736), 
            .D(n255[26]), .R(n14862));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1272_15 (.CI(n22268), .I0(n1797), .I1(n1829), .CO(n22269));
    SB_CARRY timer_1126_add_4_22 (.CI(n22352), .I0(GND_net), .I1(timer[20]), 
            .CO(n22353));
    SB_LUT4 timer_1126_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n22351), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_21 (.CI(n22351), .I0(GND_net), .I1(timer[19]), 
            .CO(n22352));
    SB_LUT4 timer_1126_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n22350), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_20 (.CI(n22350), .I0(GND_net), .I1(timer[18]), 
            .CO(n22351));
    SB_LUT4 timer_1126_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n22349), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_19 (.CI(n22349), .I0(GND_net), .I1(timer[17]), 
            .CO(n22350));
    SB_LUT4 timer_1126_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n22348), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_18 (.CI(n22348), .I0(GND_net), .I1(timer[16]), 
            .CO(n22349));
    SB_LUT4 timer_1126_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n22347), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_17 (.CI(n22347), .I0(GND_net), .I1(timer[15]), 
            .CO(n22348));
    SB_LUT4 timer_1126_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n22346), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1126_add_4_16 (.CI(n22346), .I0(GND_net), .I1(timer[14]), 
            .CO(n22347));
    SB_LUT4 timer_1126_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n22345), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1126_add_4_15_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, clk32MHz, 
            data_o, n27693, reg_B, ENCODER1_A_c_1, ENCODER1_B_c_0, 
            VCC_net, n15442, n14956) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n27693;
    output [1:0]reg_B;
    input ENCODER1_A_c_1;
    input ENCODER1_B_c_0;
    input VCC_net;
    input n15442;
    input n14956;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2424;
    
    wire n2400, n22114, n22115, n22113, n22112, n22111, n22110, 
        count_enable, B_delayed, A_delayed, n22109, n22108, count_direction, 
        n22107, n22130, n22129, n22128, n22127, n22126, n22125, 
        n22124, n22123, n22122, n22121, n22120, n22119, n22118, 
        n22117, n22116;
    
    SB_LUT4 add_528_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2400), 
            .I3(n22114), .O(n2424[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_9 (.CI(n22114), .I0(encoder1_position[7]), .I1(n2400), 
            .CO(n22115));
    SB_LUT4 add_528_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2400), 
            .I3(n22113), .O(n2424[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_8 (.CI(n22113), .I0(encoder1_position[6]), .I1(n2400), 
            .CO(n22114));
    SB_LUT4 add_528_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2400), 
            .I3(n22112), .O(n2424[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_7 (.CI(n22112), .I0(encoder1_position[5]), .I1(n2400), 
            .CO(n22113));
    SB_LUT4 add_528_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2400), 
            .I3(n22111), .O(n2424[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_6 (.CI(n22111), .I0(encoder1_position[4]), .I1(n2400), 
            .CO(n22112));
    SB_LUT4 add_528_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2400), 
            .I3(n22110), .O(n2424[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_528_5 (.CI(n22110), .I0(encoder1_position[3]), .I1(n2400), 
            .CO(n22111));
    SB_LUT4 add_528_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2400), 
            .I3(n22109), .O(n2424[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_4 (.CI(n22109), .I0(encoder1_position[2]), .I1(n2400), 
            .CO(n22110));
    SB_LUT4 add_528_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2400), 
            .I3(n22108), .O(n2424[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_3 (.CI(n22108), .I0(encoder1_position[1]), .I1(n2400), 
            .CO(n22109));
    SB_LUT4 add_528_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n22107), .O(n2424[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_2 (.CI(n22107), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n22108));
    SB_CARRY add_528_1 (.CI(GND_net), .I0(n2400), .I1(n2400), .CO(n22107));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[1]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2424[23]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_528_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2400), 
            .I3(n22130), .O(n2424[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_528_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2400), 
            .I3(n22129), .O(n2424[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_24 (.CI(n22129), .I0(encoder1_position[22]), .I1(n2400), 
            .CO(n22130));
    SB_LUT4 add_528_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2400), 
            .I3(n22128), .O(n2424[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_23 (.CI(n22128), .I0(encoder1_position[21]), .I1(n2400), 
            .CO(n22129));
    SB_LUT4 add_528_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2400), 
            .I3(n22127), .O(n2424[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_22 (.CI(n22127), .I0(encoder1_position[20]), .I1(n2400), 
            .CO(n22128));
    SB_LUT4 add_528_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2400), 
            .I3(n22126), .O(n2424[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_21 (.CI(n22126), .I0(encoder1_position[19]), .I1(n2400), 
            .CO(n22127));
    SB_LUT4 add_528_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2400), 
            .I3(n22125), .O(n2424[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_20 (.CI(n22125), .I0(encoder1_position[18]), .I1(n2400), 
            .CO(n22126));
    SB_LUT4 i863_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2400));   // quad.v(37[5] 40[8])
    defparam i863_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_528_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2400), 
            .I3(n22124), .O(n2424[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_19 (.CI(n22124), .I0(encoder1_position[17]), .I1(n2400), 
            .CO(n22125));
    SB_LUT4 add_528_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2400), 
            .I3(n22123), .O(n2424[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_18 (.CI(n22123), .I0(encoder1_position[16]), .I1(n2400), 
            .CO(n22124));
    SB_LUT4 add_528_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2400), 
            .I3(n22122), .O(n2424[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_17 (.CI(n22122), .I0(encoder1_position[15]), .I1(n2400), 
            .CO(n22123));
    SB_LUT4 add_528_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2400), 
            .I3(n22121), .O(n2424[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_16 (.CI(n22121), .I0(encoder1_position[14]), .I1(n2400), 
            .CO(n22122));
    SB_LUT4 add_528_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2400), 
            .I3(n22120), .O(n2424[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_15 (.CI(n22120), .I0(encoder1_position[13]), .I1(n2400), 
            .CO(n22121));
    SB_LUT4 add_528_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2400), 
            .I3(n22119), .O(n2424[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_14 (.CI(n22119), .I0(encoder1_position[12]), .I1(n2400), 
            .CO(n22120));
    SB_LUT4 add_528_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2400), 
            .I3(n22118), .O(n2424[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_13 (.CI(n22118), .I0(encoder1_position[11]), .I1(n2400), 
            .CO(n22119));
    SB_LUT4 add_528_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2400), 
            .I3(n22117), .O(n2424[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_12 (.CI(n22117), .I0(encoder1_position[10]), .I1(n2400), 
            .CO(n22118));
    SB_LUT4 add_528_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2400), 
            .I3(n22116), .O(n2424[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_11 (.CI(n22116), .I0(encoder1_position[9]), .I1(n2400), 
            .CO(n22117));
    SB_LUT4 add_528_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2400), 
            .I3(n22115), .O(n2424[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_528_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_528_10 (.CI(n22115), .I0(encoder1_position[8]), .I1(n2400), 
            .CO(n22116));
    \grp_debouncer(2,100)  debounce (.n27693(n27693), .reg_B({reg_B}), .GND_net(GND_net), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .VCC_net(VCC_net), .n15442(n15442), .data_o({data_o}), .n14956(n14956));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (n27693, reg_B, GND_net, ENCODER1_A_c_1, 
            clk32MHz, ENCODER1_B_c_0, VCC_net, n15442, data_o, n14956);
    output n27693;
    output [1:0]reg_B;
    input GND_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input ENCODER1_B_c_0;
    input VCC_net;
    input n15442;
    output [1:0]data_o;
    input n14956;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3576;
    wire [6:0]n33;
    
    wire n22451, n22450, n22449, n22448, n22447, n22446;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[3]), .I2(cnt_reg[6]), 
            .I3(cnt_reg[5]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(n12), .I2(cnt_reg[2]), .I3(cnt_reg[4]), 
            .O(n27693));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n27693), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1134__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1134_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n22451), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1134_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n22450), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_7 (.CI(n22450), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n22451));
    SB_LUT4 cnt_reg_1134_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n22449), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_6 (.CI(n22449), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n22450));
    SB_LUT4 cnt_reg_1134_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n22448), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_5 (.CI(n22448), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n22449));
    SB_LUT4 cnt_reg_1134_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n22447), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_4 (.CI(n22447), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n22448));
    SB_LUT4 cnt_reg_1134_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n22446), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_3 (.CI(n22446), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n22447));
    SB_LUT4 cnt_reg_1134_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1134_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1134_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n22446));
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n15442));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n14956));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1134__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1134__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1134__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1134__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1134__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1134__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3576));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[1] , GND_net, \Ki[8] , \Ki[0] , \Ki[2] , 
            PWMLimit, \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , 
            \Ki[9] , \Ki[10] , \Kp[5] , \Kp[1] , IntegralLimit, duty, 
            \Kp[9] , \Kp[6] , \Kp[4] , \Kp[3] , \Kp[2] , \Kp[0] , 
            \Kp[10] , \Kp[8] , \Kp[7] , \Kp[11] , \Kp[12] , \Kp[13] , 
            \Kp[14] , \Kp[15] , \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , 
            \Ki[15] , clk32MHz, n30253, VCC_net, setpoint, motor_state, 
            n25) /* synthesis syn_module_defined=1 */ ;
    input \Ki[1] ;
    input GND_net;
    input \Ki[8] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input [23:0]PWMLimit;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Kp[5] ;
    input \Kp[1] ;
    input [23:0]IntegralLimit;
    output [23:0]duty;
    input \Kp[9] ;
    input \Kp[6] ;
    input \Kp[4] ;
    input \Kp[3] ;
    input \Kp[2] ;
    input \Kp[0] ;
    input \Kp[10] ;
    input \Kp[8] ;
    input \Kp[7] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input clk32MHz;
    output n30253;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input n25;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n110, n606;
    wire [11:0]n6776;
    wire [10:0]n6790;
    
    wire n545, n22843, n41, n22844, n472, n22842, n183;
    wire [47:0]n155;
    
    wire n256;
    wire [23:0]n2554;
    
    wire n256_adj_3903, n39;
    wire [23:0]n1;
    
    wire n22180, n399, n22841, n329, n326, n22840, n22181, n402, 
        n253, n22839, n475, n548, n621, n694, n767;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(21[23:26])
    
    wire n13, n17, n9, n11, n29500, n29498, n31055, n29899, 
        n29766, n31037, n29764, n29762, n31031, n27, n15, n13_adj_3904, 
        n11_adj_3905, n29428, n21, n19, n17_adj_3906, n9_adj_3907, 
        n29434, n43, n16, n29407, n8, n45, n24, n7, n5, n29444, 
        n180, n22838, n29738, n29734, n25_c, n23, n30042, n31, 
        n29, n29877, n37, n35, n33, n30072, n29768, n38, n107, 
        n31024, n29756, n31019, n12, n29478, n31042, n10, n30, 
        n22179, n29971, n29486, n31022, n29893, n31048;
    wire [12:0]n6761;
    
    wire n980, n22837, n30046, n31013, n30103, n907, n22836, n31010, 
        n16_adj_3909, n22178, n834, n22835, n29446, n761, n22834, 
        n688, n22833, n615, n22832, n24_adj_3911, n6_adj_3912, n29929, 
        n29930, n29448, n542, n22831, n8_adj_3913, n31008, n29869, 
        n29712;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3467 ;
    
    wire n3, n4, n30012, n469, n22830, n30013, n12_adj_3914, n29417, 
        n10_adj_3915, n30_adj_3916, n29420, n30081, n29948, n30127, 
        n30128, n30112, n6_adj_3917, n29921, n29922, n29409, n29871, 
        n29722, n41_adj_3918, n29411, n30026, n40, n30028, n4_adj_3919, 
        n29927, n29928, n29480, n30066, n29714, n396, n22829;
    wire [5:0]n7142;
    
    wire n27773, n490, n23136;
    wire [4:0]n7150;
    
    wire n417, n23135, n344, n23134, n271, n23133, n198, n23132, 
        n56, n125;
    wire [6:0]n7133;
    
    wire n560, n23131, n487, n23130, n414, n23129, n341, n23128, 
        n268, n23127, n195, n23126, n53, n122;
    wire [7:0]n7123;
    
    wire n630, n23125, n557, n23124, n30115, n484, n23123, n411, 
        n23122, n338, n23121, n265, n23120, n192, n23119, n50, 
        n119;
    wire [8:0]n7112;
    
    wire n700, n23118, n627, n23117, n554, n23116, n481, n23115, 
        n408, n23114, n335, n23113, n262, n23112, n189, n23111, 
        n47, n116;
    wire [9:0]n7100;
    
    wire n770, n23110, n697, n23109, n624, n23108, n551, n23107, 
        n478, n23106, n405, n23105, n332, n23104, n259, n23103, 
        n186, n23102, n44, n113;
    wire [10:0]n7087;
    
    wire n840, n23101, n23100, n23099, n23098, n23097, n23096, 
        n23095, n23094, n23093, n23092;
    wire [11:0]n7073;
    
    wire n910, n23091, n837, n23090, n764, n23089, n691, n23088, 
        n618, n23087, n30116, n545_adj_3920, n23086, n472_adj_3921, 
        n23085, n399_adj_3922, n23084, n326_adj_3923, n23083, n253_adj_3924, 
        n23082, n180_adj_3925, n23081, n38_adj_3926, n107_adj_3927;
    wire [12:0]n7058;
    
    wire n980_adj_3928, n23080, n907_adj_3929, n23079, n834_adj_3930, 
        n23078, n761_adj_3931, n23077, n688_adj_3932, n23076, n615_adj_3933, 
        n23075, n30090, n542_adj_3934, n23074, n469_adj_3935, n23073, 
        n396_adj_3936, n23072, n323, n23071, n250, n23070, n177, 
        n23069, n35_adj_3937, n104;
    wire [13:0]n7042;
    
    wire n1050, n23068, n977, n23067, n904, n23066, n831, n23065, 
        n758, n23064, n685, n23063, n612, n23062, n539, n23061, 
        n29472, n466, n23060, n393, n23059, n320, n23058, n247, 
        n23057, n174, n23056, n32, n101;
    wire [14:0]n7025;
    
    wire n1120, n23055, n1047, n23054, n974, n23053, n901, n23052, 
        n828, n23051, n755, n23050, n682, n23049, n609, n23048, 
        n536, n23047, n463, n23046, n390, n23045, n317, n23044, 
        n244, n23043, n171, n23042, n29_adj_3938, n98;
    wire [15:0]n7007;
    
    wire n23041, n1117, n23040, n1044, n23039, n971, n23038, n898, 
        n23037, n825, n23036, n752, n23035, n679, n23034, n23033, 
        n533, n23032, n460, n23031, n387, n23030, n314, n23029, 
        n241, n23028, n168, n23027, n26, n95;
    wire [16:0]n6988;
    
    wire n23026, n23025, n323_adj_3939, n22828, n1114, n23024, n1041, 
        n23023, n968, n23022, n895, n23021, n822, n23020, n749, 
        n23019, n676, n23018, n603, n23017, n530, n23016, n30022, 
        n29720, \PID_CONTROLLER.integral_23__N_3466 , n457, n23015, 
        n384, n23014, n311, n23013, n238, n23012, n165, n23011, 
        n23_adj_3940, n92;
    wire [17:0]n6968;
    
    wire n23010, n23009, n23008, n1111, n23007, n1038, n23006, 
        n965, n23005, n892, n23004, n819, n23003, n30074, n746, 
        n23002, \PID_CONTROLLER.integral_23__N_3464 , n250_adj_3941, n22827, 
        n177_adj_3942, n22826, n35_adj_3943, n104_adj_3944;
    wire [13:0]n6745;
    
    wire n1050_adj_3945, n22825, n673, n23001, n977_adj_3946, n22824, 
        n600, n23000, n904_adj_3947, n22823, n831_adj_3948, n22822, 
        n527, n22999, n758_adj_3949, n22821, n685_adj_3950, n22820, 
        n612_adj_3951, n22819, n539_adj_3952, n22818, n454, n22998, 
        n466_adj_3953, n22817, n393_adj_3954, n22816, n320_adj_3955, 
        n22815, n381, n22997, n247_adj_3956, n22814, n174_adj_3958, 
        n22813, n32_adj_3959, n101_adj_3960;
    wire [14:0]n6728;
    
    wire n1120_adj_3961, n22812, n308, n22996, n1047_adj_3962, n22811, 
        n974_adj_3963, n22810;
    wire [23:0]n257;
    
    wire n29370, n700_adj_3964, n481_adj_3965, n408_adj_3966, n335_adj_3967, 
        n262_adj_3968, n189_adj_3969, n116_adj_3970, n47_adj_3971, n770_adj_3972, 
        n901_adj_3973, n22809, n697_adj_3974, n22177, n624_adj_3976, 
        n29296, n828_adj_3977, n22808, n551_adj_3978, n478_adj_3979, 
        n405_adj_3980, n332_adj_3981, n259_adj_3982, n186_adj_3983, 
        n113_adj_3984, n235, n22995, n44_adj_3985, n840_adj_3986, 
        n767_adj_3987, n694_adj_3988, n621_adj_3989, n548_adj_3990, 
        n475_adj_3991, n402_adj_3992, n755_adj_3993, n22807, n329_adj_3994, 
        n256_adj_3995, n183_adj_3996, n110_adj_3997, n41_adj_3998, n910_adj_3999, 
        n837_adj_4000, n764_adj_4001, n691_adj_4002, n682_adj_4003, 
        n22806, n77, n8_adj_4004, n150, n223, n609_adj_4005, n22805, 
        n296, n369, n442, n515, n588, n661, n734, n807, n880, 
        n953, n1026, n1099, n74, n5_adj_4006, n147, n220, n536_adj_4007, 
        n22804, n293, n366, n439, n512, n585, n658, n731, n804, 
        n877, n950, n1023, n1096, n618_adj_4008, n463_adj_4009, 
        n22803, n119_adj_4010, n50_adj_4011, n192_adj_4012, n265_adj_4013, 
        n338_adj_4014, n41_adj_4015, n39_adj_4017, n162, n22994, n45_adj_4019, 
        n43_adj_4020, n37_adj_4021, n23_adj_4022, n25_adj_4023, n29_adj_4024, 
        n390_adj_4025, n22802, n31_adj_4026, n35_adj_4027, n11_adj_4028, 
        n13_adj_4029, n20, n89, n15_adj_4030, n27_adj_4032, n9_adj_4033, 
        n17_adj_4034, n19_adj_4035, n21_adj_4037, n33_adj_4039, n29360, 
        n29354, n12_adj_4040, n10_adj_4041, n30_adj_4042, n29646, 
        n29642, n30000, n29835, n30068, n16_adj_4043, n6_adj_4044, 
        n29986, n29987, n8_adj_4045, n24_adj_4046, n29340, n29338, 
        n29875, n29958, n29248, n4_adj_4047, n29984, n29985, n29350, 
        n29348, n30085, n29960, n30131, n30132, n30108, n29342;
    wire [18:0]n6947;
    
    wire n22993, n30038, n22992, n22991, n40_adj_4048, n22990, n1108, 
        n22989, n1035, n22988, n962, n22987, n30040, n47_adj_4049, 
        n889, n22986, n18679, n816, n22985, n411_adj_4050, n743, 
        n22984, n670, n22983, n317_adj_4051, n22801, n597, n22982, 
        n244_adj_4052, n22800, n524, n22981, n451, n22980, n171_adj_4053, 
        n22799, n484_adj_4054, n557_adj_4055, n378, n22979, n305, 
        n22978, n232, n22977, n29_adj_4056, n98_adj_4057, n630_adj_4058, 
        n159, n22976, n122_adj_4059;
    wire [15:0]n6710;
    
    wire n22798, n53_adj_4060, n80, n11_adj_4061, n195_adj_4062, n17_adj_4063, 
        n86, n268_adj_4064, n341_adj_4065, n414_adj_4066, n153, n1117_adj_4068, 
        n22797, n1044_adj_4069, n22796, n487_adj_4070, n560_adj_4071, 
        n125_adj_4072, n971_adj_4073, n22795, n56_adj_4074, n198_adj_4075, 
        n271_adj_4076, n898_adj_4077, n22794, n226, n344_adj_4078, 
        n417_adj_4079, n6_adj_4080;
    wire [3:0]n6860;
    wire [4:0]n6853;
    
    wire n299, n372, n825_adj_4082, n22793, n204, n22176;
    wire [1:0]n6871;
    
    wire n752_adj_4084, n22792, n131, n62, n4_adj_4085;
    wire [2:0]n6866;
    
    wire n490_adj_4086, n12_adj_4087, n8_adj_4088, n11_adj_4089, n6_adj_4090, 
        n21745, n18, n4_adj_4091, n27329, n77_adj_4092;
    wire [19:0]n6925;
    
    wire n22975, n8_adj_4093, n150_adj_4094, n445, n223_adj_4095, 
        n296_adj_4096, n369_adj_4097, n518, n442_adj_4098, n591, n22974, 
        n679_adj_4099, n22791, n606_adj_4100, n22790, n664, n737, 
        n22973, n22972, n810, n515_adj_4102, n883, n588_adj_4103, 
        n22971, n1105, n22970, n533_adj_4104, n22789, n22175, n460_adj_4106, 
        n22788, n387_adj_4107, n22787;
    wire [23:0]duty_23__N_3368;
    wire [23:0]\PID_CONTROLLER.err_23__N_3392 ;
    
    wire n314_adj_4108, n22786, n1032, n22969, n241_adj_4109, n22785, 
        n168_adj_4110, n22784, n959, n22968, n26_adj_4111, n95_adj_4112;
    wire [16:0]n6691;
    
    wire n22783, n886, n22967, n22782, n813, n22966, n740, n22965, 
        n1114_adj_4113, n22781, n667, n22964, n594, n22963, n521, 
        n22962, n1041_adj_4114, n22780, n448, n22961, n375, n22960, 
        n302, n22959, n968_adj_4115, n22779, n229, n22958, n156, 
        n22957, n22174, n14, n83;
    wire [20:0]n6902;
    
    wire n22956, n22955, n22954, n895_adj_4118, n22778, n22953, 
        n22173, n956, n822_adj_4120, n22777, n22952, n22951, n1102, 
        n22950, n1029, n22949, n22172, n661_adj_4122, n749_adj_4123, 
        n22776, n734_adj_4124, n22171, n807_adj_4126, n880_adj_4127, 
        n956_adj_4128, n22948, n676_adj_4129, n22775, n953_adj_4130, 
        n603_adj_4131, n22774, n530_adj_4132, n22773, n457_adj_4133, 
        n22772, n384_adj_4134, n22771, n1026_adj_4135, n22170, n311_adj_4137, 
        n22770, n238_adj_4138, n22769, n1099_adj_4139, n1029_adj_4140, 
        n165_adj_4141, n22768, n23_adj_4142, n92_adj_4143, n74_adj_4144;
    wire [17:0]n6671;
    
    wire n22767, n22766, n22765, n883_adj_4145, n22947, n1111_adj_4146, 
        n22764, n5_adj_4147, n147_adj_4148, n1102_adj_4149, n220_adj_4150, 
        n83_adj_4151, n14_adj_4152, n156_adj_4153, n293_adj_4154, n229_adj_4155, 
        n366_adj_4156, n439_adj_4157, n512_adj_4158, n302_adj_4159, 
        n585_adj_4160, n375_adj_4161, n810_adj_4162, n22946, n658_adj_4163, 
        n737_adj_4164, n22945, n664_adj_4165, n22944, n731_adj_4166, 
        n448_adj_4167, n591_adj_4168, n22943, n518_adj_4169, n22942, 
        n521_adj_4170, n445_adj_4171, n22941, n372_adj_4172, n22940, 
        n1038_adj_4173, n22763, n804_adj_4174, n594_adj_4175, n965_adj_4176, 
        n22762, n299_adj_4177, n22939, n667_adj_4179, n740_adj_4180, 
        n892_adj_4181, n22761, n819_adj_4182, n22760, n746_adj_4183, 
        n22759, n813_adj_4184, n226_adj_4185, n22938, n153_adj_4186, 
        n22937, n877_adj_4187, n22169, n673_adj_4189, n22758, n11_adj_4190, 
        n80_adj_4191, n886_adj_4192, n22168;
    wire [21:0]n6878;
    
    wire n22936, n959_adj_4194, n950_adj_4195, n22935, n22934, n1032_adj_4196, 
        n600_adj_4197, n22757, n527_adj_4198, n22756, n1023_adj_4199, 
        n454_adj_4200, n22755, n1105_adj_4201, n22167, n1096_adj_4203, 
        n86_adj_4205, n17_adj_4206, n159_adj_4207, n232_adj_4208, n381_adj_4209, 
        n22754, n305_adj_4210, n22933, n308_adj_4211, n22753, n22932, 
        n235_adj_4212, n22752, n162_adj_4213, n22751, n20_adj_4214, 
        n89_adj_4215, n378_adj_4216;
    wire [18:0]n6650;
    
    wire n22750, n451_adj_4217, n22749, n524_adj_4218, n597_adj_4219, 
        n22748, n670_adj_4220, n743_adj_4221, n816_adj_4222, n889_adj_4223, 
        n22931, n962_adj_4224, n1035_adj_4225, n1108_adj_4226, n22747, 
        n22746, n22745, n22744, n22743, n22742, n22741, n22740, 
        n22739, n22738, n22737, n22736, n22735, n22734, n22733, 
        n22930, n22929;
    wire [19:0]n6628;
    
    wire n22732, n22731, n22166, n22730, n22729, n22928, n22728, 
        n22727, n22927, n22726, n22926, n22725, n6_adj_4228;
    wire [3:0]n7157;
    
    wire n22724, n204_adj_4229, n22925, n22723, n22722;
    wire [1:0]n7168;
    
    wire n22721, n22165, n22720, n22924, n22719, n22718, n22923, 
        n22922, n22717, n22921, n22716, n22920, n22919, n22918, 
        n131_adj_4233, n62_adj_4234, n22715, n22917, n22714, n22164, 
        n4_adj_4235;
    wire [2:0]n7163;
    wire [20:0]n6605;
    
    wire n22713, n22712, n22711, n22710, n22709, n22708, n22916, 
        n22707, n22915, n22914, n22913, n22912, n22911, n22910, 
        n22909, n22706, n22908, n22907, n22906, n22905, n22904, 
        n22903, n22902, n22901, n22705, n22900, n22704, n22899, 
        n22703, n22702, n22163, n22701, n22700, n22898, n22699, 
        n22897, n22896, n22895, n22698, n22894;
    wire [5:0]n6845;
    
    wire n22893, n22697, n22696, n22162, n22892, n22891, n22695, 
        n22890, n22889;
    wire [6:0]n6836;
    
    wire n22888, n22887, n22694, n22886, n22885, n22884, n22883;
    wire [7:0]n6826;
    
    wire n22882, n22881, n22880, n22879;
    wire [0:0]n5022;
    wire [21:0]n6581;
    
    wire n22693, n12_adj_4236, n8_adj_4237, n11_adj_4238, n6_adj_4239, 
        n21877, n18_adj_4240, n13_adj_4241, n4_adj_4242;
    wire [23:0]n2529;
    
    wire n22692, n22878, n22691, n22877, n22876, n22690, n22845, 
        n22689, n22688, n22687, n22686, n22685, n22684, n22683, 
        n22682, n22681, n22680, n22679, n22678;
    wire [23:0]n1_adj_4311;
    
    wire n22677, n22676, n22675, n22674, n22673, n22672, n22671, 
        n22670, n22669, n22668, n22667, n22666, n22665, n22664, 
        n22663, n22662, n22661, n22660, n22659, n22658, n22657, 
        n22656, n22655, n22654, n22653, n22652, n22651, n41_adj_4244, 
        n39_adj_4245, n45_adj_4246, n37_adj_4247, n29_adj_4248, n31_adj_4249, 
        n43_adj_4250, n23_adj_4251, n25_adj_4252, n35_adj_4253, n33_adj_4254, 
        n11_adj_4255, n13_adj_4256, n15_adj_4257, n27_adj_4258, n9_adj_4259, 
        n17_adj_4260, n19_adj_4261, n21_adj_4262, n29395, n29389, 
        n12_adj_4263, n30_adj_4264, n29405, n29680, n29676, n30010, 
        n29851, n30070, n6_adj_4265, n29992, n29993, n16_adj_4266, 
        n24_adj_4267, n29374, n22846, n22847, n22848, n22849;
    wire [9:0]n6803;
    
    wire n22850, n22851, n8_adj_4268, n29372, n29873, n29952, n4_adj_4269, 
        n29990, n29991, n29385, n10_adj_4270, n29383, n30083, n29954, 
        n22852, n22853, n22854, n30129, n22855, n22856, n22857, 
        n22858, n30130, n30110, n29376, n30032, n40_adj_4271, n30034, 
        duty_23__N_3515;
    wire [23:0]duty_23__N_3491;
    
    wire n22859;
    wire [8:0]n6815;
    
    wire n22860, n22861, n22862, n22863, n22864, n22865, n22036, 
        n22035, n22034, n22866, n22867, n22868, n22869, n22870, 
        n22871, n22872, n22873, n22875, n22033;
    wire [23:0]n28;
    
    wire n22032, n22083, n22031, n554_adj_4277, n22030, n627_adj_4278, 
        n22082, n22029, n22081, n22080, n22028, n22079, n22078, 
        n22027, n22026, n4_adj_4282, n22077, n22025, n21775, n22076, 
        n22024, n22075, n21852, n22023, n22022, n22074, n22073, 
        n22021, n22072, n22020, n22071, n22070, n22019, n22069, 
        n22018, n22207, n22206, n22068, n22017, n22205, n22067, 
        n22016, n22204, n22066, n22874, n22015, n22203, n22202, 
        n22014, n22065, n22064, n22063, n22201, n22200, n22062, 
        n22199, n22424, n22423, n22422, n22421, n22420, n22419, 
        n22418, n22417, n22416, n22415, n22414, n22413, n22412, 
        n22061, n22411, n22410, n22409, n22198, n22408, n22407, 
        n22406, n22405, n22197, n22404, n22403, n22402, n22196, 
        n4_adj_4309, n22195, n22194, n21643, n22193, n22192, n22191, 
        n22190, n22189, n22188, n22187, n22186, n21720, n22185, 
        n22184, n22183, n22182;
    
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3394_8_lut (.I0(GND_net), .I1(n6790[5]), .I2(n545), .I3(n22843), 
            .O(n6776[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3394_8 (.CI(n22843), .I0(n6790[5]), .I1(n545), .CO(n22844));
    SB_LUT4 add_3394_7_lut (.I0(GND_net), .I1(n6790[4]), .I2(n472), .I3(n22842), 
            .O(n6776[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i19_3_lut (.I0(n155[18]), .I1(PWMLimit[18]), .I2(n256), 
            .I3(GND_net), .O(n2554[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i19_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3903));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3394_7 (.CI(n22842), .I0(n6790[4]), .I1(n472), .CO(n22843));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n22180), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3394_6_lut (.I0(GND_net), .I1(n6790[3]), .I2(n399), .I3(n22841), 
            .O(n6776[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3394_6 (.CI(n22841), .I0(n6790[3]), .I1(n399), .CO(n22842));
    SB_LUT4 add_3394_5_lut (.I0(GND_net), .I1(n6790[2]), .I2(n326), .I3(n22840), 
            .O(n6776[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n22180), .I0(GND_net), .I1(n1[19]), 
            .CO(n22181));
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3394_5 (.CI(n22840), .I0(n6790[2]), .I1(n326), .CO(n22841));
    SB_LUT4 add_3394_4_lut (.I0(GND_net), .I1(n6790[1]), .I2(n253), .I3(n22839), 
            .O(n6776[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13));   // verilog/motorControl.v(34[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3394_4 (.CI(n22839), .I0(n6790[1]), .I1(n253), .CO(n22840));
    SB_LUT4 mux_561_i20_3_lut (.I0(n155[19]), .I1(PWMLimit[19]), .I2(n256), 
            .I3(GND_net), .O(n2554[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24410_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n29500));
    defparam i24410_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i24408_3_lut (.I0(n11), .I1(n9), .I2(n29500), .I3(GND_net), 
            .O(n29498));
    defparam i24408_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_115_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n31055));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_115_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24807_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n31055), 
            .I2(IntegralLimit[7]), .I3(n29498), .O(n29899));
    defparam i24807_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i24674_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n29899), .O(n29766));
    defparam i24674_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_97_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n31037));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_97_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24672_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n9), .O(n29764));
    defparam i24672_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i24670_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n31037), 
            .I2(IntegralLimit[11]), .I3(n29764), .O(n29762));
    defparam i24670_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_91_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n31031));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_91_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24338_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_3904), .I3(n11_adj_3905), 
            .O(n29428));
    defparam i24338_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24344_4_lut (.I0(n21), .I1(n19), .I2(n17_adj_3906), .I3(n9_adj_3907), 
            .O(n29434));
    defparam i24344_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24317_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n29407));
    defparam i24317_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3906), .I3(GND_net), 
            .O(n8));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n45), .I3(GND_net), .O(n24));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24354_2_lut (.I0(n7), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n29444));
    defparam i24354_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_3394_3_lut (.I0(GND_net), .I1(n6790[0]), .I2(n180), .I3(n22838), 
            .O(n6776[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24646_4_lut (.I0(n13_adj_3904), .I1(n11_adj_3905), .I2(n9_adj_3907), 
            .I3(n29444), .O(n29738));
    defparam i24646_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24642_4_lut (.I0(n19), .I1(n17_adj_3906), .I2(n15), .I3(n29738), 
            .O(n29734));
    defparam i24642_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24950_4_lut (.I0(n25_c), .I1(n23), .I2(n21), .I3(n29734), 
            .O(n30042));
    defparam i24950_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24785_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n30042), 
            .O(n29877));
    defparam i24785_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24980_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n29877), 
            .O(n30072));
    defparam i24980_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24676_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n31055), 
            .I2(IntegralLimit[7]), .I3(n11), .O(n29768));
    defparam i24676_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_3394_3 (.CI(n22838), .I0(n6790[0]), .I1(n180), .CO(n22839));
    SB_LUT4 add_3394_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n6776[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_84_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n31024));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_84_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24664_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n31024), 
            .I2(IntegralLimit[14]), .I3(n29768), .O(n29756));
    defparam i24664_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_79_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n31019));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_79_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24388_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n29478));
    defparam i24388_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_102_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n31042));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_102_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n22179), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24879_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n31037), 
            .I2(IntegralLimit[11]), .I3(n29766), .O(n29971));
    defparam i24879_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i24396_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n31031), 
            .I2(IntegralLimit[13]), .I3(n29971), .O(n29486));
    defparam i24396_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_3394_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n22838));
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_82_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n31022));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_82_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24801_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n31022), 
            .I2(IntegralLimit[15]), .I3(n29486), .O(n29893));
    defparam i24801_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_108_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n31048));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_108_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3393_14_lut (.I0(GND_net), .I1(n6776[11]), .I2(n980), 
            .I3(n22837), .O(n6761[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24954_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n31048), 
            .I2(IntegralLimit[17]), .I3(n29893), .O(n30046));
    defparam i24954_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_73_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n31013));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_73_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n22179), .I0(GND_net), .I1(n1[18]), 
            .CO(n22180));
    SB_LUT4 i25011_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n31013), 
            .I2(IntegralLimit[19]), .I3(n30046), .O(n30103));
    defparam i25011_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_3393_13_lut (.I0(GND_net), .I1(n6776[10]), .I2(n907), 
            .I3(n22836), .O(n6761[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_70_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n31010));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_70_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3909));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3393_13 (.CI(n22836), .I0(n6776[10]), .I1(n907), .CO(n22837));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n22178), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3393_12_lut (.I0(GND_net), .I1(n6776[9]), .I2(n834), .I3(n22835), 
            .O(n6761[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24356_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n29446));
    defparam i24356_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_3393_12 (.CI(n22835), .I0(n6776[9]), .I1(n834), .CO(n22836));
    SB_LUT4 add_3393_11_lut (.I0(GND_net), .I1(n6776[8]), .I2(n761), .I3(n22834), 
            .O(n6761[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_11 (.CI(n22834), .I0(n6776[8]), .I1(n761), .CO(n22835));
    SB_LUT4 add_3393_10_lut (.I0(GND_net), .I1(n6776[7]), .I2(n688), .I3(n22833), 
            .O(n6761[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_10 (.CI(n22833), .I0(n6776[7]), .I1(n688), .CO(n22834));
    SB_LUT4 add_3393_9_lut (.I0(GND_net), .I1(n6776[6]), .I2(n615), .I3(n22832), 
            .O(n6761[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_9 (.CI(n22832), .I0(n6776[6]), .I1(n615), .CO(n22833));
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3909), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3911));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3912));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24837_3_lut (.I0(n6_adj_3912), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n29929));   // verilog/motorControl.v(31[10:34])
    defparam i24837_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24838_3_lut (.I0(n29929), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n29930));   // verilog/motorControl.v(31[10:34])
    defparam i24838_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24358_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n31031), 
            .I2(IntegralLimit[21]), .I3(n29762), .O(n29448));
    defparam i24358_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_3393_8_lut (.I0(GND_net), .I1(n6776[5]), .I2(n542), .I3(n22831), 
            .O(n6761[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_8 (.CI(n22831), .I0(n6776[5]), .I1(n542), .CO(n22832));
    SB_LUT4 i24777_4_lut (.I0(n24_adj_3911), .I1(n8_adj_3913), .I2(n31008), 
            .I3(n29446), .O(n29869));   // verilog/motorControl.v(31[10:34])
    defparam i24777_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24620_3_lut (.I0(n29930), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n29712));   // verilog/motorControl.v(31[10:34])
    defparam i24620_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3467 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n22178), .I0(GND_net), .I1(n1[17]), 
            .CO(n22179));
    SB_LUT4 i24920_3_lut (.I0(n4), .I1(\PID_CONTROLLER.integral [13]), .I2(n27), 
            .I3(GND_net), .O(n30012));   // verilog/motorControl.v(31[38:63])
    defparam i24920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3393_7_lut (.I0(GND_net), .I1(n6776[4]), .I2(n469), .I3(n22830), 
            .O(n6761[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24921_3_lut (.I0(n30012), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n30013));   // verilog/motorControl.v(31[38:63])
    defparam i24921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_3914));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24327_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n29417));
    defparam i24327_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3904), .I3(GND_net), 
            .O(n10_adj_3915));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3914), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_3916));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24330_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n29428), 
            .O(n29420));
    defparam i24330_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24989_4_lut (.I0(n30_adj_3916), .I1(n10_adj_3915), .I2(n35), 
            .I3(n29417), .O(n30081));   // verilog/motorControl.v(31[38:63])
    defparam i24989_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24856_3_lut (.I0(n30013), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n29948));   // verilog/motorControl.v(31[38:63])
    defparam i24856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25035_4_lut (.I0(n29948), .I1(n30081), .I2(n35), .I3(n29420), 
            .O(n30127));   // verilog/motorControl.v(31[38:63])
    defparam i25035_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25036_3_lut (.I0(n30127), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n30128));   // verilog/motorControl.v(31[38:63])
    defparam i25036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25020_3_lut (.I0(n30128), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n30112));   // verilog/motorControl.v(31[38:63])
    defparam i25020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7), .I3(GND_net), 
            .O(n6_adj_3917));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i24829_3_lut (.I0(n6_adj_3917), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21), .I3(GND_net), .O(n29921));   // verilog/motorControl.v(31[38:63])
    defparam i24829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24830_3_lut (.I0(n29921), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23), .I3(GND_net), .O(n29922));   // verilog/motorControl.v(31[38:63])
    defparam i24830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24319_4_lut (.I0(n43), .I1(n25_c), .I2(n23), .I3(n29434), 
            .O(n29409));
    defparam i24319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24779_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n29407), 
            .O(n29871));   // verilog/motorControl.v(31[38:63])
    defparam i24779_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24630_3_lut (.I0(n29922), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_c), .I3(GND_net), .O(n29722));   // verilog/motorControl.v(31[38:63])
    defparam i24630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24321_4_lut (.I0(n43), .I1(n41_adj_3918), .I2(n39), .I3(n30072), 
            .O(n29411));
    defparam i24321_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24934_4_lut (.I0(n29722), .I1(n29871), .I2(n45), .I3(n29409), 
            .O(n30026));   // verilog/motorControl.v(31[38:63])
    defparam i24934_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25006_3_lut (.I0(n30112), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_3918), .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[38:63])
    defparam i25006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24936_4_lut (.I0(n40), .I1(n30026), .I2(n45), .I3(n29411), 
            .O(n30028));   // verilog/motorControl.v(31[38:63])
    defparam i24936_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3919));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i24835_3_lut (.I0(n4_adj_3919), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n29927));   // verilog/motorControl.v(31[10:34])
    defparam i24835_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24836_3_lut (.I0(n29927), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n29928));   // verilog/motorControl.v(31[10:34])
    defparam i24836_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24390_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n31019), 
            .I2(IntegralLimit[16]), .I3(n29756), .O(n29480));
    defparam i24390_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i24974_4_lut (.I0(n30), .I1(n10), .I2(n31042), .I3(n29478), 
            .O(n30066));   // verilog/motorControl.v(31[10:34])
    defparam i24974_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24622_3_lut (.I0(n29928), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n29714));   // verilog/motorControl.v(31[10:34])
    defparam i24622_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3393_7 (.CI(n22830), .I0(n6776[4]), .I1(n469), .CO(n22831));
    SB_LUT4 add_3393_6_lut (.I0(GND_net), .I1(n6776[3]), .I2(n396), .I3(n22829), 
            .O(n6761[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3422_7_lut (.I0(GND_net), .I1(n27773), .I2(n490), .I3(n23136), 
            .O(n7142[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3422_6_lut (.I0(GND_net), .I1(n7150[3]), .I2(n417), .I3(n23135), 
            .O(n7142[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3422_6 (.CI(n23135), .I0(n7150[3]), .I1(n417), .CO(n23136));
    SB_LUT4 add_3422_5_lut (.I0(GND_net), .I1(n7150[2]), .I2(n344), .I3(n23134), 
            .O(n7142[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3422_5 (.CI(n23134), .I0(n7150[2]), .I1(n344), .CO(n23135));
    SB_LUT4 add_3422_4_lut (.I0(GND_net), .I1(n7150[1]), .I2(n271), .I3(n23133), 
            .O(n7142[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3422_4 (.CI(n23133), .I0(n7150[1]), .I1(n271), .CO(n23134));
    SB_LUT4 add_3422_3_lut (.I0(GND_net), .I1(n7150[0]), .I2(n198), .I3(n23132), 
            .O(n7142[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3422_3 (.CI(n23132), .I0(n7150[0]), .I1(n198), .CO(n23133));
    SB_LUT4 add_3422_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n7142[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3422_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3422_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n23132));
    SB_LUT4 add_3421_8_lut (.I0(GND_net), .I1(n7142[5]), .I2(n560), .I3(n23131), 
            .O(n7133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3421_7_lut (.I0(GND_net), .I1(n7142[4]), .I2(n487), .I3(n23130), 
            .O(n7133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_7 (.CI(n23130), .I0(n7142[4]), .I1(n487), .CO(n23131));
    SB_LUT4 add_3421_6_lut (.I0(GND_net), .I1(n7142[3]), .I2(n414), .I3(n23129), 
            .O(n7133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_6 (.CI(n23129), .I0(n7142[3]), .I1(n414), .CO(n23130));
    SB_LUT4 add_3421_5_lut (.I0(GND_net), .I1(n7142[2]), .I2(n341), .I3(n23128), 
            .O(n7133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_5 (.CI(n23128), .I0(n7142[2]), .I1(n341), .CO(n23129));
    SB_LUT4 add_3421_4_lut (.I0(GND_net), .I1(n7142[1]), .I2(n268), .I3(n23127), 
            .O(n7133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_4 (.CI(n23127), .I0(n7142[1]), .I1(n268), .CO(n23128));
    SB_LUT4 add_3421_3_lut (.I0(GND_net), .I1(n7142[0]), .I2(n195), .I3(n23126), 
            .O(n7133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_3 (.CI(n23126), .I0(n7142[0]), .I1(n195), .CO(n23127));
    SB_LUT4 add_3421_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n7133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3421_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3421_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n23126));
    SB_LUT4 add_3420_9_lut (.I0(GND_net), .I1(n7133[6]), .I2(n630), .I3(n23125), 
            .O(n7123[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3420_8_lut (.I0(GND_net), .I1(n7133[5]), .I2(n557), .I3(n23124), 
            .O(n7123[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_8 (.CI(n23124), .I0(n7133[5]), .I1(n557), .CO(n23125));
    SB_LUT4 i25023_4_lut (.I0(n29714), .I1(n30066), .I2(n31042), .I3(n29480), 
            .O(n30115));   // verilog/motorControl.v(31[10:34])
    defparam i25023_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3420_7_lut (.I0(GND_net), .I1(n7133[4]), .I2(n484), .I3(n23123), 
            .O(n7123[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_7 (.CI(n23123), .I0(n7133[4]), .I1(n484), .CO(n23124));
    SB_LUT4 add_3420_6_lut (.I0(GND_net), .I1(n7133[3]), .I2(n411), .I3(n23122), 
            .O(n7123[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_6 (.CI(n23122), .I0(n7133[3]), .I1(n411), .CO(n23123));
    SB_LUT4 add_3420_5_lut (.I0(GND_net), .I1(n7133[2]), .I2(n338), .I3(n23121), 
            .O(n7123[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_5 (.CI(n23121), .I0(n7133[2]), .I1(n338), .CO(n23122));
    SB_LUT4 add_3420_4_lut (.I0(GND_net), .I1(n7133[1]), .I2(n265), .I3(n23120), 
            .O(n7123[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_4 (.CI(n23120), .I0(n7133[1]), .I1(n265), .CO(n23121));
    SB_LUT4 add_3420_3_lut (.I0(GND_net), .I1(n7133[0]), .I2(n192), .I3(n23119), 
            .O(n7123[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_3 (.CI(n23119), .I0(n7133[0]), .I1(n192), .CO(n23120));
    SB_LUT4 add_3420_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n7123[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3420_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3420_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n23119));
    SB_LUT4 add_3419_10_lut (.I0(GND_net), .I1(n7123[7]), .I2(n700), .I3(n23118), 
            .O(n7112[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3419_9_lut (.I0(GND_net), .I1(n7123[6]), .I2(n627), .I3(n23117), 
            .O(n7112[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_9 (.CI(n23117), .I0(n7123[6]), .I1(n627), .CO(n23118));
    SB_LUT4 add_3419_8_lut (.I0(GND_net), .I1(n7123[5]), .I2(n554), .I3(n23116), 
            .O(n7112[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_8 (.CI(n23116), .I0(n7123[5]), .I1(n554), .CO(n23117));
    SB_LUT4 add_3419_7_lut (.I0(GND_net), .I1(n7123[4]), .I2(n481), .I3(n23115), 
            .O(n7112[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_7 (.CI(n23115), .I0(n7123[4]), .I1(n481), .CO(n23116));
    SB_LUT4 add_3419_6_lut (.I0(GND_net), .I1(n7123[3]), .I2(n408), .I3(n23114), 
            .O(n7112[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_6 (.CI(n23114), .I0(n7123[3]), .I1(n408), .CO(n23115));
    SB_LUT4 add_3419_5_lut (.I0(GND_net), .I1(n7123[2]), .I2(n335), .I3(n23113), 
            .O(n7112[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_5 (.CI(n23113), .I0(n7123[2]), .I1(n335), .CO(n23114));
    SB_LUT4 add_3419_4_lut (.I0(GND_net), .I1(n7123[1]), .I2(n262), .I3(n23112), 
            .O(n7112[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_4 (.CI(n23112), .I0(n7123[1]), .I1(n262), .CO(n23113));
    SB_LUT4 add_3419_3_lut (.I0(GND_net), .I1(n7123[0]), .I2(n189), .I3(n23111), 
            .O(n7112[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_3 (.CI(n23111), .I0(n7123[0]), .I1(n189), .CO(n23112));
    SB_LUT4 add_3419_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n7112[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3419_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3419_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n23111));
    SB_LUT4 add_3418_11_lut (.I0(GND_net), .I1(n7112[8]), .I2(n770), .I3(n23110), 
            .O(n7100[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3418_10_lut (.I0(GND_net), .I1(n7112[7]), .I2(n697), .I3(n23109), 
            .O(n7100[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_10 (.CI(n23109), .I0(n7112[7]), .I1(n697), .CO(n23110));
    SB_LUT4 add_3418_9_lut (.I0(GND_net), .I1(n7112[6]), .I2(n624), .I3(n23108), 
            .O(n7100[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_9 (.CI(n23108), .I0(n7112[6]), .I1(n624), .CO(n23109));
    SB_LUT4 add_3418_8_lut (.I0(GND_net), .I1(n7112[5]), .I2(n551), .I3(n23107), 
            .O(n7100[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_8 (.CI(n23107), .I0(n7112[5]), .I1(n551), .CO(n23108));
    SB_LUT4 add_3418_7_lut (.I0(GND_net), .I1(n7112[4]), .I2(n478), .I3(n23106), 
            .O(n7100[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_7 (.CI(n23106), .I0(n7112[4]), .I1(n478), .CO(n23107));
    SB_LUT4 add_3418_6_lut (.I0(GND_net), .I1(n7112[3]), .I2(n405), .I3(n23105), 
            .O(n7100[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_6 (.CI(n23105), .I0(n7112[3]), .I1(n405), .CO(n23106));
    SB_LUT4 add_3418_5_lut (.I0(GND_net), .I1(n7112[2]), .I2(n332), .I3(n23104), 
            .O(n7100[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_5 (.CI(n23104), .I0(n7112[2]), .I1(n332), .CO(n23105));
    SB_LUT4 add_3418_4_lut (.I0(GND_net), .I1(n7112[1]), .I2(n259), .I3(n23103), 
            .O(n7100[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_4 (.CI(n23103), .I0(n7112[1]), .I1(n259), .CO(n23104));
    SB_LUT4 add_3418_3_lut (.I0(GND_net), .I1(n7112[0]), .I2(n186), .I3(n23102), 
            .O(n7100[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_3 (.CI(n23102), .I0(n7112[0]), .I1(n186), .CO(n23103));
    SB_LUT4 add_3418_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n7100[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3418_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3418_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n23102));
    SB_LUT4 add_3417_12_lut (.I0(GND_net), .I1(n7100[9]), .I2(n840), .I3(n23101), 
            .O(n7087[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_11_lut (.I0(GND_net), .I1(n7100[8]), .I2(n767), .I3(n23100), 
            .O(n7087[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_11 (.CI(n23100), .I0(n7100[8]), .I1(n767), .CO(n23101));
    SB_LUT4 add_3417_10_lut (.I0(GND_net), .I1(n7100[7]), .I2(n694), .I3(n23099), 
            .O(n7087[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_10 (.CI(n23099), .I0(n7100[7]), .I1(n694), .CO(n23100));
    SB_LUT4 add_3417_9_lut (.I0(GND_net), .I1(n7100[6]), .I2(n621), .I3(n23098), 
            .O(n7087[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_9 (.CI(n23098), .I0(n7100[6]), .I1(n621), .CO(n23099));
    SB_LUT4 add_3417_8_lut (.I0(GND_net), .I1(n7100[5]), .I2(n548), .I3(n23097), 
            .O(n7087[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_8 (.CI(n23097), .I0(n7100[5]), .I1(n548), .CO(n23098));
    SB_LUT4 add_3417_7_lut (.I0(GND_net), .I1(n7100[4]), .I2(n475), .I3(n23096), 
            .O(n7087[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_7 (.CI(n23096), .I0(n7100[4]), .I1(n475), .CO(n23097));
    SB_LUT4 add_3417_6_lut (.I0(GND_net), .I1(n7100[3]), .I2(n402), .I3(n23095), 
            .O(n7087[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_6 (.CI(n23095), .I0(n7100[3]), .I1(n402), .CO(n23096));
    SB_LUT4 add_3417_5_lut (.I0(GND_net), .I1(n7100[2]), .I2(n329), .I3(n23094), 
            .O(n7087[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_5 (.CI(n23094), .I0(n7100[2]), .I1(n329), .CO(n23095));
    SB_LUT4 add_3417_4_lut (.I0(GND_net), .I1(n7100[1]), .I2(n256_adj_3903), 
            .I3(n23093), .O(n7087[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_4 (.CI(n23093), .I0(n7100[1]), .I1(n256_adj_3903), 
            .CO(n23094));
    SB_LUT4 add_3417_3_lut (.I0(GND_net), .I1(n7100[0]), .I2(n183), .I3(n23092), 
            .O(n7087[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_3 (.CI(n23092), .I0(n7100[0]), .I1(n183), .CO(n23093));
    SB_LUT4 add_3417_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n7087[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n23092));
    SB_LUT4 add_3416_13_lut (.I0(GND_net), .I1(n7087[10]), .I2(n910), 
            .I3(n23091), .O(n7073[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_12_lut (.I0(GND_net), .I1(n7087[9]), .I2(n837), .I3(n23090), 
            .O(n7073[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_12 (.CI(n23090), .I0(n7087[9]), .I1(n837), .CO(n23091));
    SB_LUT4 add_3416_11_lut (.I0(GND_net), .I1(n7087[8]), .I2(n764), .I3(n23089), 
            .O(n7073[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_11 (.CI(n23089), .I0(n7087[8]), .I1(n764), .CO(n23090));
    SB_LUT4 add_3416_10_lut (.I0(GND_net), .I1(n7087[7]), .I2(n691), .I3(n23088), 
            .O(n7073[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_10 (.CI(n23088), .I0(n7087[7]), .I1(n691), .CO(n23089));
    SB_LUT4 add_3416_9_lut (.I0(GND_net), .I1(n7087[6]), .I2(n618), .I3(n23087), 
            .O(n7073[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25024_3_lut (.I0(n30115), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n30116));   // verilog/motorControl.v(31[10:34])
    defparam i25024_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3416_9 (.CI(n23087), .I0(n7087[6]), .I1(n618), .CO(n23088));
    SB_LUT4 add_3416_8_lut (.I0(GND_net), .I1(n7087[5]), .I2(n545_adj_3920), 
            .I3(n23086), .O(n7073[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_8 (.CI(n23086), .I0(n7087[5]), .I1(n545_adj_3920), 
            .CO(n23087));
    SB_LUT4 add_3416_7_lut (.I0(GND_net), .I1(n7087[4]), .I2(n472_adj_3921), 
            .I3(n23085), .O(n7073[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_7 (.CI(n23085), .I0(n7087[4]), .I1(n472_adj_3921), 
            .CO(n23086));
    SB_LUT4 add_3416_6_lut (.I0(GND_net), .I1(n7087[3]), .I2(n399_adj_3922), 
            .I3(n23084), .O(n7073[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_6 (.CI(n23084), .I0(n7087[3]), .I1(n399_adj_3922), 
            .CO(n23085));
    SB_LUT4 add_3416_5_lut (.I0(GND_net), .I1(n7087[2]), .I2(n326_adj_3923), 
            .I3(n23083), .O(n7073[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_5 (.CI(n23083), .I0(n7087[2]), .I1(n326_adj_3923), 
            .CO(n23084));
    SB_LUT4 add_3416_4_lut (.I0(GND_net), .I1(n7087[1]), .I2(n253_adj_3924), 
            .I3(n23082), .O(n7073[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_4 (.CI(n23082), .I0(n7087[1]), .I1(n253_adj_3924), 
            .CO(n23083));
    SB_LUT4 add_3416_3_lut (.I0(GND_net), .I1(n7087[0]), .I2(n180_adj_3925), 
            .I3(n23081), .O(n7073[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_3 (.CI(n23081), .I0(n7087[0]), .I1(n180_adj_3925), 
            .CO(n23082));
    SB_LUT4 add_3416_2_lut (.I0(GND_net), .I1(n38_adj_3926), .I2(n107_adj_3927), 
            .I3(GND_net), .O(n7073[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_2 (.CI(GND_net), .I0(n38_adj_3926), .I1(n107_adj_3927), 
            .CO(n23081));
    SB_LUT4 add_3415_14_lut (.I0(GND_net), .I1(n7073[11]), .I2(n980_adj_3928), 
            .I3(n23080), .O(n7058[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3415_13_lut (.I0(GND_net), .I1(n7073[10]), .I2(n907_adj_3929), 
            .I3(n23079), .O(n7058[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_13 (.CI(n23079), .I0(n7073[10]), .I1(n907_adj_3929), 
            .CO(n23080));
    SB_LUT4 add_3415_12_lut (.I0(GND_net), .I1(n7073[9]), .I2(n834_adj_3930), 
            .I3(n23078), .O(n7058[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_12 (.CI(n23078), .I0(n7073[9]), .I1(n834_adj_3930), 
            .CO(n23079));
    SB_LUT4 add_3415_11_lut (.I0(GND_net), .I1(n7073[8]), .I2(n761_adj_3931), 
            .I3(n23077), .O(n7058[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_11 (.CI(n23077), .I0(n7073[8]), .I1(n761_adj_3931), 
            .CO(n23078));
    SB_LUT4 add_3415_10_lut (.I0(GND_net), .I1(n7073[7]), .I2(n688_adj_3932), 
            .I3(n23076), .O(n7058[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_10 (.CI(n23076), .I0(n7073[7]), .I1(n688_adj_3932), 
            .CO(n23077));
    SB_LUT4 add_3415_9_lut (.I0(GND_net), .I1(n7073[6]), .I2(n615_adj_3933), 
            .I3(n23075), .O(n7058[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24998_3_lut (.I0(n30116), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n30090));   // verilog/motorControl.v(31[10:34])
    defparam i24998_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3415_9 (.CI(n23075), .I0(n7073[6]), .I1(n615_adj_3933), 
            .CO(n23076));
    SB_LUT4 add_3415_8_lut (.I0(GND_net), .I1(n7073[5]), .I2(n542_adj_3934), 
            .I3(n23074), .O(n7058[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_8 (.CI(n23074), .I0(n7073[5]), .I1(n542_adj_3934), 
            .CO(n23075));
    SB_LUT4 add_3415_7_lut (.I0(GND_net), .I1(n7073[4]), .I2(n469_adj_3935), 
            .I3(n23073), .O(n7058[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_7 (.CI(n23073), .I0(n7073[4]), .I1(n469_adj_3935), 
            .CO(n23074));
    SB_LUT4 add_3415_6_lut (.I0(GND_net), .I1(n7073[3]), .I2(n396_adj_3936), 
            .I3(n23072), .O(n7058[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_6 (.CI(n23072), .I0(n7073[3]), .I1(n396_adj_3936), 
            .CO(n23073));
    SB_LUT4 add_3415_5_lut (.I0(GND_net), .I1(n7073[2]), .I2(n323), .I3(n23071), 
            .O(n7058[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_5 (.CI(n23071), .I0(n7073[2]), .I1(n323), .CO(n23072));
    SB_LUT4 add_3415_4_lut (.I0(GND_net), .I1(n7073[1]), .I2(n250), .I3(n23070), 
            .O(n7058[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_4 (.CI(n23070), .I0(n7073[1]), .I1(n250), .CO(n23071));
    SB_LUT4 add_3415_3_lut (.I0(GND_net), .I1(n7073[0]), .I2(n177), .I3(n23069), 
            .O(n7058[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_3 (.CI(n23069), .I0(n7073[0]), .I1(n177), .CO(n23070));
    SB_LUT4 add_3415_2_lut (.I0(GND_net), .I1(n35_adj_3937), .I2(n104), 
            .I3(GND_net), .O(n7058[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3415_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3415_2 (.CI(GND_net), .I0(n35_adj_3937), .I1(n104), .CO(n23069));
    SB_LUT4 add_3414_15_lut (.I0(GND_net), .I1(n7058[12]), .I2(n1050), 
            .I3(n23068), .O(n7042[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3414_14_lut (.I0(GND_net), .I1(n7058[11]), .I2(n977), 
            .I3(n23067), .O(n7042[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_14 (.CI(n23067), .I0(n7058[11]), .I1(n977), .CO(n23068));
    SB_LUT4 add_3414_13_lut (.I0(GND_net), .I1(n7058[10]), .I2(n904), 
            .I3(n23066), .O(n7042[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_13 (.CI(n23066), .I0(n7058[10]), .I1(n904), .CO(n23067));
    SB_LUT4 add_3414_12_lut (.I0(GND_net), .I1(n7058[9]), .I2(n831), .I3(n23065), 
            .O(n7042[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_12 (.CI(n23065), .I0(n7058[9]), .I1(n831), .CO(n23066));
    SB_LUT4 add_3414_11_lut (.I0(GND_net), .I1(n7058[8]), .I2(n758), .I3(n23064), 
            .O(n7042[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_11 (.CI(n23064), .I0(n7058[8]), .I1(n758), .CO(n23065));
    SB_LUT4 add_3414_10_lut (.I0(GND_net), .I1(n7058[7]), .I2(n685), .I3(n23063), 
            .O(n7042[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_10 (.CI(n23063), .I0(n7058[7]), .I1(n685), .CO(n23064));
    SB_LUT4 add_3414_9_lut (.I0(GND_net), .I1(n7058[6]), .I2(n612), .I3(n23062), 
            .O(n7042[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_9 (.CI(n23062), .I0(n7058[6]), .I1(n612), .CO(n23063));
    SB_LUT4 add_3414_8_lut (.I0(GND_net), .I1(n7058[5]), .I2(n539), .I3(n23061), 
            .O(n7042[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24382_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n31010), 
            .I2(IntegralLimit[21]), .I3(n30103), .O(n29472));
    defparam i24382_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_3414_8 (.CI(n23061), .I0(n7058[5]), .I1(n539), .CO(n23062));
    SB_LUT4 add_3414_7_lut (.I0(GND_net), .I1(n7058[4]), .I2(n466), .I3(n23060), 
            .O(n7042[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_7 (.CI(n23060), .I0(n7058[4]), .I1(n466), .CO(n23061));
    SB_LUT4 add_3414_6_lut (.I0(GND_net), .I1(n7058[3]), .I2(n393), .I3(n23059), 
            .O(n7042[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_6 (.CI(n23059), .I0(n7058[3]), .I1(n393), .CO(n23060));
    SB_LUT4 add_3414_5_lut (.I0(GND_net), .I1(n7058[2]), .I2(n320), .I3(n23058), 
            .O(n7042[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_5 (.CI(n23058), .I0(n7058[2]), .I1(n320), .CO(n23059));
    SB_LUT4 add_3414_4_lut (.I0(GND_net), .I1(n7058[1]), .I2(n247), .I3(n23057), 
            .O(n7042[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_4 (.CI(n23057), .I0(n7058[1]), .I1(n247), .CO(n23058));
    SB_LUT4 add_3414_3_lut (.I0(GND_net), .I1(n7058[0]), .I2(n174), .I3(n23056), 
            .O(n7042[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_3 (.CI(n23056), .I0(n7058[0]), .I1(n174), .CO(n23057));
    SB_LUT4 add_3414_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n7042[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3414_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3414_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n23056));
    SB_LUT4 add_3413_16_lut (.I0(GND_net), .I1(n7042[13]), .I2(n1120), 
            .I3(n23055), .O(n7025[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3413_15_lut (.I0(GND_net), .I1(n7042[12]), .I2(n1047), 
            .I3(n23054), .O(n7025[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_15 (.CI(n23054), .I0(n7042[12]), .I1(n1047), .CO(n23055));
    SB_LUT4 add_3413_14_lut (.I0(GND_net), .I1(n7042[11]), .I2(n974), 
            .I3(n23053), .O(n7025[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_14 (.CI(n23053), .I0(n7042[11]), .I1(n974), .CO(n23054));
    SB_LUT4 add_3413_13_lut (.I0(GND_net), .I1(n7042[10]), .I2(n901), 
            .I3(n23052), .O(n7025[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_13 (.CI(n23052), .I0(n7042[10]), .I1(n901), .CO(n23053));
    SB_LUT4 add_3413_12_lut (.I0(GND_net), .I1(n7042[9]), .I2(n828), .I3(n23051), 
            .O(n7025[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_12 (.CI(n23051), .I0(n7042[9]), .I1(n828), .CO(n23052));
    SB_LUT4 add_3413_11_lut (.I0(GND_net), .I1(n7042[8]), .I2(n755), .I3(n23050), 
            .O(n7025[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_11 (.CI(n23050), .I0(n7042[8]), .I1(n755), .CO(n23051));
    SB_LUT4 add_3413_10_lut (.I0(GND_net), .I1(n7042[7]), .I2(n682), .I3(n23049), 
            .O(n7025[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_10 (.CI(n23049), .I0(n7042[7]), .I1(n682), .CO(n23050));
    SB_LUT4 add_3413_9_lut (.I0(GND_net), .I1(n7042[6]), .I2(n609), .I3(n23048), 
            .O(n7025[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_9 (.CI(n23048), .I0(n7042[6]), .I1(n609), .CO(n23049));
    SB_CARRY add_3393_6 (.CI(n22829), .I0(n6776[3]), .I1(n396), .CO(n22830));
    SB_LUT4 add_3413_8_lut (.I0(GND_net), .I1(n7042[5]), .I2(n536), .I3(n23047), 
            .O(n7025[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_8 (.CI(n23047), .I0(n7042[5]), .I1(n536), .CO(n23048));
    SB_LUT4 add_3413_7_lut (.I0(GND_net), .I1(n7042[4]), .I2(n463), .I3(n23046), 
            .O(n7025[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_7 (.CI(n23046), .I0(n7042[4]), .I1(n463), .CO(n23047));
    SB_LUT4 add_3413_6_lut (.I0(GND_net), .I1(n7042[3]), .I2(n390), .I3(n23045), 
            .O(n7025[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_6 (.CI(n23045), .I0(n7042[3]), .I1(n390), .CO(n23046));
    SB_LUT4 add_3413_5_lut (.I0(GND_net), .I1(n7042[2]), .I2(n317), .I3(n23044), 
            .O(n7025[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_5 (.CI(n23044), .I0(n7042[2]), .I1(n317), .CO(n23045));
    SB_LUT4 add_3413_4_lut (.I0(GND_net), .I1(n7042[1]), .I2(n244), .I3(n23043), 
            .O(n7025[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_4 (.CI(n23043), .I0(n7042[1]), .I1(n244), .CO(n23044));
    SB_LUT4 add_3413_3_lut (.I0(GND_net), .I1(n7042[0]), .I2(n171), .I3(n23042), 
            .O(n7025[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_3 (.CI(n23042), .I0(n7042[0]), .I1(n171), .CO(n23043));
    SB_LUT4 add_3413_2_lut (.I0(GND_net), .I1(n29_adj_3938), .I2(n98), 
            .I3(GND_net), .O(n7025[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3413_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3413_2 (.CI(GND_net), .I0(n29_adj_3938), .I1(n98), .CO(n23042));
    SB_LUT4 add_3412_17_lut (.I0(GND_net), .I1(n7025[14]), .I2(GND_net), 
            .I3(n23041), .O(n7007[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3412_16_lut (.I0(GND_net), .I1(n7025[13]), .I2(n1117), 
            .I3(n23040), .O(n7007[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_16 (.CI(n23040), .I0(n7025[13]), .I1(n1117), .CO(n23041));
    SB_LUT4 add_3412_15_lut (.I0(GND_net), .I1(n7025[12]), .I2(n1044), 
            .I3(n23039), .O(n7007[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_15 (.CI(n23039), .I0(n7025[12]), .I1(n1044), .CO(n23040));
    SB_LUT4 add_3412_14_lut (.I0(GND_net), .I1(n7025[11]), .I2(n971), 
            .I3(n23038), .O(n7007[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_14 (.CI(n23038), .I0(n7025[11]), .I1(n971), .CO(n23039));
    SB_LUT4 add_3412_13_lut (.I0(GND_net), .I1(n7025[10]), .I2(n898), 
            .I3(n23037), .O(n7007[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_13 (.CI(n23037), .I0(n7025[10]), .I1(n898), .CO(n23038));
    SB_LUT4 add_3412_12_lut (.I0(GND_net), .I1(n7025[9]), .I2(n825), .I3(n23036), 
            .O(n7007[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_12 (.CI(n23036), .I0(n7025[9]), .I1(n825), .CO(n23037));
    SB_LUT4 add_3412_11_lut (.I0(GND_net), .I1(n7025[8]), .I2(n752), .I3(n23035), 
            .O(n7007[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_11 (.CI(n23035), .I0(n7025[8]), .I1(n752), .CO(n23036));
    SB_LUT4 add_3412_10_lut (.I0(GND_net), .I1(n7025[7]), .I2(n679), .I3(n23034), 
            .O(n7007[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_10 (.CI(n23034), .I0(n7025[7]), .I1(n679), .CO(n23035));
    SB_LUT4 add_3412_9_lut (.I0(GND_net), .I1(n7025[6]), .I2(n606), .I3(n23033), 
            .O(n7007[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_9 (.CI(n23033), .I0(n7025[6]), .I1(n606), .CO(n23034));
    SB_LUT4 add_3412_8_lut (.I0(GND_net), .I1(n7025[5]), .I2(n533), .I3(n23032), 
            .O(n7007[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_8 (.CI(n23032), .I0(n7025[5]), .I1(n533), .CO(n23033));
    SB_LUT4 add_3412_7_lut (.I0(GND_net), .I1(n7025[4]), .I2(n460), .I3(n23031), 
            .O(n7007[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_7 (.CI(n23031), .I0(n7025[4]), .I1(n460), .CO(n23032));
    SB_LUT4 add_3412_6_lut (.I0(GND_net), .I1(n7025[3]), .I2(n387), .I3(n23030), 
            .O(n7007[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_6 (.CI(n23030), .I0(n7025[3]), .I1(n387), .CO(n23031));
    SB_LUT4 add_3412_5_lut (.I0(GND_net), .I1(n7025[2]), .I2(n314), .I3(n23029), 
            .O(n7007[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_5 (.CI(n23029), .I0(n7025[2]), .I1(n314), .CO(n23030));
    SB_LUT4 add_3412_4_lut (.I0(GND_net), .I1(n7025[1]), .I2(n241), .I3(n23028), 
            .O(n7007[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_4 (.CI(n23028), .I0(n7025[1]), .I1(n241), .CO(n23029));
    SB_LUT4 add_3412_3_lut (.I0(GND_net), .I1(n7025[0]), .I2(n168), .I3(n23027), 
            .O(n7007[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_3 (.CI(n23027), .I0(n7025[0]), .I1(n168), .CO(n23028));
    SB_LUT4 add_3412_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7007[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3412_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3412_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n23027));
    SB_LUT4 add_3411_18_lut (.I0(GND_net), .I1(n7007[15]), .I2(GND_net), 
            .I3(n23026), .O(n6988[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3411_17_lut (.I0(GND_net), .I1(n7007[14]), .I2(GND_net), 
            .I3(n23025), .O(n6988[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3393_5_lut (.I0(GND_net), .I1(n6776[2]), .I2(n323_adj_3939), 
            .I3(n22828), .O(n6761[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_5 (.CI(n22828), .I0(n6776[2]), .I1(n323_adj_3939), 
            .CO(n22829));
    SB_CARRY add_3411_17 (.CI(n23025), .I0(n7007[14]), .I1(GND_net), .CO(n23026));
    SB_LUT4 add_3411_16_lut (.I0(GND_net), .I1(n7007[13]), .I2(n1114), 
            .I3(n23024), .O(n6988[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_16 (.CI(n23024), .I0(n7007[13]), .I1(n1114), .CO(n23025));
    SB_LUT4 add_3411_15_lut (.I0(GND_net), .I1(n7007[12]), .I2(n1041), 
            .I3(n23023), .O(n6988[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_15 (.CI(n23023), .I0(n7007[12]), .I1(n1041), .CO(n23024));
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_68_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n31008));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_68_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3411_14_lut (.I0(GND_net), .I1(n7007[11]), .I2(n968), 
            .I3(n23022), .O(n6988[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_14 (.CI(n23022), .I0(n7007[11]), .I1(n968), .CO(n23023));
    SB_LUT4 add_3411_13_lut (.I0(GND_net), .I1(n7007[10]), .I2(n895), 
            .I3(n23021), .O(n6988[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_13 (.CI(n23021), .I0(n7007[10]), .I1(n895), .CO(n23022));
    SB_LUT4 add_3411_12_lut (.I0(GND_net), .I1(n7007[9]), .I2(n822), .I3(n23020), 
            .O(n6988[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_12 (.CI(n23020), .I0(n7007[9]), .I1(n822), .CO(n23021));
    SB_LUT4 add_3411_11_lut (.I0(GND_net), .I1(n7007[8]), .I2(n749), .I3(n23019), 
            .O(n6988[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_11 (.CI(n23019), .I0(n7007[8]), .I1(n749), .CO(n23020));
    SB_LUT4 add_3411_10_lut (.I0(GND_net), .I1(n7007[7]), .I2(n676), .I3(n23018), 
            .O(n6988[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_10 (.CI(n23018), .I0(n7007[7]), .I1(n676), .CO(n23019));
    SB_LUT4 add_3411_9_lut (.I0(GND_net), .I1(n7007[6]), .I2(n603), .I3(n23017), 
            .O(n6988[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_9 (.CI(n23017), .I0(n7007[6]), .I1(n603), .CO(n23018));
    SB_LUT4 add_3411_8_lut (.I0(GND_net), .I1(n7007[5]), .I2(n530), .I3(n23016), 
            .O(n6988[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24930_4_lut (.I0(n29712), .I1(n29869), .I2(n31008), .I3(n29448), 
            .O(n30022));   // verilog/motorControl.v(31[10:34])
    defparam i24930_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24628_3_lut (.I0(n30090), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n29720));   // verilog/motorControl.v(31[10:34])
    defparam i24628_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24937_3_lut (.I0(n30028), .I1(\PID_CONTROLLER.integral_23__N_3467 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3466 ));   // verilog/motorControl.v(31[38:63])
    defparam i24937_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3411_8 (.CI(n23016), .I0(n7007[5]), .I1(n530), .CO(n23017));
    SB_LUT4 add_3411_7_lut (.I0(GND_net), .I1(n7007[4]), .I2(n457), .I3(n23015), 
            .O(n6988[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_7 (.CI(n23015), .I0(n7007[4]), .I1(n457), .CO(n23016));
    SB_LUT4 add_3411_6_lut (.I0(GND_net), .I1(n7007[3]), .I2(n384), .I3(n23014), 
            .O(n6988[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_6 (.CI(n23014), .I0(n7007[3]), .I1(n384), .CO(n23015));
    SB_LUT4 add_3411_5_lut (.I0(GND_net), .I1(n7007[2]), .I2(n311), .I3(n23013), 
            .O(n6988[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_5 (.CI(n23013), .I0(n7007[2]), .I1(n311), .CO(n23014));
    SB_LUT4 add_3411_4_lut (.I0(GND_net), .I1(n7007[1]), .I2(n238), .I3(n23012), 
            .O(n6988[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_4 (.CI(n23012), .I0(n7007[1]), .I1(n238), .CO(n23013));
    SB_LUT4 add_3411_3_lut (.I0(GND_net), .I1(n7007[0]), .I2(n165), .I3(n23011), 
            .O(n6988[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_3 (.CI(n23011), .I0(n7007[0]), .I1(n165), .CO(n23012));
    SB_LUT4 add_3411_2_lut (.I0(GND_net), .I1(n23_adj_3940), .I2(n92), 
            .I3(GND_net), .O(n6988[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3411_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3411_2 (.CI(GND_net), .I0(n23_adj_3940), .I1(n92), .CO(n23011));
    SB_LUT4 add_3410_19_lut (.I0(GND_net), .I1(n6988[16]), .I2(GND_net), 
            .I3(n23010), .O(n6968[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3410_18_lut (.I0(GND_net), .I1(n6988[15]), .I2(GND_net), 
            .I3(n23009), .O(n6968[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_18 (.CI(n23009), .I0(n6988[15]), .I1(GND_net), .CO(n23010));
    SB_LUT4 add_3410_17_lut (.I0(GND_net), .I1(n6988[14]), .I2(GND_net), 
            .I3(n23008), .O(n6968[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_17 (.CI(n23008), .I0(n6988[14]), .I1(GND_net), .CO(n23009));
    SB_LUT4 add_3410_16_lut (.I0(GND_net), .I1(n6988[13]), .I2(n1111), 
            .I3(n23007), .O(n6968[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_16 (.CI(n23007), .I0(n6988[13]), .I1(n1111), .CO(n23008));
    SB_LUT4 add_3410_15_lut (.I0(GND_net), .I1(n6988[12]), .I2(n1038), 
            .I3(n23006), .O(n6968[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_15 (.CI(n23006), .I0(n6988[12]), .I1(n1038), .CO(n23007));
    SB_LUT4 add_3410_14_lut (.I0(GND_net), .I1(n6988[11]), .I2(n965), 
            .I3(n23005), .O(n6968[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_14 (.CI(n23005), .I0(n6988[11]), .I1(n965), .CO(n23006));
    SB_LUT4 add_3410_13_lut (.I0(GND_net), .I1(n6988[10]), .I2(n892), 
            .I3(n23004), .O(n6968[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_13 (.CI(n23004), .I0(n6988[10]), .I1(n892), .CO(n23005));
    SB_LUT4 add_3410_12_lut (.I0(GND_net), .I1(n6988[9]), .I2(n819), .I3(n23003), 
            .O(n6968[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_12 (.CI(n23003), .I0(n6988[9]), .I1(n819), .CO(n23004));
    SB_LUT4 i24982_4_lut (.I0(n29720), .I1(n30022), .I2(n31008), .I3(n29472), 
            .O(n30074));   // verilog/motorControl.v(31[10:34])
    defparam i24982_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3410_11_lut (.I0(GND_net), .I1(n6988[8]), .I2(n746), .I3(n23002), 
            .O(n6968[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n30074), .I1(\PID_CONTROLLER.integral_23__N_3466 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3464 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3393_4_lut (.I0(GND_net), .I1(n6776[1]), .I2(n250_adj_3941), 
            .I3(n22827), .O(n6761[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_4 (.CI(n22827), .I0(n6776[1]), .I1(n250_adj_3941), 
            .CO(n22828));
    SB_LUT4 add_3393_3_lut (.I0(GND_net), .I1(n6776[0]), .I2(n177_adj_3942), 
            .I3(n22826), .O(n6761[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_3 (.CI(n22826), .I0(n6776[0]), .I1(n177_adj_3942), 
            .CO(n22827));
    SB_LUT4 add_3393_2_lut (.I0(GND_net), .I1(n35_adj_3943), .I2(n104_adj_3944), 
            .I3(GND_net), .O(n6761[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3393_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3393_2 (.CI(GND_net), .I0(n35_adj_3943), .I1(n104_adj_3944), 
            .CO(n22826));
    SB_LUT4 add_3392_15_lut (.I0(GND_net), .I1(n6761[12]), .I2(n1050_adj_3945), 
            .I3(n22825), .O(n6745[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_11 (.CI(n23002), .I0(n6988[8]), .I1(n746), .CO(n23003));
    SB_LUT4 add_3410_10_lut (.I0(GND_net), .I1(n6988[7]), .I2(n673), .I3(n23001), 
            .O(n6968[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3392_14_lut (.I0(GND_net), .I1(n6761[11]), .I2(n977_adj_3946), 
            .I3(n22824), .O(n6745[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_10 (.CI(n23001), .I0(n6988[7]), .I1(n673), .CO(n23002));
    SB_LUT4 add_3410_9_lut (.I0(GND_net), .I1(n6988[6]), .I2(n600), .I3(n23000), 
            .O(n6968[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_14 (.CI(n22824), .I0(n6761[11]), .I1(n977_adj_3946), 
            .CO(n22825));
    SB_CARRY add_3410_9 (.CI(n23000), .I0(n6988[6]), .I1(n600), .CO(n23001));
    SB_LUT4 add_3392_13_lut (.I0(GND_net), .I1(n6761[10]), .I2(n904_adj_3947), 
            .I3(n22823), .O(n6745[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_13 (.CI(n22823), .I0(n6761[10]), .I1(n904_adj_3947), 
            .CO(n22824));
    SB_LUT4 add_3392_12_lut (.I0(GND_net), .I1(n6761[9]), .I2(n831_adj_3948), 
            .I3(n22822), .O(n6745[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3410_8_lut (.I0(GND_net), .I1(n6988[5]), .I2(n527), .I3(n22999), 
            .O(n6968[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_12 (.CI(n22822), .I0(n6761[9]), .I1(n831_adj_3948), 
            .CO(n22823));
    SB_CARRY add_3410_8 (.CI(n22999), .I0(n6988[5]), .I1(n527), .CO(n23000));
    SB_LUT4 add_3392_11_lut (.I0(GND_net), .I1(n6761[8]), .I2(n758_adj_3949), 
            .I3(n22821), .O(n6745[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_11 (.CI(n22821), .I0(n6761[8]), .I1(n758_adj_3949), 
            .CO(n22822));
    SB_LUT4 add_3392_10_lut (.I0(GND_net), .I1(n6761[7]), .I2(n685_adj_3950), 
            .I3(n22820), .O(n6745[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_10 (.CI(n22820), .I0(n6761[7]), .I1(n685_adj_3950), 
            .CO(n22821));
    SB_LUT4 add_3392_9_lut (.I0(GND_net), .I1(n6761[6]), .I2(n612_adj_3951), 
            .I3(n22819), .O(n6745[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_9 (.CI(n22819), .I0(n6761[6]), .I1(n612_adj_3951), 
            .CO(n22820));
    SB_LUT4 add_3392_8_lut (.I0(GND_net), .I1(n6761[5]), .I2(n539_adj_3952), 
            .I3(n22818), .O(n6745[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3410_7_lut (.I0(GND_net), .I1(n6988[4]), .I2(n454), .I3(n22998), 
            .O(n6968[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_8 (.CI(n22818), .I0(n6761[5]), .I1(n539_adj_3952), 
            .CO(n22819));
    SB_LUT4 add_3392_7_lut (.I0(GND_net), .I1(n6761[4]), .I2(n466_adj_3953), 
            .I3(n22817), .O(n6745[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_7 (.CI(n22817), .I0(n6761[4]), .I1(n466_adj_3953), 
            .CO(n22818));
    SB_LUT4 add_3392_6_lut (.I0(GND_net), .I1(n6761[3]), .I2(n393_adj_3954), 
            .I3(n22816), .O(n6745[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_6 (.CI(n22816), .I0(n6761[3]), .I1(n393_adj_3954), 
            .CO(n22817));
    SB_LUT4 add_3392_5_lut (.I0(GND_net), .I1(n6761[2]), .I2(n320_adj_3955), 
            .I3(n22815), .O(n6745[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_5 (.CI(n22815), .I0(n6761[2]), .I1(n320_adj_3955), 
            .CO(n22816));
    SB_CARRY add_3410_7 (.CI(n22998), .I0(n6988[4]), .I1(n454), .CO(n22999));
    SB_LUT4 add_3410_6_lut (.I0(GND_net), .I1(n6988[3]), .I2(n381), .I3(n22997), 
            .O(n6968[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3392_4_lut (.I0(GND_net), .I1(n6761[1]), .I2(n247_adj_3956), 
            .I3(n22814), .O(n6745[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_561_i21_3_lut (.I0(n155[20]), .I1(PWMLimit[20]), .I2(n256), 
            .I3(GND_net), .O(n2554[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i21_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3410_6 (.CI(n22997), .I0(n6988[3]), .I1(n381), .CO(n22998));
    SB_CARRY add_3392_4 (.CI(n22814), .I0(n6761[1]), .I1(n247_adj_3956), 
            .CO(n22815));
    SB_LUT4 add_3392_3_lut (.I0(GND_net), .I1(n6761[0]), .I2(n174_adj_3958), 
            .I3(n22813), .O(n6745[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_3 (.CI(n22813), .I0(n6761[0]), .I1(n174_adj_3958), 
            .CO(n22814));
    SB_LUT4 add_3392_2_lut (.I0(GND_net), .I1(n32_adj_3959), .I2(n101_adj_3960), 
            .I3(GND_net), .O(n6745[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3392_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3392_2 (.CI(GND_net), .I0(n32_adj_3959), .I1(n101_adj_3960), 
            .CO(n22813));
    SB_LUT4 add_3391_16_lut (.I0(GND_net), .I1(n6745[13]), .I2(n1120_adj_3961), 
            .I3(n22812), .O(n6728[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3410_5_lut (.I0(GND_net), .I1(n6988[2]), .I2(n308), .I3(n22996), 
            .O(n6968[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3391_15_lut (.I0(GND_net), .I1(n6745[12]), .I2(n1047_adj_3962), 
            .I3(n22811), .O(n6728[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3410_5 (.CI(n22996), .I0(n6988[2]), .I1(n308), .CO(n22997));
    SB_CARRY add_3391_15 (.CI(n22811), .I0(n6745[12]), .I1(n1047_adj_3962), 
            .CO(n22812));
    SB_LUT4 add_3391_14_lut (.I0(GND_net), .I1(n6745[11]), .I2(n974_adj_3963), 
            .I3(n22810), .O(n6728[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24280_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n29370));   // verilog/motorControl.v(38[19:35])
    defparam i24280_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_3964));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3965));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3966));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3967));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3968));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3969));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3970));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3971));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_3972));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3391_14 (.CI(n22810), .I0(n6745[11]), .I1(n974_adj_3963), 
            .CO(n22811));
    SB_LUT4 add_3391_13_lut (.I0(GND_net), .I1(n6745[10]), .I2(n901_adj_3973), 
            .I3(n22809), .O(n6728[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_3974));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n22177), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_3976));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i22_3_lut (.I0(n155[21]), .I1(PWMLimit[21]), .I2(n256), 
            .I3(GND_net), .O(n2554[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3391_13 (.CI(n22809), .I0(n6745[10]), .I1(n901_adj_3973), 
            .CO(n22810));
    SB_LUT4 mux_561_i23_3_lut (.I0(n155[22]), .I1(PWMLimit[22]), .I2(n256), 
            .I3(GND_net), .O(n2554[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_561_i24_3_lut (.I0(n29296), .I1(PWMLimit[23]), .I2(n256), 
            .I3(GND_net), .O(n2554[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3391_12_lut (.I0(GND_net), .I1(n6745[9]), .I2(n828_adj_3977), 
            .I3(n22808), .O(n6728[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3978));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3979));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3980));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3981));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3982));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3983));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3984));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3410_4_lut (.I0(GND_net), .I1(n6988[1]), .I2(n235), .I3(n22995), 
            .O(n6968[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3985));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_3986));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_3987));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_3988));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_3989));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3410_4 (.CI(n22995), .I0(n6988[1]), .I1(n235), .CO(n22996));
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3990));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3991));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3992));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3391_12 (.CI(n22808), .I0(n6745[9]), .I1(n828_adj_3977), 
            .CO(n22809));
    SB_LUT4 add_3391_11_lut (.I0(GND_net), .I1(n6745[8]), .I2(n755_adj_3993), 
            .I3(n22807), .O(n6728[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_11 (.CI(n22807), .I0(n6745[8]), .I1(n755_adj_3993), 
            .CO(n22808));
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3994));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3995));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3996));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3997));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3998));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_3999));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4000));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4001));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4002));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n22177), .I0(GND_net), .I1(n1[16]), 
            .CO(n22178));
    SB_LUT4 add_3391_10_lut (.I0(GND_net), .I1(n6745[7]), .I2(n682_adj_4003), 
            .I3(n22806), .O(n6728[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_10 (.CI(n22806), .I0(n6745[7]), .I1(n682_adj_4003), 
            .CO(n22807));
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4004));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3391_9_lut (.I0(GND_net), .I1(n6745[6]), .I2(n609_adj_4005), 
            .I3(n22805), .O(n6728[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_9 (.CI(n22805), .I0(n6745[6]), .I1(n609_adj_4005), 
            .CO(n22806));
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4006));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3391_8_lut (.I0(GND_net), .I1(n6745[5]), .I2(n536_adj_4007), 
            .I3(n22804), .O(n6728[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3391_8 (.CI(n22804), .I0(n6745[5]), .I1(n536_adj_4007), 
            .CO(n22805));
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256), 
            .I3(GND_net), .O(n2554[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4008));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3391_7_lut (.I0(GND_net), .I1(n6745[4]), .I2(n463_adj_4009), 
            .I3(n22803), .O(n6728[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4010));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4011));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4012));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4013));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4014));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4015));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4017));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3410_3_lut (.I0(GND_net), .I1(n6988[0]), .I2(n162), .I3(n22994), 
            .O(n6968[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4019));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3410_3 (.CI(n22994), .I0(n6988[0]), .I1(n162), .CO(n22995));
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4020));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4021));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3391_7 (.CI(n22803), .I0(n6745[4]), .I1(n463_adj_4009), 
            .CO(n22804));
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4022));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4023));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4024));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3391_6_lut (.I0(GND_net), .I1(n6745[3]), .I2(n390_adj_4025), 
            .I3(n22802), .O(n6728[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4026));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4027));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4028));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4029));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3410_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n6968[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3410_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4030));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4032));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4033));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4034));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4035));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4037));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4039));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24270_4_lut (.I0(n21_adj_4037), .I1(n19_adj_4035), .I2(n17_adj_4034), 
            .I3(n9_adj_4033), .O(n29360));
    defparam i24270_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24264_4_lut (.I0(n27_adj_4032), .I1(n15_adj_4030), .I2(n13_adj_4029), 
            .I3(n11_adj_4028), .O(n29354));
    defparam i24264_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4039), 
            .I3(GND_net), .O(n12_adj_4040));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4029), 
            .I3(GND_net), .O(n10_adj_4041));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4040), .I1(n257[17]), .I2(n35_adj_4027), 
            .I3(GND_net), .O(n30_adj_4042));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24554_4_lut (.I0(n13_adj_4029), .I1(n11_adj_4028), .I2(n9_adj_4033), 
            .I3(n29370), .O(n29646));
    defparam i24554_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24550_4_lut (.I0(n19_adj_4035), .I1(n17_adj_4034), .I2(n15_adj_4030), 
            .I3(n29646), .O(n29642));
    defparam i24550_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24908_4_lut (.I0(n25_adj_4023), .I1(n23_adj_4022), .I2(n21_adj_4037), 
            .I3(n29642), .O(n30000));
    defparam i24908_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24743_4_lut (.I0(n31_adj_4026), .I1(n29_adj_4024), .I2(n27_adj_4032), 
            .I3(n30000), .O(n29835));
    defparam i24743_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24976_4_lut (.I0(n37_adj_4021), .I1(n35_adj_4027), .I2(n33_adj_4039), 
            .I3(n29835), .O(n30068));
    defparam i24976_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4020), 
            .I3(GND_net), .O(n16_adj_4043));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24894_3_lut (.I0(n6_adj_4044), .I1(n257[10]), .I2(n21_adj_4037), 
            .I3(GND_net), .O(n29986));   // verilog/motorControl.v(38[19:35])
    defparam i24894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24895_3_lut (.I0(n29986), .I1(n257[11]), .I2(n23_adj_4022), 
            .I3(GND_net), .O(n29987));   // verilog/motorControl.v(38[19:35])
    defparam i24895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4034), 
            .I3(GND_net), .O(n8_adj_4045));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4043), .I1(n257[22]), .I2(n45_adj_4019), 
            .I3(GND_net), .O(n24_adj_4046));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24250_4_lut (.I0(n43_adj_4020), .I1(n25_adj_4023), .I2(n23_adj_4022), 
            .I3(n29360), .O(n29340));
    defparam i24250_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24783_4_lut (.I0(n24_adj_4046), .I1(n8_adj_4045), .I2(n45_adj_4019), 
            .I3(n29338), .O(n29875));   // verilog/motorControl.v(38[19:35])
    defparam i24783_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24866_3_lut (.I0(n29987), .I1(n257[12]), .I2(n25_adj_4023), 
            .I3(GND_net), .O(n29958));   // verilog/motorControl.v(38[19:35])
    defparam i24866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n29248), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_4047));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24892_3_lut (.I0(n4_adj_4047), .I1(n257[13]), .I2(n27_adj_4032), 
            .I3(GND_net), .O(n29984));   // verilog/motorControl.v(38[19:35])
    defparam i24892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24893_3_lut (.I0(n29984), .I1(n257[14]), .I2(n29_adj_4024), 
            .I3(GND_net), .O(n29985));   // verilog/motorControl.v(38[19:35])
    defparam i24893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24260_4_lut (.I0(n33_adj_4039), .I1(n31_adj_4026), .I2(n29_adj_4024), 
            .I3(n29354), .O(n29350));
    defparam i24260_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24993_4_lut (.I0(n30_adj_4042), .I1(n10_adj_4041), .I2(n35_adj_4027), 
            .I3(n29348), .O(n30085));   // verilog/motorControl.v(38[19:35])
    defparam i24993_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24868_3_lut (.I0(n29985), .I1(n257[15]), .I2(n31_adj_4026), 
            .I3(GND_net), .O(n29960));   // verilog/motorControl.v(38[19:35])
    defparam i24868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25039_4_lut (.I0(n29960), .I1(n30085), .I2(n35_adj_4027), 
            .I3(n29350), .O(n30131));   // verilog/motorControl.v(38[19:35])
    defparam i25039_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25040_3_lut (.I0(n30131), .I1(n257[18]), .I2(n37_adj_4021), 
            .I3(GND_net), .O(n30132));   // verilog/motorControl.v(38[19:35])
    defparam i25040_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3410_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n22994));
    SB_LUT4 i25016_3_lut (.I0(n30132), .I1(n257[19]), .I2(n39_adj_4017), 
            .I3(GND_net), .O(n30108));   // verilog/motorControl.v(38[19:35])
    defparam i25016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24252_4_lut (.I0(n43_adj_4020), .I1(n41_adj_4015), .I2(n39_adj_4017), 
            .I3(n30068), .O(n29342));
    defparam i24252_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3409_20_lut (.I0(GND_net), .I1(n6968[17]), .I2(GND_net), 
            .I3(n22993), .O(n6947[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24946_4_lut (.I0(n29958), .I1(n29875), .I2(n45_adj_4019), 
            .I3(n29340), .O(n30038));   // verilog/motorControl.v(38[19:35])
    defparam i24946_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3409_19_lut (.I0(GND_net), .I1(n6968[16]), .I2(GND_net), 
            .I3(n22992), .O(n6947[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_19 (.CI(n22992), .I0(n6968[16]), .I1(GND_net), .CO(n22993));
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_4044));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_3409_18_lut (.I0(GND_net), .I1(n6968[15]), .I2(GND_net), 
            .I3(n22991), .O(n6947[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25010_3_lut (.I0(n30108), .I1(n257[20]), .I2(n41_adj_4015), 
            .I3(GND_net), .O(n40_adj_4048));   // verilog/motorControl.v(38[19:35])
    defparam i25010_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3409_18 (.CI(n22991), .I0(n6968[15]), .I1(GND_net), .CO(n22992));
    SB_LUT4 add_3409_17_lut (.I0(GND_net), .I1(n6968[14]), .I2(GND_net), 
            .I3(n22990), .O(n6947[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_17 (.CI(n22990), .I0(n6968[14]), .I1(GND_net), .CO(n22991));
    SB_LUT4 add_3409_16_lut (.I0(GND_net), .I1(n6968[13]), .I2(n1108), 
            .I3(n22989), .O(n6947[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_16 (.CI(n22989), .I0(n6968[13]), .I1(n1108), .CO(n22990));
    SB_LUT4 add_3409_15_lut (.I0(GND_net), .I1(n6968[12]), .I2(n1035), 
            .I3(n22988), .O(n6947[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_6 (.CI(n22802), .I0(n6745[3]), .I1(n390_adj_4025), 
            .CO(n22803));
    SB_CARRY add_3409_15 (.CI(n22988), .I0(n6968[12]), .I1(n1035), .CO(n22989));
    SB_LUT4 add_3409_14_lut (.I0(GND_net), .I1(n6968[11]), .I2(n962), 
            .I3(n22987), .O(n6947[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24948_4_lut (.I0(n40_adj_4048), .I1(n30038), .I2(n45_adj_4019), 
            .I3(n29342), .O(n30040));   // verilog/motorControl.v(38[19:35])
    defparam i24948_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3409_14 (.CI(n22987), .I0(n6968[11]), .I1(n962), .CO(n22988));
    SB_LUT4 i24949_3_lut (.I0(n30040), .I1(duty[23]), .I2(n47_adj_4049), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i24949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3409_13_lut (.I0(GND_net), .I1(n6968[10]), .I2(n889), 
            .I3(n22986), .O(n6947[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_13 (.CI(n22986), .I0(n6968[10]), .I1(n889), .CO(n22987));
    SB_LUT4 i14854_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n18679));   // verilog/motorControl.v(38[19:35])
    defparam i14854_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3409_12_lut (.I0(GND_net), .I1(n6968[9]), .I2(n816), .I3(n22985), 
            .O(n6947[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_12 (.CI(n22985), .I0(n6968[9]), .I1(n816), .CO(n22986));
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4050));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3409_11_lut (.I0(GND_net), .I1(n6968[8]), .I2(n743), .I3(n22984), 
            .O(n6947[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_11 (.CI(n22984), .I0(n6968[8]), .I1(n743), .CO(n22985));
    SB_LUT4 add_3409_10_lut (.I0(GND_net), .I1(n6968[7]), .I2(n670), .I3(n22983), 
            .O(n6947[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_10 (.CI(n22983), .I0(n6968[7]), .I1(n670), .CO(n22984));
    SB_LUT4 add_3391_5_lut (.I0(GND_net), .I1(n6745[2]), .I2(n317_adj_4051), 
            .I3(n22801), .O(n6728[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_5 (.CI(n22801), .I0(n6745[2]), .I1(n317_adj_4051), 
            .CO(n22802));
    SB_LUT4 add_3409_9_lut (.I0(GND_net), .I1(n6968[6]), .I2(n597), .I3(n22982), 
            .O(n6947[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3391_4_lut (.I0(GND_net), .I1(n6745[1]), .I2(n244_adj_4052), 
            .I3(n22800), .O(n6728[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_4 (.CI(n22800), .I0(n6745[1]), .I1(n244_adj_4052), 
            .CO(n22801));
    SB_CARRY add_3409_9 (.CI(n22982), .I0(n6968[6]), .I1(n597), .CO(n22983));
    SB_LUT4 add_3409_8_lut (.I0(GND_net), .I1(n6968[5]), .I2(n524), .I3(n22981), 
            .O(n6947[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_8 (.CI(n22981), .I0(n6968[5]), .I1(n524), .CO(n22982));
    SB_LUT4 add_3409_7_lut (.I0(GND_net), .I1(n6968[4]), .I2(n451), .I3(n22980), 
            .O(n6947[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3391_3_lut (.I0(GND_net), .I1(n6745[0]), .I2(n171_adj_4053), 
            .I3(n22799), .O(n6728[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4054));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3409_7 (.CI(n22980), .I0(n6968[4]), .I1(n451), .CO(n22981));
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4055));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3409_6_lut (.I0(GND_net), .I1(n6968[3]), .I2(n378), .I3(n22979), 
            .O(n6947[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_6 (.CI(n22979), .I0(n6968[3]), .I1(n378), .CO(n22980));
    SB_LUT4 add_3409_5_lut (.I0(GND_net), .I1(n6968[2]), .I2(n305), .I3(n22978), 
            .O(n6947[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3409_5 (.CI(n22978), .I0(n6968[2]), .I1(n305), .CO(n22979));
    SB_LUT4 add_3409_4_lut (.I0(GND_net), .I1(n6968[1]), .I2(n232), .I3(n22977), 
            .O(n6947[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3391_3 (.CI(n22799), .I0(n6745[0]), .I1(n171_adj_4053), 
            .CO(n22800));
    SB_LUT4 add_3391_2_lut (.I0(GND_net), .I1(n29_adj_4056), .I2(n98_adj_4057), 
            .I3(GND_net), .O(n6728[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3391_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3391_2 (.CI(GND_net), .I0(n29_adj_4056), .I1(n98_adj_4057), 
            .CO(n22799));
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4058));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3409_4 (.CI(n22977), .I0(n6968[1]), .I1(n232), .CO(n22978));
    SB_LUT4 add_3409_3_lut (.I0(GND_net), .I1(n6968[0]), .I2(n159), .I3(n22976), 
            .O(n6947[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4059));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_17_lut (.I0(GND_net), .I1(n6728[14]), .I2(GND_net), 
            .I3(n22798), .O(n6710[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4060));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3409_3 (.CI(n22976), .I0(n6968[0]), .I1(n159), .CO(n22977));
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4061));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4062));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3409_2_lut (.I0(GND_net), .I1(n17_adj_4063), .I2(n86), 
            .I3(GND_net), .O(n6947[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3409_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4064));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4065));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4066));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3390_16_lut (.I0(GND_net), .I1(n6728[13]), .I2(n1117_adj_4068), 
            .I3(n22797), .O(n6710[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_16 (.CI(n22797), .I0(n6728[13]), .I1(n1117_adj_4068), 
            .CO(n22798));
    SB_LUT4 add_3390_15_lut (.I0(GND_net), .I1(n6728[12]), .I2(n1044_adj_4069), 
            .I3(n22796), .O(n6710[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_15 (.CI(n22796), .I0(n6728[12]), .I1(n1044_adj_4069), 
            .CO(n22797));
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4070));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4071));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4072));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_14_lut (.I0(GND_net), .I1(n6728[11]), .I2(n971_adj_4073), 
            .I3(n22795), .O(n6710[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_14 (.CI(n22795), .I0(n6728[11]), .I1(n971_adj_4073), 
            .CO(n22796));
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4074));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4075));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4076));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_13_lut (.I0(GND_net), .I1(n6728[10]), .I2(n898_adj_4077), 
            .I3(n22794), .O(n6710[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4078));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4079));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4080), .I1(\Kp[4] ), .I2(n6860[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n6853[3]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3390_13 (.CI(n22794), .I0(n6728[10]), .I1(n898_adj_4077), 
            .CO(n22795));
    SB_LUT4 add_3390_12_lut (.I0(GND_net), .I1(n6728[9]), .I2(n825_adj_4082), 
            .I3(n22793), .O(n6710[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n22176), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17932_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n6871[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17932_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3390_12 (.CI(n22793), .I0(n6728[9]), .I1(n825_adj_4082), 
            .CO(n22794));
    SB_LUT4 add_3390_11_lut (.I0(GND_net), .I1(n6728[8]), .I2(n752_adj_4084), 
            .I3(n22792), .O(n6710[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_3961));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1462 (.I0(n4_adj_4085), .I1(\Kp[3] ), .I2(n6866[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6860[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1462.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4086));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1463 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12_adj_4087));   // verilog/motorControl.v(34[17:23])
    defparam i2_4_lut_adj_1463.LUT_INIT = 16'h9c50;
    SB_LUT4 i17868_4_lut (.I0(n6860[2]), .I1(\Kp[4] ), .I2(n6_adj_4080), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_4088));   // verilog/motorControl.v(34[17:23])
    defparam i17868_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_4089));   // verilog/motorControl.v(34[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i17899_4_lut (.I0(n6866[1]), .I1(\Kp[3] ), .I2(n4_adj_4085), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_4090));   // verilog/motorControl.v(34[17:23])
    defparam i17899_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17934_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n21745));   // verilog/motorControl.v(34[17:23])
    defparam i17934_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n21745), .I3(n4_adj_4091), 
            .O(n27329));   // verilog/motorControl.v(34[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3409_2 (.CI(GND_net), .I0(n17_adj_4063), .I1(n86), .CO(n22976));
    SB_LUT4 mux_561_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256), 
            .I3(GND_net), .O(n2554[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4092));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3408_21_lut (.I0(GND_net), .I1(n6947[18]), .I2(GND_net), 
            .I3(n22975), .O(n6925[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4093));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4094));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3960));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3959));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4095));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_3958));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4096));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_3956));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4097));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_3955));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4098));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3390_11 (.CI(n22792), .I0(n6728[8]), .I1(n752_adj_4084), 
            .CO(n22793));
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3408_20_lut (.I0(GND_net), .I1(n6947[17]), .I2(GND_net), 
            .I3(n22974), .O(n6925[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3390_10_lut (.I0(GND_net), .I1(n6728[7]), .I2(n679_adj_4099), 
            .I3(n22791), .O(n6710[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_10 (.CI(n22791), .I0(n6728[7]), .I1(n679_adj_4099), 
            .CO(n22792));
    SB_LUT4 add_3390_9_lut (.I0(GND_net), .I1(n6728[6]), .I2(n606_adj_4100), 
            .I3(n22790), .O(n6710[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3408_20 (.CI(n22974), .I0(n6947[17]), .I1(GND_net), .CO(n22975));
    SB_CARRY add_3390_9 (.CI(n22790), .I0(n6728[6]), .I1(n606_adj_4100), 
            .CO(n22791));
    SB_LUT4 add_3408_19_lut (.I0(GND_net), .I1(n6947[16]), .I2(GND_net), 
            .I3(n22973), .O(n6925[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_19 (.CI(n22973), .I0(n6947[16]), .I1(GND_net), .CO(n22974));
    SB_LUT4 add_3408_18_lut (.I0(GND_net), .I1(n6947[15]), .I2(GND_net), 
            .I3(n22972), .O(n6925[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3408_18 (.CI(n22972), .I0(n6947[15]), .I1(GND_net), .CO(n22973));
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4102));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4103));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3408_17_lut (.I0(GND_net), .I1(n6947[14]), .I2(GND_net), 
            .I3(n22971), .O(n6925[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_17 (.CI(n22971), .I0(n6947[14]), .I1(GND_net), .CO(n22972));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n22176), .I0(GND_net), .I1(n1[15]), 
            .CO(n22177));
    SB_LUT4 add_3408_16_lut (.I0(GND_net), .I1(n6947[13]), .I2(n1105), 
            .I3(n22970), .O(n6925[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3390_8_lut (.I0(GND_net), .I1(n6728[5]), .I2(n533_adj_4104), 
            .I3(n22789), .O(n6710[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_16 (.CI(n22970), .I0(n6947[13]), .I1(n1105), .CO(n22971));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n22175), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3390_8 (.CI(n22789), .I0(n6728[5]), .I1(n533_adj_4104), 
            .CO(n22790));
    SB_LUT4 add_3390_7_lut (.I0(GND_net), .I1(n6728[4]), .I2(n460_adj_4106), 
            .I3(n22788), .O(n6710[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_7 (.CI(n22788), .I0(n6728[4]), .I1(n460_adj_4106), 
            .CO(n22789));
    SB_LUT4 add_3390_6_lut (.I0(GND_net), .I1(n6728[3]), .I2(n387_adj_4107), 
            .I3(n22787), .O(n6710[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3368[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_3390_6 (.CI(n22787), .I0(n6728[3]), .I1(n387_adj_4107), 
            .CO(n22788));
    SB_LUT4 add_3390_5_lut (.I0(GND_net), .I1(n6728[2]), .I2(n314_adj_4108), 
            .I3(n22786), .O(n6710[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3408_15_lut (.I0(GND_net), .I1(n6947[12]), .I2(n1032), 
            .I3(n22969), .O(n6925[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n22175), .I0(GND_net), .I1(n1[14]), 
            .CO(n22176));
    SB_CARRY add_3390_5 (.CI(n22786), .I0(n6728[2]), .I1(n314_adj_4108), 
            .CO(n22787));
    SB_CARRY add_3408_15 (.CI(n22969), .I0(n6947[12]), .I1(n1032), .CO(n22970));
    SB_LUT4 add_3390_4_lut (.I0(GND_net), .I1(n6728[1]), .I2(n241_adj_4109), 
            .I3(n22785), .O(n6710[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_3954));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_3953));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3390_4 (.CI(n22785), .I0(n6728[1]), .I1(n241_adj_4109), 
            .CO(n22786));
    SB_LUT4 add_3390_3_lut (.I0(GND_net), .I1(n6728[0]), .I2(n168_adj_4110), 
            .I3(n22784), .O(n6710[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3390_3 (.CI(n22784), .I0(n6728[0]), .I1(n168_adj_4110), 
            .CO(n22785));
    SB_LUT4 add_3408_14_lut (.I0(GND_net), .I1(n6947[11]), .I2(n959), 
            .I3(n22968), .O(n6925[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3390_2_lut (.I0(GND_net), .I1(n26_adj_4111), .I2(n95_adj_4112), 
            .I3(GND_net), .O(n6710[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3390_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3938));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3390_2 (.CI(GND_net), .I0(n26_adj_4111), .I1(n95_adj_4112), 
            .CO(n22784));
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3389_18_lut (.I0(GND_net), .I1(n6710[15]), .I2(GND_net), 
            .I3(n22783), .O(n6691[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_14 (.CI(n22968), .I0(n6947[11]), .I1(n959), .CO(n22969));
    SB_LUT4 add_3408_13_lut (.I0(GND_net), .I1(n6947[10]), .I2(n886), 
            .I3(n22967), .O(n6925[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_17_lut (.I0(GND_net), .I1(n6710[14]), .I2(GND_net), 
            .I3(n22782), .O(n6691[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_13 (.CI(n22967), .I0(n6947[10]), .I1(n886), .CO(n22968));
    SB_LUT4 add_3408_12_lut (.I0(GND_net), .I1(n6947[9]), .I2(n813), .I3(n22966), 
            .O(n6925[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_17 (.CI(n22782), .I0(n6710[14]), .I1(GND_net), .CO(n22783));
    SB_CARRY add_3408_12 (.CI(n22966), .I0(n6947[9]), .I1(n813), .CO(n22967));
    SB_LUT4 add_3408_11_lut (.I0(GND_net), .I1(n6947[8]), .I2(n740), .I3(n22965), 
            .O(n6925[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_16_lut (.I0(GND_net), .I1(n6710[13]), .I2(n1114_adj_4113), 
            .I3(n22781), .O(n6691[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_11 (.CI(n22965), .I0(n6947[8]), .I1(n740), .CO(n22966));
    SB_LUT4 add_3408_10_lut (.I0(GND_net), .I1(n6947[7]), .I2(n667), .I3(n22964), 
            .O(n6925[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_10 (.CI(n22964), .I0(n6947[7]), .I1(n667), .CO(n22965));
    SB_LUT4 add_3408_9_lut (.I0(GND_net), .I1(n6947[6]), .I2(n594), .I3(n22963), 
            .O(n6925[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_9 (.CI(n22963), .I0(n6947[6]), .I1(n594), .CO(n22964));
    SB_CARRY add_3389_16 (.CI(n22781), .I0(n6710[13]), .I1(n1114_adj_4113), 
            .CO(n22782));
    SB_LUT4 add_3408_8_lut (.I0(GND_net), .I1(n6947[5]), .I2(n521), .I3(n22962), 
            .O(n6925[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_15_lut (.I0(GND_net), .I1(n6710[12]), .I2(n1041_adj_4114), 
            .I3(n22780), .O(n6691[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_8 (.CI(n22962), .I0(n6947[5]), .I1(n521), .CO(n22963));
    SB_LUT4 add_3408_7_lut (.I0(GND_net), .I1(n6947[4]), .I2(n448), .I3(n22961), 
            .O(n6925[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_15 (.CI(n22780), .I0(n6710[12]), .I1(n1041_adj_4114), 
            .CO(n22781));
    SB_CARRY add_3408_7 (.CI(n22961), .I0(n6947[4]), .I1(n448), .CO(n22962));
    SB_LUT4 add_3408_6_lut (.I0(GND_net), .I1(n6947[3]), .I2(n375), .I3(n22960), 
            .O(n6925[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_6 (.CI(n22960), .I0(n6947[3]), .I1(n375), .CO(n22961));
    SB_LUT4 add_3408_5_lut (.I0(GND_net), .I1(n6947[2]), .I2(n302), .I3(n22959), 
            .O(n6925[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_5 (.CI(n22959), .I0(n6947[2]), .I1(n302), .CO(n22960));
    SB_LUT4 add_3389_14_lut (.I0(GND_net), .I1(n6710[11]), .I2(n968_adj_4115), 
            .I3(n22779), .O(n6691[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3408_4_lut (.I0(GND_net), .I1(n6947[1]), .I2(n229), .I3(n22958), 
            .O(n6925[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_4 (.CI(n22958), .I0(n6947[1]), .I1(n229), .CO(n22959));
    SB_LUT4 add_3408_3_lut (.I0(GND_net), .I1(n6947[0]), .I2(n156), .I3(n22957), 
            .O(n6925[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3408_3 (.CI(n22957), .I0(n6947[0]), .I1(n156), .CO(n22958));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n22174), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3408_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n6925[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3408_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n22174), .I0(GND_net), .I1(n1[13]), 
            .CO(n22175));
    SB_CARRY add_3408_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n22957));
    SB_LUT4 add_3407_22_lut (.I0(GND_net), .I1(n6925[19]), .I2(GND_net), 
            .I3(n22956), .O(n6902[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_14 (.CI(n22779), .I0(n6710[11]), .I1(n968_adj_4115), 
            .CO(n22780));
    SB_LUT4 mux_561_i18_3_lut (.I0(n155[17]), .I1(PWMLimit[17]), .I2(n256), 
            .I3(GND_net), .O(n2554[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_3952));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_21_lut (.I0(GND_net), .I1(n6925[18]), .I2(GND_net), 
            .I3(n22955), .O(n6902[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_21 (.CI(n22955), .I0(n6925[18]), .I1(GND_net), .CO(n22956));
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_3951));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_20_lut (.I0(GND_net), .I1(n6925[17]), .I2(GND_net), 
            .I3(n22954), .O(n6902[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_20 (.CI(n22954), .I0(n6925[17]), .I1(GND_net), .CO(n22955));
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_3950));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_3949));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3389_13_lut (.I0(GND_net), .I1(n6710[10]), .I2(n895_adj_4118), 
            .I3(n22778), .O(n6691[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_19_lut (.I0(GND_net), .I1(n6925[16]), .I2(GND_net), 
            .I3(n22953), .O(n6902[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n22173), .O(n25_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_13 (.CI(n22778), .I0(n6710[10]), .I1(n895_adj_4118), 
            .CO(n22779));
    SB_LUT4 add_3389_12_lut (.I0(GND_net), .I1(n6710[9]), .I2(n822_adj_4120), 
            .I3(n22777), .O(n6691[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_3948));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_19 (.CI(n22953), .I0(n6925[16]), .I1(GND_net), .CO(n22954));
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_18_lut (.I0(GND_net), .I1(n6925[15]), .I2(GND_net), 
            .I3(n22952), .O(n6902[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_18 (.CI(n22952), .I0(n6925[15]), .I1(GND_net), .CO(n22953));
    SB_LUT4 add_3407_17_lut (.I0(GND_net), .I1(n6925[14]), .I2(GND_net), 
            .I3(n22951), .O(n6902[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_17 (.CI(n22951), .I0(n6925[14]), .I1(GND_net), .CO(n22952));
    SB_CARRY unary_minus_5_add_3_14 (.CI(n22173), .I0(GND_net), .I1(n1[12]), 
            .CO(n22174));
    SB_LUT4 add_3407_16_lut (.I0(GND_net), .I1(n6925[13]), .I2(n1102), 
            .I3(n22950), .O(n6902[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_12 (.CI(n22777), .I0(n6710[9]), .I1(n822_adj_4120), 
            .CO(n22778));
    SB_CARRY add_3407_16 (.CI(n22950), .I0(n6925[13]), .I1(n1102), .CO(n22951));
    SB_LUT4 add_3407_15_lut (.I0(GND_net), .I1(n6925[12]), .I2(n1029), 
            .I3(n22949), .O(n6902[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_3947));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n22172), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4122));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3389_11_lut (.I0(GND_net), .I1(n6710[8]), .I2(n749_adj_4123), 
            .I3(n22776), .O(n6691[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4124));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n22172), .I0(GND_net), .I1(n1[11]), 
            .CO(n22173));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n22171), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4126));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_11 (.CI(n22776), .I0(n6710[8]), .I1(n749_adj_4123), 
            .CO(n22777));
    SB_CARRY add_3407_15 (.CI(n22949), .I0(n6925[12]), .I1(n1029), .CO(n22950));
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4127));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_14_lut (.I0(GND_net), .I1(n6925[11]), .I2(n956_adj_4128), 
            .I3(n22948), .O(n6902[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_10_lut (.I0(GND_net), .I1(n6710[7]), .I2(n676_adj_4129), 
            .I3(n22775), .O(n6691[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n22171), .I0(GND_net), .I1(n1[10]), 
            .CO(n22172));
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_3946));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4130));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_10 (.CI(n22775), .I0(n6710[7]), .I1(n676_adj_4129), 
            .CO(n22776));
    SB_LUT4 add_3389_9_lut (.I0(GND_net), .I1(n6710[6]), .I2(n603_adj_4131), 
            .I3(n22774), .O(n6691[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_9 (.CI(n22774), .I0(n6710[6]), .I1(n603_adj_4131), 
            .CO(n22775));
    SB_LUT4 add_3389_8_lut (.I0(GND_net), .I1(n6710[5]), .I2(n530_adj_4132), 
            .I3(n22773), .O(n6691[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_8 (.CI(n22773), .I0(n6710[5]), .I1(n530_adj_4132), 
            .CO(n22774));
    SB_LUT4 add_3389_7_lut (.I0(GND_net), .I1(n6710[4]), .I2(n457_adj_4133), 
            .I3(n22772), .O(n6691[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_7 (.CI(n22772), .I0(n6710[4]), .I1(n457_adj_4133), 
            .CO(n22773));
    SB_LUT4 add_3389_6_lut (.I0(GND_net), .I1(n6710[3]), .I2(n384_adj_4134), 
            .I3(n22771), .O(n6691[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4135));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_3945));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_6 (.CI(n22771), .I0(n6710[3]), .I1(n384_adj_4134), 
            .CO(n22772));
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n22170), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3389_5_lut (.I0(GND_net), .I1(n6710[2]), .I2(n311_adj_4137), 
            .I3(n22770), .O(n6691[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_5 (.CI(n22770), .I0(n6710[2]), .I1(n311_adj_4137), 
            .CO(n22771));
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3389_4_lut (.I0(GND_net), .I1(n6710[1]), .I2(n238_adj_4138), 
            .I3(n22769), .O(n6691[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4139));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3944));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4140));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3943));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_4 (.CI(n22769), .I0(n6710[1]), .I1(n238_adj_4138), 
            .CO(n22770));
    SB_LUT4 add_3389_3_lut (.I0(GND_net), .I1(n6710[0]), .I2(n165_adj_4141), 
            .I3(n22768), .O(n6691[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_3 (.CI(n22768), .I0(n6710[0]), .I1(n165_adj_4141), 
            .CO(n22769));
    SB_LUT4 add_3389_2_lut (.I0(GND_net), .I1(n23_adj_4142), .I2(n92_adj_4143), 
            .I3(GND_net), .O(n6691[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_2 (.CI(GND_net), .I0(n23_adj_4142), .I1(n92_adj_4143), 
            .CO(n22768));
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4144));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_19_lut (.I0(GND_net), .I1(n6691[16]), .I2(GND_net), 
            .I3(n22767), .O(n6671[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3388_18_lut (.I0(GND_net), .I1(n6691[15]), .I2(GND_net), 
            .I3(n22766), .O(n6671[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_18 (.CI(n22766), .I0(n6691[15]), .I1(GND_net), .CO(n22767));
    SB_CARRY add_3407_14 (.CI(n22948), .I0(n6925[11]), .I1(n956_adj_4128), 
            .CO(n22949));
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_17_lut (.I0(GND_net), .I1(n6691[14]), .I2(GND_net), 
            .I3(n22765), .O(n6671[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_13_lut (.I0(GND_net), .I1(n6925[10]), .I2(n883_adj_4145), 
            .I3(n22947), .O(n6902[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_3942));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_17 (.CI(n22765), .I0(n6691[14]), .I1(GND_net), .CO(n22766));
    SB_LUT4 add_3388_16_lut (.I0(GND_net), .I1(n6691[13]), .I2(n1111_adj_4146), 
            .I3(n22764), .O(n6671[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4147));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4148));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_3941));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4149));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4150));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4151));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4152));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4153));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4154));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4155));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4156));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4157));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4158));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4090), .I1(n11_adj_4089), .I2(n8_adj_4088), 
            .I3(n12_adj_4087), .O(n18));   // verilog/motorControl.v(34[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4159));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4160));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4161));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_13 (.CI(n22947), .I0(n6925[10]), .I1(n883_adj_4145), 
            .CO(n22948));
    SB_LUT4 add_3407_12_lut (.I0(GND_net), .I1(n6925[9]), .I2(n810_adj_4162), 
            .I3(n22946), .O(n6902[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_12 (.CI(n22946), .I0(n6925[9]), .I1(n810_adj_4162), 
            .CO(n22947));
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4163));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_11_lut (.I0(GND_net), .I1(n6925[8]), .I2(n737_adj_4164), 
            .I3(n22945), .O(n6902[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_11 (.CI(n22945), .I0(n6925[8]), .I1(n737_adj_4164), 
            .CO(n22946));
    SB_LUT4 add_3407_10_lut (.I0(GND_net), .I1(n6925[7]), .I2(n664_adj_4165), 
            .I3(n22944), .O(n6902[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4166));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_10 (.CI(n22944), .I0(n6925[7]), .I1(n664_adj_4165), 
            .CO(n22945));
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4167));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_9_lut (.I0(GND_net), .I1(n6925[6]), .I2(n591_adj_4168), 
            .I3(n22943), .O(n6902[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_9 (.CI(n22943), .I0(n6925[6]), .I1(n591_adj_4168), 
            .CO(n22944));
    SB_LUT4 add_3407_8_lut (.I0(GND_net), .I1(n6925[5]), .I2(n518_adj_4169), 
            .I3(n22942), .O(n6902[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_8 (.CI(n22942), .I0(n6925[5]), .I1(n518_adj_4169), 
            .CO(n22943));
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4170));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_7_lut (.I0(GND_net), .I1(n6925[4]), .I2(n445_adj_4171), 
            .I3(n22941), .O(n6902[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_7 (.CI(n22941), .I0(n6925[4]), .I1(n445_adj_4171), 
            .CO(n22942));
    SB_LUT4 add_3407_6_lut (.I0(GND_net), .I1(n6925[3]), .I2(n372_adj_4172), 
            .I3(n22940), .O(n6902[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_16 (.CI(n22764), .I0(n6691[13]), .I1(n1111_adj_4146), 
            .CO(n22765));
    SB_LUT4 add_3388_15_lut (.I0(GND_net), .I1(n6691[12]), .I2(n1038_adj_4173), 
            .I3(n22763), .O(n6671[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_6 (.CI(n22940), .I0(n6925[3]), .I1(n372_adj_4172), 
            .CO(n22941));
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4174));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4175));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_15 (.CI(n22763), .I0(n6691[12]), .I1(n1038_adj_4173), 
            .CO(n22764));
    SB_LUT4 add_3388_14_lut (.I0(GND_net), .I1(n6691[11]), .I2(n965_adj_4176), 
            .I3(n22762), .O(n6671[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_5_lut (.I0(GND_net), .I1(n6925[2]), .I2(n299_adj_4177), 
            .I3(n22939), .O(n6902[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n22170), .I0(GND_net), .I1(n1[9]), 
            .CO(n22171));
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4179));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4180));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_14 (.CI(n22762), .I0(n6691[11]), .I1(n965_adj_4176), 
            .CO(n22763));
    SB_LUT4 add_3388_13_lut (.I0(GND_net), .I1(n6691[10]), .I2(n892_adj_4181), 
            .I3(n22761), .O(n6671[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_13 (.CI(n22761), .I0(n6691[10]), .I1(n892_adj_4181), 
            .CO(n22762));
    SB_LUT4 add_3388_12_lut (.I0(GND_net), .I1(n6691[9]), .I2(n819_adj_4182), 
            .I3(n22760), .O(n6671[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_12 (.CI(n22760), .I0(n6691[9]), .I1(n819_adj_4182), 
            .CO(n22761));
    SB_LUT4 add_3388_11_lut (.I0(GND_net), .I1(n6691[8]), .I2(n746_adj_4183), 
            .I3(n22759), .O(n6671[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_5 (.CI(n22939), .I0(n6925[2]), .I1(n299_adj_4177), 
            .CO(n22940));
    SB_CARRY add_3388_11 (.CI(n22759), .I0(n6691[8]), .I1(n746_adj_4183), 
            .CO(n22760));
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4184));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_4_lut (.I0(GND_net), .I1(n6925[1]), .I2(n226_adj_4185), 
            .I3(n22938), .O(n6902[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_4 (.CI(n22938), .I0(n6925[1]), .I1(n226_adj_4185), 
            .CO(n22939));
    SB_LUT4 add_3407_3_lut (.I0(GND_net), .I1(n6925[0]), .I2(n153_adj_4186), 
            .I3(n22937), .O(n6902[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_3 (.CI(n22937), .I0(n6925[0]), .I1(n153_adj_4186), 
            .CO(n22938));
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4187));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n22169), .O(n17_adj_3906)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3388_10_lut (.I0(GND_net), .I1(n6691[7]), .I2(n673_adj_4189), 
            .I3(n22758), .O(n6671[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_2_lut (.I0(GND_net), .I1(n11_adj_4190), .I2(n80_adj_4191), 
            .I3(GND_net), .O(n6902[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_10 (.CI(n22758), .I0(n6691[7]), .I1(n673_adj_4189), 
            .CO(n22759));
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4192));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n22169), .I0(GND_net), .I1(n1[8]), 
            .CO(n22170));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n22168), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3407_2 (.CI(GND_net), .I0(n11_adj_4190), .I1(n80_adj_4191), 
            .CO(n22937));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n6878[21]), 
            .I2(GND_net), .I3(n22936), .O(n29296)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4194));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4195));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n6878[20]), .I2(GND_net), 
            .I3(n22935), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n22935), .I0(n6878[20]), .I1(GND_net), 
            .CO(n22936));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n6878[19]), .I2(GND_net), 
            .I3(n22934), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n22168), .I0(GND_net), .I1(n1[7]), 
            .CO(n22169));
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4196));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_9_lut (.I0(GND_net), .I1(n6691[6]), .I2(n600_adj_4197), 
            .I3(n22757), .O(n6671[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_9 (.CI(n22757), .I0(n6691[6]), .I1(n600_adj_4197), 
            .CO(n22758));
    SB_LUT4 add_3388_8_lut (.I0(GND_net), .I1(n6691[5]), .I2(n527_adj_4198), 
            .I3(n22756), .O(n6671[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_8 (.CI(n22756), .I0(n6691[5]), .I1(n527_adj_4198), 
            .CO(n22757));
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4199));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_7_lut (.I0(GND_net), .I1(n6691[4]), .I2(n454_adj_4200), 
            .I3(n22755), .O(n6671[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4201));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n22167), .O(n13_adj_3904)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4203));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_22 (.CI(n22934), .I0(n6878[19]), .I1(GND_net), 
            .CO(n22935));
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4205));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_7 (.CI(n22755), .I0(n6691[4]), .I1(n454_adj_4200), 
            .CO(n22756));
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4206));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4207));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4208));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_6_lut (.I0(GND_net), .I1(n6691[3]), .I2(n381_adj_4209), 
            .I3(n22754), .O(n6671[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4210));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n6878[18]), .I2(GND_net), 
            .I3(n22933), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n22933), .I0(n6878[18]), .I1(GND_net), 
            .CO(n22934));
    SB_CARRY add_3388_6 (.CI(n22754), .I0(n6691[3]), .I1(n381_adj_4209), 
            .CO(n22755));
    SB_LUT4 add_3388_5_lut (.I0(GND_net), .I1(n6691[2]), .I2(n308_adj_4211), 
            .I3(n22753), .O(n6671[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n6878[17]), .I2(GND_net), 
            .I3(n22932), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3388_5 (.CI(n22753), .I0(n6691[2]), .I1(n308_adj_4211), 
            .CO(n22754));
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3388_4_lut (.I0(GND_net), .I1(n6691[1]), .I2(n235_adj_4212), 
            .I3(n22752), .O(n6671[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_4 (.CI(n22752), .I0(n6691[1]), .I1(n235_adj_4212), 
            .CO(n22753));
    SB_LUT4 add_3388_3_lut (.I0(GND_net), .I1(n6691[0]), .I2(n162_adj_4213), 
            .I3(n22751), .O(n6671[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_3 (.CI(n22751), .I0(n6691[0]), .I1(n162_adj_4213), 
            .CO(n22752));
    SB_LUT4 add_3388_2_lut (.I0(GND_net), .I1(n20_adj_4214), .I2(n89_adj_4215), 
            .I3(GND_net), .O(n6671[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3388_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3388_2 (.CI(GND_net), .I0(n20_adj_4214), .I1(n89_adj_4215), 
            .CO(n22751));
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4216));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3387_20_lut (.I0(GND_net), .I1(n6671[17]), .I2(GND_net), 
            .I3(n22750), .O(n6650[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4217));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3387_19_lut (.I0(GND_net), .I1(n6671[16]), .I2(GND_net), 
            .I3(n22749), .O(n6650[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4218));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_20 (.CI(n22932), .I0(n6878[17]), .I1(GND_net), 
            .CO(n22933));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4219));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_19 (.CI(n22749), .I0(n6671[16]), .I1(GND_net), .CO(n22750));
    SB_LUT4 add_3387_18_lut (.I0(GND_net), .I1(n6671[15]), .I2(GND_net), 
            .I3(n22748), .O(n6650[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4220));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4221));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4222));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4223));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n6878[16]), .I2(GND_net), 
            .I3(n22931), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4224));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4225));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4226));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4215));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_18 (.CI(n22748), .I0(n6671[15]), .I1(GND_net), .CO(n22749));
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4214));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3387_17_lut (.I0(GND_net), .I1(n6671[14]), .I2(GND_net), 
            .I3(n22747), .O(n6650[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4213));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3940));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4212));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_17 (.CI(n22747), .I0(n6671[14]), .I1(GND_net), .CO(n22748));
    SB_LUT4 add_3387_16_lut (.I0(GND_net), .I1(n6671[13]), .I2(n1108_adj_4226), 
            .I3(n22746), .O(n6650[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_16 (.CI(n22746), .I0(n6671[13]), .I1(n1108_adj_4226), 
            .CO(n22747));
    SB_LUT4 add_3387_15_lut (.I0(GND_net), .I1(n6671[12]), .I2(n1035_adj_4225), 
            .I3(n22745), .O(n6650[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_15 (.CI(n22745), .I0(n6671[12]), .I1(n1035_adj_4225), 
            .CO(n22746));
    SB_LUT4 add_3387_14_lut (.I0(GND_net), .I1(n6671[11]), .I2(n962_adj_4224), 
            .I3(n22744), .O(n6650[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_14 (.CI(n22744), .I0(n6671[11]), .I1(n962_adj_4224), 
            .CO(n22745));
    SB_LUT4 add_3387_13_lut (.I0(GND_net), .I1(n6671[10]), .I2(n889_adj_4223), 
            .I3(n22743), .O(n6650[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_13 (.CI(n22743), .I0(n6671[10]), .I1(n889_adj_4223), 
            .CO(n22744));
    SB_LUT4 add_3387_12_lut (.I0(GND_net), .I1(n6671[9]), .I2(n816_adj_4222), 
            .I3(n22742), .O(n6650[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_12 (.CI(n22742), .I0(n6671[9]), .I1(n816_adj_4222), 
            .CO(n22743));
    SB_LUT4 add_3387_11_lut (.I0(GND_net), .I1(n6671[8]), .I2(n743_adj_4221), 
            .I3(n22741), .O(n6650[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_11 (.CI(n22741), .I0(n6671[8]), .I1(n743_adj_4221), 
            .CO(n22742));
    SB_LUT4 add_3387_10_lut (.I0(GND_net), .I1(n6671[7]), .I2(n670_adj_4220), 
            .I3(n22740), .O(n6650[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_10 (.CI(n22740), .I0(n6671[7]), .I1(n670_adj_4220), 
            .CO(n22741));
    SB_LUT4 add_3387_9_lut (.I0(GND_net), .I1(n6671[6]), .I2(n597_adj_4219), 
            .I3(n22739), .O(n6650[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_9 (.CI(n22739), .I0(n6671[6]), .I1(n597_adj_4219), 
            .CO(n22740));
    SB_LUT4 add_3387_8_lut (.I0(GND_net), .I1(n6671[5]), .I2(n524_adj_4218), 
            .I3(n22738), .O(n6650[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_8 (.CI(n22738), .I0(n6671[5]), .I1(n524_adj_4218), 
            .CO(n22739));
    SB_LUT4 add_3387_7_lut (.I0(GND_net), .I1(n6671[4]), .I2(n451_adj_4217), 
            .I3(n22737), .O(n6650[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_7 (.CI(n22737), .I0(n6671[4]), .I1(n451_adj_4217), 
            .CO(n22738));
    SB_LUT4 add_3387_6_lut (.I0(GND_net), .I1(n6671[3]), .I2(n378_adj_4216), 
            .I3(n22736), .O(n6650[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n22167), .I0(GND_net), .I1(n1[6]), 
            .CO(n22168));
    SB_CARRY add_3387_6 (.CI(n22736), .I0(n6671[3]), .I1(n378_adj_4216), 
            .CO(n22737));
    SB_LUT4 add_3387_5_lut (.I0(GND_net), .I1(n6671[2]), .I2(n305_adj_4210), 
            .I3(n22735), .O(n6650[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_5 (.CI(n22735), .I0(n6671[2]), .I1(n305_adj_4210), 
            .CO(n22736));
    SB_LUT4 add_3387_4_lut (.I0(GND_net), .I1(n6671[1]), .I2(n232_adj_4208), 
            .I3(n22734), .O(n6650[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_4 (.CI(n22734), .I0(n6671[1]), .I1(n232_adj_4208), 
            .CO(n22735));
    SB_LUT4 add_3387_3_lut (.I0(GND_net), .I1(n6671[0]), .I2(n159_adj_4207), 
            .I3(n22733), .O(n6650[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4211));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3387_3 (.CI(n22733), .I0(n6671[0]), .I1(n159_adj_4207), 
            .CO(n22734));
    SB_CARRY mult_11_add_1225_19 (.CI(n22931), .I0(n6878[16]), .I1(GND_net), 
            .CO(n22932));
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4209));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n6878[15]), .I2(GND_net), 
            .I3(n22930), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n22930), .I0(n6878[15]), .I1(GND_net), 
            .CO(n22931));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n6878[14]), .I2(GND_net), 
            .I3(n22929), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n22929), .I0(n6878[14]), .I1(GND_net), 
            .CO(n22930));
    SB_LUT4 add_3387_2_lut (.I0(GND_net), .I1(n17_adj_4206), .I2(n86_adj_4205), 
            .I3(GND_net), .O(n6650[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_2 (.CI(GND_net), .I0(n17_adj_4206), .I1(n86_adj_4205), 
            .CO(n22733));
    SB_LUT4 add_3386_21_lut (.I0(GND_net), .I1(n6650[18]), .I2(GND_net), 
            .I3(n22732), .O(n6628[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_20_lut (.I0(GND_net), .I1(n6650[17]), .I2(GND_net), 
            .I3(n22731), .O(n6628[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_20 (.CI(n22731), .I0(n6650[17]), .I1(GND_net), .CO(n22732));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n22166), .O(n11_adj_3905)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n22166), .I0(GND_net), .I1(n1[5]), 
            .CO(n22167));
    SB_LUT4 i25163_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n30253));   // verilog/motorControl.v(29[14] 48[8])
    defparam i25163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3386_19_lut (.I0(GND_net), .I1(n6650[16]), .I2(GND_net), 
            .I3(n22730), .O(n6628[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_19 (.CI(n22730), .I0(n6650[16]), .I1(GND_net), .CO(n22731));
    SB_LUT4 add_3386_18_lut (.I0(GND_net), .I1(n6650[15]), .I2(GND_net), 
            .I3(n22729), .O(n6628[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_18 (.CI(n22729), .I0(n6650[15]), .I1(GND_net), .CO(n22730));
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n6878[13]), .I2(n1096_adj_4203), 
            .I3(n22928), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3386_17_lut (.I0(GND_net), .I1(n6650[14]), .I2(GND_net), 
            .I3(n22728), .O(n6628[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_17 (.CI(n22728), .I0(n6650[14]), .I1(GND_net), .CO(n22729));
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_16 (.CI(n22928), .I0(n6878[13]), .I1(n1096_adj_4203), 
            .CO(n22929));
    SB_LUT4 add_3386_16_lut (.I0(GND_net), .I1(n6650[13]), .I2(n1105_adj_4201), 
            .I3(n22727), .O(n6628[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n6878[12]), .I2(n1023_adj_4199), 
            .I3(n22927), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_16 (.CI(n22727), .I0(n6650[13]), .I1(n1105_adj_4201), 
            .CO(n22728));
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4200));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_15 (.CI(n22927), .I0(n6878[12]), .I1(n1023_adj_4199), 
            .CO(n22928));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4198));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_15_lut (.I0(GND_net), .I1(n6650[12]), .I2(n1032_adj_4196), 
            .I3(n22726), .O(n6628[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n6878[11]), .I2(n950_adj_4195), 
            .I3(n22926), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_15 (.CI(n22726), .I0(n6650[12]), .I1(n1032_adj_4196), 
            .CO(n22727));
    SB_LUT4 add_3386_14_lut (.I0(GND_net), .I1(n6650[11]), .I2(n959_adj_4194), 
            .I3(n22725), .O(n6628[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4197));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1464 (.I0(n6_adj_4228), .I1(\Ki[4] ), .I2(n7157[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n7150[3]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1464.LUT_INIT = 16'h965a;
    SB_CARRY add_3386_14 (.CI(n22725), .I0(n6650[11]), .I1(n959_adj_4194), 
            .CO(n22726));
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3386_13_lut (.I0(GND_net), .I1(n6650[10]), .I2(n886_adj_4192), 
            .I3(n22724), .O(n6628[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_13 (.CI(n22724), .I0(n6650[10]), .I1(n886_adj_4192), 
            .CO(n22725));
    SB_CARRY mult_11_add_1225_14 (.CI(n22926), .I0(n6878[11]), .I1(n950_adj_4195), 
            .CO(n22927));
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_4229));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4191));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4190));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n6878[10]), .I2(n877_adj_4187), 
            .I3(n22925), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4189));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_12_lut (.I0(GND_net), .I1(n6650[9]), .I2(n813_adj_4184), 
            .I3(n22723), .O(n6628[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4186));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_12 (.CI(n22723), .I0(n6650[9]), .I1(n813_adj_4184), 
            .CO(n22724));
    SB_CARRY mult_11_add_1225_13 (.CI(n22925), .I0(n6878[10]), .I1(n877_adj_4187), 
            .CO(n22926));
    SB_LUT4 add_3386_11_lut (.I0(GND_net), .I1(n6650[8]), .I2(n740_adj_4180), 
            .I3(n22722), .O(n6628[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18054_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n7168[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18054_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_3386_11 (.CI(n22722), .I0(n6650[8]), .I1(n740_adj_4180), 
            .CO(n22723));
    SB_LUT4 add_3386_10_lut (.I0(GND_net), .I1(n6650[7]), .I2(n667_adj_4179), 
            .I3(n22721), .O(n6628[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4185));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n22165), .O(n9_adj_3907)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3386_10 (.CI(n22721), .I0(n6650[7]), .I1(n667_adj_4179), 
            .CO(n22722));
    SB_LUT4 add_3386_9_lut (.I0(GND_net), .I1(n6650[6]), .I2(n594_adj_4175), 
            .I3(n22720), .O(n6628[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n6878[9]), .I2(n804_adj_4174), 
            .I3(n22924), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_9 (.CI(n22720), .I0(n6650[6]), .I1(n594_adj_4175), 
            .CO(n22721));
    SB_LUT4 add_3386_8_lut (.I0(GND_net), .I1(n6650[5]), .I2(n521_adj_4170), 
            .I3(n22719), .O(n6628[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_8 (.CI(n22719), .I0(n6650[5]), .I1(n521_adj_4170), 
            .CO(n22720));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n22165), .I0(GND_net), .I1(n1[4]), 
            .CO(n22166));
    SB_LUT4 add_3386_7_lut (.I0(GND_net), .I1(n6650[4]), .I2(n448_adj_4167), 
            .I3(n22718), .O(n6628[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4183));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_12 (.CI(n22924), .I0(n6878[9]), .I1(n804_adj_4174), 
            .CO(n22925));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n6878[8]), .I2(n731_adj_4166), 
            .I3(n22923), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4182));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4181));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_11 (.CI(n22923), .I0(n6878[8]), .I1(n731_adj_4166), 
            .CO(n22924));
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n6878[7]), .I2(n658_adj_4163), 
            .I3(n22922), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_7 (.CI(n22718), .I0(n6650[4]), .I1(n448_adj_4167), 
            .CO(n22719));
    SB_CARRY mult_11_add_1225_10 (.CI(n22922), .I0(n6878[7]), .I1(n658_adj_4163), 
            .CO(n22923));
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4177));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4176));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_6_lut (.I0(GND_net), .I1(n6650[3]), .I2(n375_adj_4161), 
            .I3(n22717), .O(n6628[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_6 (.CI(n22717), .I0(n6650[3]), .I1(n375_adj_4161), 
            .CO(n22718));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n6878[6]), .I2(n585_adj_4160), 
            .I3(n22921), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3386_5_lut (.I0(GND_net), .I1(n6650[2]), .I2(n302_adj_4159), 
            .I3(n22716), .O(n6628[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n22921), .I0(n6878[6]), .I1(n585_adj_4160), 
            .CO(n22922));
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n6878[5]), .I2(n512_adj_4158), 
            .I3(n22920), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n22920), .I0(n6878[5]), .I1(n512_adj_4158), 
            .CO(n22921));
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4173));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4172));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n6878[4]), .I2(n439_adj_4157), 
            .I3(n22919), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n22919), .I0(n6878[4]), .I1(n439_adj_4157), 
            .CO(n22920));
    SB_CARRY add_3386_5 (.CI(n22716), .I0(n6650[2]), .I1(n302_adj_4159), 
            .CO(n22717));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n6878[3]), .I2(n366_adj_4156), 
            .I3(n22918), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n22918), .I0(n6878[3]), .I1(n366_adj_4156), 
            .CO(n22919));
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4171));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_4233));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_4234));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3386_4_lut (.I0(GND_net), .I1(n6650[1]), .I2(n229_adj_4155), 
            .I3(n22715), .O(n6628[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n6878[2]), .I2(n293_adj_4154), 
            .I3(n22917), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_4 (.CI(n22715), .I0(n6650[1]), .I1(n229_adj_4155), 
            .CO(n22716));
    SB_LUT4 add_3386_3_lut (.I0(GND_net), .I1(n6650[0]), .I2(n156_adj_4153), 
            .I3(n22714), .O(n6628[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3386_3 (.CI(n22714), .I0(n6650[0]), .I1(n156_adj_4153), 
            .CO(n22715));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n22164), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3386_2_lut (.I0(GND_net), .I1(n14_adj_4152), .I2(n83_adj_4151), 
            .I3(GND_net), .O(n6628[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3386_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4169));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3386_2 (.CI(GND_net), .I0(n14_adj_4152), .I1(n83_adj_4151), 
            .CO(n22714));
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4168));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4165));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1465 (.I0(n4_adj_4235), .I1(\Ki[3] ), .I2(n7163[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n7157[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1465.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4164));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_22_lut (.I0(GND_net), .I1(n6628[19]), .I2(GND_net), 
            .I3(n22713), .O(n6605[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4162));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_21_lut (.I0(GND_net), .I1(n6628[18]), .I2(GND_net), 
            .I3(n22712), .O(n6605[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_21 (.CI(n22712), .I0(n6628[18]), .I1(GND_net), .CO(n22713));
    SB_LUT4 add_3385_20_lut (.I0(GND_net), .I1(n6628[17]), .I2(GND_net), 
            .I3(n22711), .O(n6605[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_20 (.CI(n22711), .I0(n6628[17]), .I1(GND_net), .CO(n22712));
    SB_LUT4 add_3385_19_lut (.I0(GND_net), .I1(n6628[16]), .I2(GND_net), 
            .I3(n22710), .O(n6605[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_19 (.CI(n22710), .I0(n6628[16]), .I1(GND_net), .CO(n22711));
    SB_LUT4 add_3385_18_lut (.I0(GND_net), .I1(n6628[15]), .I2(GND_net), 
            .I3(n22709), .O(n6605[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_18 (.CI(n22709), .I0(n6628[15]), .I1(GND_net), .CO(n22710));
    SB_CARRY mult_11_add_1225_5 (.CI(n22917), .I0(n6878[2]), .I1(n293_adj_4154), 
            .CO(n22918));
    SB_LUT4 add_3385_17_lut (.I0(GND_net), .I1(n6628[14]), .I2(GND_net), 
            .I3(n22708), .O(n6605[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n6878[1]), .I2(n220_adj_4150), 
            .I3(n22916), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_17 (.CI(n22708), .I0(n6628[14]), .I1(GND_net), .CO(n22709));
    SB_CARRY mult_11_add_1225_4 (.CI(n22916), .I0(n6878[1]), .I1(n220_adj_4150), 
            .CO(n22917));
    SB_LUT4 add_3385_16_lut (.I0(GND_net), .I1(n6628[13]), .I2(n1102_adj_4149), 
            .I3(n22707), .O(n6605[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n6878[0]), .I2(n147_adj_4148), 
            .I3(n22915), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n22915), .I0(n6878[0]), .I1(n147_adj_4148), 
            .CO(n22916));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4147), .I2(n74_adj_4144), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4147), .I1(n74_adj_4144), 
            .CO(n22915));
    SB_LUT4 add_3406_23_lut (.I0(GND_net), .I1(n6902[20]), .I2(GND_net), 
            .I3(n22914), .O(n6878[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3406_22_lut (.I0(GND_net), .I1(n6902[19]), .I2(GND_net), 
            .I3(n22913), .O(n6878[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_22 (.CI(n22913), .I0(n6902[19]), .I1(GND_net), .CO(n22914));
    SB_LUT4 add_3406_21_lut (.I0(GND_net), .I1(n6902[18]), .I2(GND_net), 
            .I3(n22912), .O(n6878[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_21 (.CI(n22912), .I0(n6902[18]), .I1(GND_net), .CO(n22913));
    SB_LUT4 add_3406_20_lut (.I0(GND_net), .I1(n6902[17]), .I2(GND_net), 
            .I3(n22911), .O(n6878[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_20 (.CI(n22911), .I0(n6902[17]), .I1(GND_net), .CO(n22912));
    SB_LUT4 add_3406_19_lut (.I0(GND_net), .I1(n6902[16]), .I2(GND_net), 
            .I3(n22910), .O(n6878[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_19 (.CI(n22910), .I0(n6902[16]), .I1(GND_net), .CO(n22911));
    SB_LUT4 add_3406_18_lut (.I0(GND_net), .I1(n6902[15]), .I2(GND_net), 
            .I3(n22909), .O(n6878[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4146));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3385_16 (.CI(n22707), .I0(n6628[13]), .I1(n1102_adj_4149), 
            .CO(n22708));
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4145));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_15_lut (.I0(GND_net), .I1(n6628[12]), .I2(n1029_adj_4140), 
            .I3(n22706), .O(n6605[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_18 (.CI(n22909), .I0(n6902[15]), .I1(GND_net), .CO(n22910));
    SB_LUT4 add_3406_17_lut (.I0(GND_net), .I1(n6902[14]), .I2(GND_net), 
            .I3(n22908), .O(n6878[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_17 (.CI(n22908), .I0(n6902[14]), .I1(GND_net), .CO(n22909));
    SB_LUT4 add_3406_16_lut (.I0(GND_net), .I1(n6902[13]), .I2(n1099_adj_4139), 
            .I3(n22907), .O(n6878[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_16 (.CI(n22907), .I0(n6902[13]), .I1(n1099_adj_4139), 
            .CO(n22908));
    SB_LUT4 add_3406_15_lut (.I0(GND_net), .I1(n6902[12]), .I2(n1026_adj_4135), 
            .I3(n22906), .O(n6878[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_15 (.CI(n22906), .I0(n6902[12]), .I1(n1026_adj_4135), 
            .CO(n22907));
    SB_LUT4 add_3406_14_lut (.I0(GND_net), .I1(n6902[11]), .I2(n953_adj_4130), 
            .I3(n22905), .O(n6878[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_14 (.CI(n22905), .I0(n6902[11]), .I1(n953_adj_4130), 
            .CO(n22906));
    SB_LUT4 add_3406_13_lut (.I0(GND_net), .I1(n6902[10]), .I2(n880_adj_4127), 
            .I3(n22904), .O(n6878[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_13 (.CI(n22904), .I0(n6902[10]), .I1(n880_adj_4127), 
            .CO(n22905));
    SB_LUT4 add_3406_12_lut (.I0(GND_net), .I1(n6902[9]), .I2(n807_adj_4126), 
            .I3(n22903), .O(n6878[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_12 (.CI(n22903), .I0(n6902[9]), .I1(n807_adj_4126), 
            .CO(n22904));
    SB_LUT4 add_3406_11_lut (.I0(GND_net), .I1(n6902[8]), .I2(n734_adj_4124), 
            .I3(n22902), .O(n6878[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_11 (.CI(n22902), .I0(n6902[8]), .I1(n734_adj_4124), 
            .CO(n22903));
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4143));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4142));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4141));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4138));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4137));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3385_15 (.CI(n22706), .I0(n6628[12]), .I1(n1029_adj_4140), 
            .CO(n22707));
    SB_LUT4 add_3406_10_lut (.I0(GND_net), .I1(n6902[7]), .I2(n661_adj_4122), 
            .I3(n22901), .O(n6878[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_10 (.CI(n22901), .I0(n6902[7]), .I1(n661_adj_4122), 
            .CO(n22902));
    SB_LUT4 add_3385_14_lut (.I0(GND_net), .I1(n6628[11]), .I2(n956), 
            .I3(n22705), .O(n6605[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3406_9_lut (.I0(GND_net), .I1(n6902[6]), .I2(n588_adj_4103), 
            .I3(n22900), .O(n6878[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_14 (.CI(n22705), .I0(n6628[11]), .I1(n956), .CO(n22706));
    SB_LUT4 add_3385_13_lut (.I0(GND_net), .I1(n6628[10]), .I2(n883), 
            .I3(n22704), .O(n6605[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_13 (.CI(n22704), .I0(n6628[10]), .I1(n883), .CO(n22705));
    SB_CARRY add_3406_9 (.CI(n22900), .I0(n6902[6]), .I1(n588_adj_4103), 
            .CO(n22901));
    SB_LUT4 add_3406_8_lut (.I0(GND_net), .I1(n6902[5]), .I2(n515_adj_4102), 
            .I3(n22899), .O(n6878[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3385_12_lut (.I0(GND_net), .I1(n6628[9]), .I2(n810), .I3(n22703), 
            .O(n6605[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_12 (.CI(n22703), .I0(n6628[9]), .I1(n810), .CO(n22704));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n22164), .I0(GND_net), .I1(n1[3]), 
            .CO(n22165));
    SB_LUT4 add_3385_11_lut (.I0(GND_net), .I1(n6628[8]), .I2(n737), .I3(n22702), 
            .O(n6605[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n22163), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3385_11 (.CI(n22702), .I0(n6628[8]), .I1(n737), .CO(n22703));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n22163), .I0(GND_net), .I1(n1[2]), 
            .CO(n22164));
    SB_LUT4 add_3385_10_lut (.I0(GND_net), .I1(n6628[7]), .I2(n664), .I3(n22701), 
            .O(n6605[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_10 (.CI(n22701), .I0(n6628[7]), .I1(n664), .CO(n22702));
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4134));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_8 (.CI(n22899), .I0(n6902[5]), .I1(n515_adj_4102), 
            .CO(n22900));
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4133));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4132));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4131));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_9_lut (.I0(GND_net), .I1(n6628[6]), .I2(n591), .I3(n22700), 
            .O(n6605[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3406_7_lut (.I0(GND_net), .I1(n6902[4]), .I2(n442_adj_4098), 
            .I3(n22898), .O(n6878[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4129));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3406_7 (.CI(n22898), .I0(n6902[4]), .I1(n442_adj_4098), 
            .CO(n22899));
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4128));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3385_9 (.CI(n22700), .I0(n6628[6]), .I1(n591), .CO(n22701));
    SB_LUT4 add_3385_8_lut (.I0(GND_net), .I1(n6628[5]), .I2(n518), .I3(n22699), 
            .O(n6605[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3406_6_lut (.I0(GND_net), .I1(n6902[3]), .I2(n369_adj_4097), 
            .I3(n22897), .O(n6878[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3406_6 (.CI(n22897), .I0(n6902[3]), .I1(n369_adj_4097), 
            .CO(n22898));
    SB_LUT4 add_3406_5_lut (.I0(GND_net), .I1(n6902[2]), .I2(n296_adj_4096), 
            .I3(n22896), .O(n6878[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_5 (.CI(n22896), .I0(n6902[2]), .I1(n296_adj_4096), 
            .CO(n22897));
    SB_LUT4 add_3406_4_lut (.I0(GND_net), .I1(n6902[1]), .I2(n223_adj_4095), 
            .I3(n22895), .O(n6878[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_8 (.CI(n22699), .I0(n6628[5]), .I1(n518), .CO(n22700));
    SB_LUT4 add_3385_7_lut (.I0(GND_net), .I1(n6628[4]), .I2(n445), .I3(n22698), 
            .O(n6605[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_7 (.CI(n22698), .I0(n6628[4]), .I1(n445), .CO(n22699));
    SB_CARRY add_3406_4 (.CI(n22895), .I0(n6902[1]), .I1(n223_adj_4095), 
            .CO(n22896));
    SB_LUT4 add_3406_3_lut (.I0(GND_net), .I1(n6902[0]), .I2(n150_adj_4094), 
            .I3(n22894), .O(n6878[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_3 (.CI(n22894), .I0(n6902[0]), .I1(n150_adj_4094), 
            .CO(n22895));
    SB_LUT4 add_3406_2_lut (.I0(GND_net), .I1(n8_adj_4093), .I2(n77_adj_4092), 
            .I3(GND_net), .O(n6878[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3406_2 (.CI(GND_net), .I0(n8_adj_4093), .I1(n77_adj_4092), 
            .CO(n22894));
    SB_LUT4 add_3400_7_lut (.I0(GND_net), .I1(n27329), .I2(n490_adj_4086), 
            .I3(n22893), .O(n6845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4123));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3385_6_lut (.I0(GND_net), .I1(n6628[3]), .I2(n372), .I3(n22697), 
            .O(n6605[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_6 (.CI(n22697), .I0(n6628[3]), .I1(n372), .CO(n22698));
    SB_LUT4 add_3385_5_lut (.I0(GND_net), .I1(n6628[2]), .I2(n299), .I3(n22696), 
            .O(n6605[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_5 (.CI(n22696), .I0(n6628[2]), .I1(n299), .CO(n22697));
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n22162), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3400_6_lut (.I0(GND_net), .I1(n6853[3]), .I2(n417_adj_4079), 
            .I3(n22892), .O(n6845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_6 (.CI(n22892), .I0(n6853[3]), .I1(n417_adj_4079), 
            .CO(n22893));
    SB_LUT4 add_3400_5_lut (.I0(GND_net), .I1(n6853[2]), .I2(n344_adj_4078), 
            .I3(n22891), .O(n6845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3385_4_lut (.I0(GND_net), .I1(n6628[1]), .I2(n226), .I3(n22695), 
            .O(n6605[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_5 (.CI(n22891), .I0(n6853[2]), .I1(n344_adj_4078), 
            .CO(n22892));
    SB_LUT4 add_3400_4_lut (.I0(GND_net), .I1(n6853[1]), .I2(n271_adj_4076), 
            .I3(n22890), .O(n6845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_4 (.CI(n22890), .I0(n6853[1]), .I1(n271_adj_4076), 
            .CO(n22891));
    SB_LUT4 add_3400_3_lut (.I0(GND_net), .I1(n6853[0]), .I2(n198_adj_4075), 
            .I3(n22889), .O(n6845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n22162), .I0(GND_net), .I1(n1[1]), 
            .CO(n22163));
    SB_CARRY add_3400_3 (.CI(n22889), .I0(n6853[0]), .I1(n198_adj_4075), 
            .CO(n22890));
    SB_LUT4 add_3400_2_lut (.I0(GND_net), .I1(n56_adj_4074), .I2(n125_adj_4072), 
            .I3(GND_net), .O(n6845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_2 (.CI(GND_net), .I0(n56_adj_4074), .I1(n125_adj_4072), 
            .CO(n22889));
    SB_LUT4 add_3399_8_lut (.I0(GND_net), .I1(n6845[5]), .I2(n560_adj_4071), 
            .I3(n22888), .O(n6836[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3399_7_lut (.I0(GND_net), .I1(n6845[4]), .I2(n487_adj_4070), 
            .I3(n22887), .O(n6836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3467 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_4 (.CI(n22695), .I0(n6628[1]), .I1(n226), .CO(n22696));
    SB_LUT4 add_3385_3_lut (.I0(GND_net), .I1(n6628[0]), .I2(n153), .I3(n22694), 
            .O(n6605[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_7 (.CI(n22887), .I0(n6845[4]), .I1(n487_adj_4070), 
            .CO(n22888));
    SB_LUT4 add_3399_6_lut (.I0(GND_net), .I1(n6845[3]), .I2(n414_adj_4066), 
            .I3(n22886), .O(n6836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_6 (.CI(n22886), .I0(n6845[3]), .I1(n414_adj_4066), 
            .CO(n22887));
    SB_CARRY add_3385_3 (.CI(n22694), .I0(n6628[0]), .I1(n153), .CO(n22695));
    SB_LUT4 add_3399_5_lut (.I0(GND_net), .I1(n6845[2]), .I2(n341_adj_4065), 
            .I3(n22885), .O(n6836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n22162));
    SB_CARRY add_3399_5 (.CI(n22885), .I0(n6845[2]), .I1(n341_adj_4065), 
            .CO(n22886));
    SB_LUT4 add_3399_4_lut (.I0(GND_net), .I1(n6845[1]), .I2(n268_adj_4064), 
            .I3(n22884), .O(n6836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_4 (.CI(n22884), .I0(n6845[1]), .I1(n268_adj_4064), 
            .CO(n22885));
    SB_LUT4 add_3399_3_lut (.I0(GND_net), .I1(n6845[0]), .I2(n195_adj_4062), 
            .I3(n22883), .O(n6836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_3 (.CI(n22883), .I0(n6845[0]), .I1(n195_adj_4062), 
            .CO(n22884));
    SB_LUT4 add_3385_2_lut (.I0(GND_net), .I1(n11_adj_4061), .I2(n80), 
            .I3(GND_net), .O(n6605[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3385_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3399_2_lut (.I0(GND_net), .I1(n53_adj_4060), .I2(n122_adj_4059), 
            .I3(GND_net), .O(n6836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3399_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3399_2 (.CI(GND_net), .I0(n53_adj_4060), .I1(n122_adj_4059), 
            .CO(n22883));
    SB_LUT4 add_3398_9_lut (.I0(GND_net), .I1(n6836[6]), .I2(n630_adj_4058), 
            .I3(n22882), .O(n6826[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3398_8_lut (.I0(GND_net), .I1(n6836[5]), .I2(n557_adj_4055), 
            .I3(n22881), .O(n6826[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3398_8 (.CI(n22881), .I0(n6836[5]), .I1(n557_adj_4055), 
            .CO(n22882));
    SB_LUT4 add_3398_7_lut (.I0(GND_net), .I1(n6836[4]), .I2(n484_adj_4054), 
            .I3(n22880), .O(n6826[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3385_2 (.CI(GND_net), .I0(n11_adj_4061), .I1(n80), .CO(n22694));
    SB_CARRY add_3398_7 (.CI(n22880), .I0(n6836[4]), .I1(n484_adj_4054), 
            .CO(n22881));
    SB_LUT4 add_3398_6_lut (.I0(GND_net), .I1(n6836[3]), .I2(n411_adj_4050), 
            .I3(n22879), .O(n6826[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3398_6 (.CI(n22879), .I0(n6836[3]), .I1(n411_adj_4050), 
            .CO(n22880));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n6581[21]), 
            .I2(GND_net), .I3(n22693), .O(n5022[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1466 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4236));   // verilog/motorControl.v(34[26:37])
    defparam i2_4_lut_adj_1466.LUT_INIT = 16'h9c50;
    SB_LUT4 i17990_4_lut (.I0(n7157[2]), .I1(\Ki[4] ), .I2(n6_adj_4228), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4237));   // verilog/motorControl.v(34[26:37])
    defparam i17990_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1467 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4238));   // verilog/motorControl.v(34[26:37])
    defparam i1_4_lut_adj_1467.LUT_INIT = 16'h6ca0;
    SB_LUT4 i18021_4_lut (.I0(n7163[1]), .I1(\Ki[3] ), .I2(n4_adj_4235), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4239));   // verilog/motorControl.v(34[26:37])
    defparam i18021_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i18056_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n21877));   // verilog/motorControl.v(34[26:37])
    defparam i18056_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1468 (.I0(n6_adj_4239), .I1(n11_adj_4238), .I2(n8_adj_4237), 
            .I3(n12_adj_4236), .O(n18_adj_4240));   // verilog/motorControl.v(34[26:37])
    defparam i8_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1469 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4241));   // verilog/motorControl.v(34[26:37])
    defparam i3_4_lut_adj_1469.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1470 (.I0(n13_adj_4241), .I1(n18_adj_4240), .I2(n21877), 
            .I3(n4_adj_4242), .O(n27773));   // verilog/motorControl.v(34[26:37])
    defparam i9_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4120));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n18679), .I1(n6581[20]), .I2(GND_net), 
            .I3(n22692), .O(n2529[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_23 (.CI(n22692), .I0(n6581[20]), .I1(GND_net), 
            .CO(n22693));
    SB_LUT4 add_3398_5_lut (.I0(GND_net), .I1(n6836[2]), .I2(n338_adj_4014), 
            .I3(n22878), .O(n6826[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n18679), .I1(n6581[19]), .I2(GND_net), 
            .I3(n22691), .O(n2529[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3398_5 (.CI(n22878), .I0(n6836[2]), .I1(n338_adj_4014), 
            .CO(n22879));
    SB_LUT4 add_3398_4_lut (.I0(GND_net), .I1(n6836[1]), .I2(n265_adj_4013), 
            .I3(n22877), .O(n6826[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3398_4 (.CI(n22877), .I0(n6836[1]), .I1(n265_adj_4013), 
            .CO(n22878));
    SB_LUT4 add_3398_3_lut (.I0(GND_net), .I1(n6836[0]), .I2(n192_adj_4012), 
            .I3(n22876), .O(n6826[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n22691), .I0(n6581[19]), .I1(GND_net), 
            .CO(n22692));
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4118));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n18679), .I1(n6581[18]), .I2(GND_net), 
            .I3(n22690), .O(n2529[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3398_3 (.CI(n22876), .I0(n6836[0]), .I1(n192_adj_4012), 
            .CO(n22877));
    SB_LUT4 add_3398_2_lut (.I0(GND_net), .I1(n50_adj_4011), .I2(n119_adj_4010), 
            .I3(GND_net), .O(n6826[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3398_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3398_2 (.CI(GND_net), .I0(n50_adj_4011), .I1(n119_adj_4010), 
            .CO(n22876));
    SB_CARRY add_3394_9 (.CI(n22844), .I0(n6790[6]), .I1(n618_adj_4008), 
            .CO(n22845));
    SB_CARRY mult_10_add_1225_21 (.CI(n22690), .I0(n6581[18]), .I1(GND_net), 
            .CO(n22691));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n18679), .I1(n6581[17]), .I2(GND_net), 
            .I3(n22689), .O(n2529[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_20 (.CI(n22689), .I0(n6581[17]), .I1(GND_net), 
            .CO(n22690));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n18679), .I1(n6581[16]), .I2(GND_net), 
            .I3(n22688), .O(n2529[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_19 (.CI(n22688), .I0(n6581[16]), .I1(GND_net), 
            .CO(n22689));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n18679), .I1(n6581[15]), .I2(GND_net), 
            .I3(n22687), .O(n2529[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_18 (.CI(n22687), .I0(n6581[15]), .I1(GND_net), 
            .CO(n22688));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n18679), .I1(n6581[14]), .I2(GND_net), 
            .I3(n22686), .O(n2529[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_17 (.CI(n22686), .I0(n6581[14]), .I1(GND_net), 
            .CO(n22687));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n18679), .I1(n6581[13]), .I2(n1096), 
            .I3(n22685), .O(n2529[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_16 (.CI(n22685), .I0(n6581[13]), .I1(n1096), 
            .CO(n22686));
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n18679), .I1(n6581[12]), .I2(n1023), 
            .I3(n22684), .O(n2529[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_15 (.CI(n22684), .I0(n6581[12]), .I1(n1023), 
            .CO(n22685));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n18679), .I1(n6581[11]), .I2(n950), 
            .I3(n22683), .O(n2529[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_14 (.CI(n22683), .I0(n6581[11]), .I1(n950), 
            .CO(n22684));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n18679), .I1(n6581[10]), .I2(n877), 
            .I3(n22682), .O(n2529[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n22682), .I0(n6581[10]), .I1(n877), 
            .CO(n22683));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n18679), .I1(n6581[9]), .I2(n804), 
            .I3(n22681), .O(n2529[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_12 (.CI(n22681), .I0(n6581[9]), .I1(n804), 
            .CO(n22682));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n18679), .I1(n6581[8]), .I2(n731), 
            .I3(n22680), .O(n2529[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_11 (.CI(n22680), .I0(n6581[8]), .I1(n731), 
            .CO(n22681));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n18679), .I1(n6581[7]), .I2(n658), 
            .I3(n22679), .O(n2529[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_10 (.CI(n22679), .I0(n6581[7]), .I1(n658), 
            .CO(n22680));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n18679), .I1(n6581[6]), .I2(n585), 
            .I3(n22678), .O(n2529[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_9 (.CI(n22678), .I0(n6581[6]), .I1(n585), 
            .CO(n22679));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4115));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[15]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n18679), .I1(n6581[5]), .I2(n512), 
            .I3(n22677), .O(n2529[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_8 (.CI(n22677), .I0(n6581[5]), .I1(n512), 
            .CO(n22678));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n18679), .I1(n6581[4]), .I2(n439), 
            .I3(n22676), .O(n2529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_7 (.CI(n22676), .I0(n6581[4]), .I1(n439), 
            .CO(n22677));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n18679), .I1(n6581[3]), .I2(n366), 
            .I3(n22675), .O(n2529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4114));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_6 (.CI(n22675), .I0(n6581[3]), .I1(n366), 
            .CO(n22676));
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n18679), .I1(n6581[2]), .I2(n293), 
            .I3(n22674), .O(n2529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_5 (.CI(n22674), .I0(n6581[2]), .I1(n293), 
            .CO(n22675));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n18679), .I1(n6581[1]), .I2(n220), 
            .I3(n22673), .O(n2529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_4 (.CI(n22673), .I0(n6581[1]), .I1(n220), 
            .CO(n22674));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n18679), .I1(n6581[0]), .I2(n147), 
            .I3(n22672), .O(n2529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4113));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_3 (.CI(n22672), .I0(n6581[0]), .I1(n147), 
            .CO(n22673));
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n18679), .I1(n5_adj_4006), .I2(n74), 
            .I3(GND_net), .O(n2529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4006), .I1(n74), 
            .CO(n22672));
    SB_LUT4 add_3384_23_lut (.I0(GND_net), .I1(n6605[20]), .I2(GND_net), 
            .I3(n22671), .O(n6581[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3384_22_lut (.I0(GND_net), .I1(n6605[19]), .I2(GND_net), 
            .I3(n22670), .O(n6581[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_22 (.CI(n22670), .I0(n6605[19]), .I1(GND_net), .CO(n22671));
    SB_LUT4 add_3384_21_lut (.I0(GND_net), .I1(n6605[18]), .I2(GND_net), 
            .I3(n22669), .O(n6581[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_21 (.CI(n22669), .I0(n6605[18]), .I1(GND_net), .CO(n22670));
    SB_LUT4 add_3384_20_lut (.I0(GND_net), .I1(n6605[17]), .I2(GND_net), 
            .I3(n22668), .O(n6581[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_20 (.CI(n22668), .I0(n6605[17]), .I1(GND_net), .CO(n22669));
    SB_LUT4 add_3384_19_lut (.I0(GND_net), .I1(n6605[16]), .I2(GND_net), 
            .I3(n22667), .O(n6581[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_19 (.CI(n22667), .I0(n6605[16]), .I1(GND_net), .CO(n22668));
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_18_lut (.I0(GND_net), .I1(n6605[15]), .I2(GND_net), 
            .I3(n22666), .O(n6581[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_18 (.CI(n22666), .I0(n6605[15]), .I1(GND_net), .CO(n22667));
    SB_LUT4 add_3384_17_lut (.I0(GND_net), .I1(n6605[14]), .I2(GND_net), 
            .I3(n22665), .O(n6581[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_17 (.CI(n22665), .I0(n6605[14]), .I1(GND_net), .CO(n22666));
    SB_LUT4 add_3384_16_lut (.I0(GND_net), .I1(n6605[13]), .I2(n1099), 
            .I3(n22664), .O(n6581[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_16 (.CI(n22664), .I0(n6605[13]), .I1(n1099), .CO(n22665));
    SB_LUT4 add_3384_15_lut (.I0(GND_net), .I1(n6605[12]), .I2(n1026), 
            .I3(n22663), .O(n6581[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_15 (.CI(n22663), .I0(n6605[12]), .I1(n1026), .CO(n22664));
    SB_LUT4 add_3384_14_lut (.I0(GND_net), .I1(n6605[11]), .I2(n953), 
            .I3(n22662), .O(n6581[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_14 (.CI(n22662), .I0(n6605[11]), .I1(n953), .CO(n22663));
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4112));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4111));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_13_lut (.I0(GND_net), .I1(n6605[10]), .I2(n880), 
            .I3(n22661), .O(n6581[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_13 (.CI(n22661), .I0(n6605[10]), .I1(n880), .CO(n22662));
    SB_LUT4 add_3384_12_lut (.I0(GND_net), .I1(n6605[9]), .I2(n807), .I3(n22660), 
            .O(n6581[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_12 (.CI(n22660), .I0(n6605[9]), .I1(n807), .CO(n22661));
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4110));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_11_lut (.I0(GND_net), .I1(n6605[8]), .I2(n734), .I3(n22659), 
            .O(n6581[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_11 (.CI(n22659), .I0(n6605[8]), .I1(n734), .CO(n22660));
    SB_LUT4 add_3384_10_lut (.I0(GND_net), .I1(n6605[7]), .I2(n661), .I3(n22658), 
            .O(n6581[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4109));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3384_10 (.CI(n22658), .I0(n6605[7]), .I1(n661), .CO(n22659));
    SB_LUT4 add_3384_9_lut (.I0(GND_net), .I1(n6605[6]), .I2(n588), .I3(n22657), 
            .O(n6581[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_9 (.CI(n22657), .I0(n6605[6]), .I1(n588), .CO(n22658));
    SB_LUT4 add_3384_8_lut (.I0(GND_net), .I1(n6605[5]), .I2(n515), .I3(n22656), 
            .O(n6581[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_8 (.CI(n22656), .I0(n6605[5]), .I1(n515), .CO(n22657));
    SB_LUT4 add_3384_7_lut (.I0(GND_net), .I1(n6605[4]), .I2(n442), .I3(n22655), 
            .O(n6581[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_7 (.CI(n22655), .I0(n6605[4]), .I1(n442), .CO(n22656));
    SB_LUT4 add_3384_6_lut (.I0(GND_net), .I1(n6605[3]), .I2(n369), .I3(n22654), 
            .O(n6581[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_6 (.CI(n22654), .I0(n6605[3]), .I1(n369), .CO(n22655));
    SB_LUT4 add_3384_5_lut (.I0(GND_net), .I1(n6605[2]), .I2(n296), .I3(n22653), 
            .O(n6581[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_5 (.CI(n22653), .I0(n6605[2]), .I1(n296), .CO(n22654));
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3384_4_lut (.I0(GND_net), .I1(n6605[1]), .I2(n223), .I3(n22652), 
            .O(n6581[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_4 (.CI(n22652), .I0(n6605[1]), .I1(n223), .CO(n22653));
    SB_LUT4 add_3384_3_lut (.I0(GND_net), .I1(n6605[0]), .I2(n150), .I3(n22651), 
            .O(n6581[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_3 (.CI(n22651), .I0(n6605[0]), .I1(n150), .CO(n22652));
    SB_LUT4 add_3384_2_lut (.I0(GND_net), .I1(n8_adj_4004), .I2(n77), 
            .I3(GND_net), .O(n6581[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3384_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3384_2 (.CI(GND_net), .I0(n8_adj_4004), .I1(n77), .CO(n22651));
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4108));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_3939));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4244));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4245));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4246));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4247));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4248));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4249));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4250));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4251));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4252));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4253));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4254));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4255));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4256));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4257));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4258));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4259));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4260));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4261));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4262));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24305_4_lut (.I0(n21_adj_4262), .I1(n19_adj_4261), .I2(n17_adj_4260), 
            .I3(n9_adj_4259), .O(n29395));
    defparam i24305_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24299_4_lut (.I0(n27_adj_4258), .I1(n15_adj_4257), .I2(n13_adj_4256), 
            .I3(n11_adj_4255), .O(n29389));
    defparam i24299_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_4263), .I1(duty[17]), .I2(n35_adj_4253), 
            .I3(GND_net), .O(n30_adj_4264));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24588_4_lut (.I0(n13_adj_4256), .I1(n11_adj_4255), .I2(n9_adj_4259), 
            .I3(n29405), .O(n29680));
    defparam i24588_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i24584_4_lut (.I0(n19_adj_4261), .I1(n17_adj_4260), .I2(n15_adj_4257), 
            .I3(n29680), .O(n29676));
    defparam i24584_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24918_4_lut (.I0(n25_adj_4252), .I1(n23_adj_4251), .I2(n21_adj_4262), 
            .I3(n29676), .O(n30010));
    defparam i24918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24759_4_lut (.I0(n31_adj_4249), .I1(n29_adj_4248), .I2(n27_adj_4258), 
            .I3(n30010), .O(n29851));
    defparam i24759_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i24978_4_lut (.I0(n37_adj_4247), .I1(n35_adj_4253), .I2(n33_adj_4254), 
            .I3(n29851), .O(n30070));
    defparam i24978_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24900_3_lut (.I0(n6_adj_4265), .I1(duty[10]), .I2(n21_adj_4262), 
            .I3(GND_net), .O(n29992));   // verilog/motorControl.v(36[10:25])
    defparam i24900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24901_3_lut (.I0(n29992), .I1(duty[11]), .I2(n23_adj_4251), 
            .I3(GND_net), .O(n29993));   // verilog/motorControl.v(36[10:25])
    defparam i24901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_4266), .I1(duty[22]), .I2(n45_adj_4246), 
            .I3(GND_net), .O(n24_adj_4267));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24284_4_lut (.I0(n43_adj_4250), .I1(n25_adj_4252), .I2(n23_adj_4251), 
            .I3(n29395), .O(n29374));
    defparam i24284_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3394_9_lut (.I0(GND_net), .I1(n6790[6]), .I2(n618_adj_4008), 
            .I3(n22844), .O(n6776[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3394_10 (.CI(n22845), .I0(n6790[7]), .I1(n691_adj_4002), 
            .CO(n22846));
    SB_LUT4 add_3394_10_lut (.I0(GND_net), .I1(n6790[7]), .I2(n691_adj_4002), 
            .I3(n22845), .O(n6776[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3394_11 (.CI(n22846), .I0(n6790[8]), .I1(n764_adj_4001), 
            .CO(n22847));
    SB_LUT4 add_3394_11_lut (.I0(GND_net), .I1(n6790[8]), .I2(n764_adj_4001), 
            .I3(n22846), .O(n6776[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3394_12 (.CI(n22847), .I0(n6790[9]), .I1(n837_adj_4000), 
            .CO(n22848));
    SB_LUT4 add_3394_12_lut (.I0(GND_net), .I1(n6790[9]), .I2(n837_adj_4000), 
            .I3(n22847), .O(n6776[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3394_13_lut (.I0(GND_net), .I1(n6790[10]), .I2(n910_adj_3999), 
            .I3(n22848), .O(n6776[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3394_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_2 (.CI(GND_net), .I0(n41_adj_3998), .I1(n110_adj_3997), 
            .CO(n22849));
    SB_LUT4 add_3395_2_lut (.I0(GND_net), .I1(n41_adj_3998), .I2(n110_adj_3997), 
            .I3(GND_net), .O(n6790[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_3 (.CI(n22849), .I0(n6803[0]), .I1(n183_adj_3996), 
            .CO(n22850));
    SB_LUT4 add_3395_3_lut (.I0(GND_net), .I1(n6803[0]), .I2(n183_adj_3996), 
            .I3(n22849), .O(n6790[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_4 (.CI(n22850), .I0(n6803[1]), .I1(n256_adj_3995), 
            .CO(n22851));
    SB_LUT4 i24781_4_lut (.I0(n24_adj_4267), .I1(n8_adj_4268), .I2(n45_adj_4246), 
            .I3(n29372), .O(n29873));   // verilog/motorControl.v(36[10:25])
    defparam i24781_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24860_3_lut (.I0(n29993), .I1(duty[12]), .I2(n25_adj_4252), 
            .I3(GND_net), .O(n29952));   // verilog/motorControl.v(36[10:25])
    defparam i24860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4269));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i24898_3_lut (.I0(n4_adj_4269), .I1(duty[13]), .I2(n27_adj_4258), 
            .I3(GND_net), .O(n29990));   // verilog/motorControl.v(36[10:25])
    defparam i24898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24899_3_lut (.I0(n29990), .I1(duty[14]), .I2(n29_adj_4248), 
            .I3(GND_net), .O(n29991));   // verilog/motorControl.v(36[10:25])
    defparam i24899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24295_4_lut (.I0(n33_adj_4254), .I1(n31_adj_4249), .I2(n29_adj_4248), 
            .I3(n29389), .O(n29385));
    defparam i24295_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24991_4_lut (.I0(n30_adj_4264), .I1(n10_adj_4270), .I2(n35_adj_4253), 
            .I3(n29383), .O(n30083));   // verilog/motorControl.v(36[10:25])
    defparam i24991_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i24862_3_lut (.I0(n29991), .I1(duty[15]), .I2(n31_adj_4249), 
            .I3(GND_net), .O(n29954));   // verilog/motorControl.v(36[10:25])
    defparam i24862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3395_4_lut (.I0(GND_net), .I1(n6803[1]), .I2(n256_adj_3995), 
            .I3(n22850), .O(n6790[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_5 (.CI(n22851), .I0(n6803[2]), .I1(n329_adj_3994), 
            .CO(n22852));
    SB_LUT4 add_3395_5_lut (.I0(GND_net), .I1(n6803[2]), .I2(n329_adj_3994), 
            .I3(n22851), .O(n6790[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_6 (.CI(n22852), .I0(n6803[3]), .I1(n402_adj_3992), 
            .CO(n22853));
    SB_LUT4 add_3395_6_lut (.I0(GND_net), .I1(n6803[3]), .I2(n402_adj_3992), 
            .I3(n22852), .O(n6790[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_7 (.CI(n22853), .I0(n6803[4]), .I1(n475_adj_3991), 
            .CO(n22854));
    SB_LUT4 i25037_4_lut (.I0(n29954), .I1(n30083), .I2(n35_adj_4253), 
            .I3(n29385), .O(n30129));   // verilog/motorControl.v(36[10:25])
    defparam i25037_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3395_7_lut (.I0(GND_net), .I1(n6803[4]), .I2(n475_adj_3991), 
            .I3(n22853), .O(n6790[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_8 (.CI(n22854), .I0(n6803[5]), .I1(n548_adj_3990), 
            .CO(n22855));
    SB_LUT4 add_3395_8_lut (.I0(GND_net), .I1(n6803[5]), .I2(n548_adj_3990), 
            .I3(n22854), .O(n6790[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_9 (.CI(n22855), .I0(n6803[6]), .I1(n621_adj_3989), 
            .CO(n22856));
    SB_LUT4 add_3395_9_lut (.I0(GND_net), .I1(n6803[6]), .I2(n621_adj_3989), 
            .I3(n22855), .O(n6790[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_10 (.CI(n22856), .I0(n6803[7]), .I1(n694_adj_3988), 
            .CO(n22857));
    SB_LUT4 add_3395_10_lut (.I0(GND_net), .I1(n6803[7]), .I2(n694_adj_3988), 
            .I3(n22856), .O(n6790[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3395_11 (.CI(n22857), .I0(n6803[8]), .I1(n767_adj_3987), 
            .CO(n22858));
    SB_LUT4 i25038_3_lut (.I0(n30129), .I1(duty[18]), .I2(n37_adj_4247), 
            .I3(GND_net), .O(n30130));   // verilog/motorControl.v(36[10:25])
    defparam i25038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25018_3_lut (.I0(n30130), .I1(duty[19]), .I2(n39_adj_4245), 
            .I3(GND_net), .O(n30110));   // verilog/motorControl.v(36[10:25])
    defparam i25018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24286_4_lut (.I0(n43_adj_4250), .I1(n41_adj_4244), .I2(n39_adj_4245), 
            .I3(n30070), .O(n29376));
    defparam i24286_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i24940_4_lut (.I0(n29952), .I1(n29873), .I2(n45_adj_4246), 
            .I3(n29374), .O(n30032));   // verilog/motorControl.v(36[10:25])
    defparam i24940_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i25008_3_lut (.I0(n30110), .I1(duty[20]), .I2(n41_adj_4244), 
            .I3(GND_net), .O(n40_adj_4271));   // verilog/motorControl.v(36[10:25])
    defparam i25008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24942_4_lut (.I0(n40_adj_4271), .I1(n30032), .I2(n45_adj_4246), 
            .I3(n29376), .O(n30034));   // verilog/motorControl.v(36[10:25])
    defparam i24942_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24943_3_lut (.I0(n30034), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3515));   // verilog/motorControl.v(36[10:25])
    defparam i24943_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3491[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4107));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3395_11_lut (.I0(GND_net), .I1(n6803[8]), .I2(n767_adj_3987), 
            .I3(n22857), .O(n6790[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3395_12_lut (.I0(GND_net), .I1(n6803[9]), .I2(n840_adj_3986), 
            .I3(n22858), .O(n6790[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3395_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_2 (.CI(GND_net), .I0(n44_adj_3985), .I1(n113_adj_3984), 
            .CO(n22859));
    SB_LUT4 add_3396_2_lut (.I0(GND_net), .I1(n44_adj_3985), .I2(n113_adj_3984), 
            .I3(GND_net), .O(n6803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_3 (.CI(n22859), .I0(n6815[0]), .I1(n186_adj_3983), 
            .CO(n22860));
    SB_LUT4 add_3396_3_lut (.I0(GND_net), .I1(n6815[0]), .I2(n186_adj_3983), 
            .I3(n22859), .O(n6803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_4 (.CI(n22860), .I0(n6815[1]), .I1(n259_adj_3982), 
            .CO(n22861));
    SB_LUT4 add_3396_4_lut (.I0(GND_net), .I1(n6815[1]), .I2(n259_adj_3982), 
            .I3(n22860), .O(n6803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_5 (.CI(n22861), .I0(n6815[2]), .I1(n332_adj_3981), 
            .CO(n22862));
    SB_LUT4 add_3396_5_lut (.I0(GND_net), .I1(n6815[2]), .I2(n332_adj_3981), 
            .I3(n22861), .O(n6803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[16]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3396_6 (.CI(n22862), .I0(n6815[3]), .I1(n405_adj_3980), 
            .CO(n22863));
    SB_LUT4 add_3396_6_lut (.I0(GND_net), .I1(n6815[3]), .I2(n405_adj_3980), 
            .I3(n22862), .O(n6803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_7 (.CI(n22863), .I0(n6815[4]), .I1(n478_adj_3979), 
            .CO(n22864));
    SB_LUT4 add_3396_7_lut (.I0(GND_net), .I1(n6815[4]), .I2(n478_adj_3979), 
            .I3(n22863), .O(n6803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_8 (.CI(n22864), .I0(n6815[5]), .I1(n551_adj_3978), 
            .CO(n22865));
    SB_LUT4 add_563_25_lut (.I0(GND_net), .I1(n2529[23]), .I2(n2554[23]), 
            .I3(n22036), .O(duty_23__N_3491[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_24_lut (.I0(GND_net), .I1(n2529[22]), .I2(n2554[22]), 
            .I3(n22035), .O(duty_23__N_3491[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_24 (.CI(n22035), .I0(n2529[22]), .I1(n2554[22]), 
            .CO(n22036));
    SB_LUT4 add_563_23_lut (.I0(GND_net), .I1(n2529[21]), .I2(n2554[21]), 
            .I3(n22034), .O(duty_23__N_3491[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_23 (.CI(n22034), .I0(n2529[21]), .I1(n2554[21]), 
            .CO(n22035));
    SB_LUT4 add_3396_8_lut (.I0(GND_net), .I1(n6815[5]), .I2(n551_adj_3978), 
            .I3(n22864), .O(n6803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_9 (.CI(n22865), .I0(n6815[6]), .I1(n624_adj_3976), 
            .CO(n22866));
    SB_LUT4 add_3396_9_lut (.I0(GND_net), .I1(n6815[6]), .I2(n624_adj_3976), 
            .I3(n22865), .O(n6803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3396_10 (.CI(n22866), .I0(n6815[7]), .I1(n697_adj_3974), 
            .CO(n22867));
    SB_LUT4 add_3396_10_lut (.I0(GND_net), .I1(n6815[7]), .I2(n697_adj_3974), 
            .I3(n22866), .O(n6803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3396_11_lut (.I0(GND_net), .I1(n6815[8]), .I2(n770_adj_3972), 
            .I3(n22867), .O(n6803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3396_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_2 (.CI(GND_net), .I0(n47_adj_3971), .I1(n116_adj_3970), 
            .CO(n22868));
    SB_LUT4 add_3397_2_lut (.I0(GND_net), .I1(n47_adj_3971), .I2(n116_adj_3970), 
            .I3(GND_net), .O(n6815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_3 (.CI(n22868), .I0(n6826[0]), .I1(n189_adj_3969), 
            .CO(n22869));
    SB_LUT4 add_3397_3_lut (.I0(GND_net), .I1(n6826[0]), .I2(n189_adj_3969), 
            .I3(n22868), .O(n6815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_4 (.CI(n22869), .I0(n6826[1]), .I1(n262_adj_3968), 
            .CO(n22870));
    SB_LUT4 add_3397_4_lut (.I0(GND_net), .I1(n6826[1]), .I2(n262_adj_3968), 
            .I3(n22869), .O(n6815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_5 (.CI(n22870), .I0(n6826[2]), .I1(n335_adj_3967), 
            .CO(n22871));
    SB_LUT4 add_3397_5_lut (.I0(GND_net), .I1(n6826[2]), .I2(n335_adj_3967), 
            .I3(n22870), .O(n6815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_6 (.CI(n22871), .I0(n6826[3]), .I1(n408_adj_3966), 
            .CO(n22872));
    SB_LUT4 add_3397_6_lut (.I0(GND_net), .I1(n6826[3]), .I2(n408_adj_3966), 
            .I3(n22871), .O(n6815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_7 (.CI(n22872), .I0(n6826[4]), .I1(n481_adj_3965), 
            .CO(n22873));
    SB_LUT4 add_3397_10_lut (.I0(GND_net), .I1(n6826[7]), .I2(n700_adj_3964), 
            .I3(n22875), .O(n6815[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3397_7_lut (.I0(GND_net), .I1(n6826[4]), .I2(n481_adj_3965), 
            .I3(n22872), .O(n6815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[17]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_22_lut (.I0(GND_net), .I1(n2529[20]), .I2(n2554[20]), 
            .I3(n22033), .O(duty_23__N_3491[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \PID_CONTROLLER.integral_1128__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[0]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4106));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_22 (.CI(n22033), .I0(n2529[20]), .I1(n2554[20]), 
            .CO(n22034));
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4104));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_21_lut (.I0(GND_net), .I1(n2529[19]), .I2(n2554[19]), 
            .I3(n22032), .O(duty_23__N_3491[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_21 (.CI(n22032), .I0(n2529[19]), .I1(n2554[19]), 
            .CO(n22033));
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4100));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4099));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3937));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4084));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4082));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4077));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4073));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4069));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4068));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4063));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 setpoint_23__I_0_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), 
            .I2(motor_state[23]), .I3(n22083), .O(\PID_CONTROLLER.err_23__N_3392 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_20_lut (.I0(GND_net), .I1(n2529[18]), .I2(n2554[18]), 
            .I3(n22031), .O(duty_23__N_3491[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4057));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4056));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_20 (.CI(n22031), .I0(n2529[18]), .I1(n2554[18]), 
            .CO(n22032));
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4053));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4052));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4051));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n2554[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14631_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n2529[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam i14631_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256), 
            .I3(GND_net), .O(n2554[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[18]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[19]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4025));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4009));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4007));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4277));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256), 
            .I3(GND_net), .O(n2554[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_563_19_lut (.I0(GND_net), .I1(n2529[17]), .I2(n2554[17]), 
            .I3(n22030), .O(duty_23__N_3491[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_3936));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4278));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4005));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4003));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[20]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 setpoint_23__I_0_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), 
            .I2(motor_state[22]), .I3(n22082), .O(\PID_CONTROLLER.err_23__N_3392 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_24 (.CI(n22082), .I0(setpoint[22]), 
            .I1(motor_state[22]), .CO(n22083));
    SB_CARRY add_563_19 (.CI(n22030), .I0(n2529[17]), .I1(n2554[17]), 
            .CO(n22031));
    SB_LUT4 add_563_18_lut (.I0(GND_net), .I1(n2529[16]), .I2(n2554[16]), 
            .I3(n22029), .O(duty_23__N_3491[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_561_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256), 
            .I3(GND_net), .O(n2554[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_563_18 (.CI(n22029), .I0(n2529[16]), .I1(n2554[16]), 
            .CO(n22030));
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[21]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 setpoint_23__I_0_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), 
            .I2(motor_state[21]), .I3(n22081), .O(\PID_CONTROLLER.err_23__N_3392 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_23 (.CI(n22081), .I0(setpoint[21]), 
            .I1(motor_state[21]), .CO(n22082));
    SB_LUT4 setpoint_23__I_0_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), 
            .I2(motor_state[20]), .I3(n22080), .O(\PID_CONTROLLER.err_23__N_3392 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_561_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256), 
            .I3(GND_net), .O(n2554[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_563_17_lut (.I0(GND_net), .I1(n2529[15]), .I2(n2554[15]), 
            .I3(n22028), .O(duty_23__N_3491[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[22]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[23]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_561_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256), 
            .I3(GND_net), .O(n2554[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_561_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256), 
            .I3(GND_net), .O(n2554[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3491[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3491[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3491[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3491[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_3935));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3491[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_3934));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_3933));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3491[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_3932));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_17 (.CI(n22028), .I0(n2529[15]), .I1(n2554[15]), 
            .CO(n22029));
    SB_CARRY setpoint_23__I_0_add_2_22 (.CI(n22080), .I0(setpoint[20]), 
            .I1(motor_state[20]), .CO(n22081));
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3491[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3491[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3491[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3491[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3491[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3491[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3491[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3491[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3491[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3491[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3491[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3491[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3491[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3491[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3491[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24315_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n29405));   // verilog/motorControl.v(36[10:25])
    defparam i24315_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3368[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_4265));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 setpoint_23__I_0_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), 
            .I2(motor_state[19]), .I3(n22079), .O(\PID_CONTROLLER.err_23__N_3392 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_21 (.CI(n22079), .I0(setpoint[19]), 
            .I1(motor_state[19]), .CO(n22080));
    SB_LUT4 setpoint_23__I_0_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), 
            .I2(motor_state[18]), .I3(n22078), .O(\PID_CONTROLLER.err_23__N_3392 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_16_lut (.I0(GND_net), .I1(n2529[14]), .I2(n2554[14]), 
            .I3(n22027), .O(duty_23__N_3491[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3491[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_561_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256), 
            .I3(GND_net), .O(n2554[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256), 
            .I3(GND_net), .O(n2554[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_563_16 (.CI(n22027), .I0(n2529[14]), .I1(n2554[14]), 
            .CO(n22028));
    SB_LUT4 add_563_15_lut (.I0(GND_net), .I1(n2529[13]), .I2(n2554[13]), 
            .I3(n22026), .O(duty_23__N_3491[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_20 (.CI(n22078), .I0(setpoint[18]), 
            .I1(motor_state[18]), .CO(n22079));
    SB_CARRY add_563_15 (.CI(n22026), .I0(n2529[13]), .I1(n2554[13]), 
            .CO(n22027));
    SB_LUT4 i17982_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_4282), .I3(n7157[1]), .O(n6_adj_4228));   // verilog/motorControl.v(34[26:37])
    defparam i17982_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 setpoint_23__I_0_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), 
            .I2(motor_state[17]), .I3(n22077), .O(\PID_CONTROLLER.err_23__N_3392 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_14_lut (.I0(GND_net), .I1(n2529[12]), .I2(n2554[12]), 
            .I3(n22025), .O(duty_23__N_3491[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n7157[1]), .I3(n4_adj_4282), .O(n7150[2]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_CARRY setpoint_23__I_0_add_2_19 (.CI(n22077), .I0(setpoint[17]), 
            .I1(motor_state[17]), .CO(n22078));
    SB_CARRY add_563_14 (.CI(n22025), .I0(n2529[12]), .I1(n2554[12]), 
            .CO(n22026));
    SB_LUT4 i2_3_lut_4_lut_adj_1471 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n7157[0]), .I3(n21775), .O(n7150[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1471.LUT_INIT = 16'h8778;
    SB_LUT4 setpoint_23__I_0_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), 
            .I2(motor_state[16]), .I3(n22076), .O(\PID_CONTROLLER.err_23__N_3392 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_13_lut (.I0(GND_net), .I1(n2529[11]), .I2(n2554[11]), 
            .I3(n22024), .O(duty_23__N_3491[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_18 (.CI(n22076), .I0(setpoint[16]), 
            .I1(motor_state[16]), .CO(n22077));
    SB_CARRY add_563_13 (.CI(n22024), .I0(n2529[11]), .I1(n2554[11]), 
            .CO(n22025));
    SB_LUT4 i17974_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n21775), .I3(n7157[0]), .O(n4_adj_4282));   // verilog/motorControl.v(34[26:37])
    defparam i17974_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 setpoint_23__I_0_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), 
            .I2(motor_state[15]), .I3(n22075), .O(\PID_CONTROLLER.err_23__N_3392 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17963_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n21775));   // verilog/motorControl.v(34[26:37])
    defparam i17963_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i17961_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n7150[0]));   // verilog/motorControl.v(34[26:37])
    defparam i17961_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_561_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256), 
            .I3(GND_net), .O(n2554[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_561_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256), 
            .I3(GND_net), .O(n2554[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_3931));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18044_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n21852), .I3(n7168[0]), .O(n4_adj_4242));   // verilog/motorControl.v(34[26:37])
    defparam i18044_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_563_12_lut (.I0(GND_net), .I1(n2529[10]), .I2(n2554[10]), 
            .I3(n22023), .O(duty_23__N_3491[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_17 (.CI(n22075), .I0(setpoint[15]), 
            .I1(motor_state[15]), .CO(n22076));
    SB_LUT4 i2_3_lut_4_lut_adj_1472 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n7168[0]), .I3(n21852), .O(n7163[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1472.LUT_INIT = 16'h8778;
    SB_CARRY add_563_12 (.CI(n22023), .I0(n2529[10]), .I1(n2554[10]), 
            .CO(n22024));
    SB_LUT4 i2_3_lut_4_lut_adj_1473 (.I0(n62_adj_4234), .I1(n131_adj_4233), 
            .I2(n7163[0]), .I3(n204_adj_4229), .O(n7157[1]));   // verilog/motorControl.v(34[26:37])
    defparam i2_3_lut_4_lut_adj_1473.LUT_INIT = 16'h8778;
    SB_LUT4 i18013_3_lut_4_lut (.I0(n62_adj_4234), .I1(n131_adj_4233), .I2(n204_adj_4229), 
            .I3(n7163[0]), .O(n4_adj_4235));   // verilog/motorControl.v(34[26:37])
    defparam i18013_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_563_11_lut (.I0(GND_net), .I1(n2529[9]), .I2(n2554[9]), 
            .I3(n22022), .O(duty_23__N_3491[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18033_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n21852));   // verilog/motorControl.v(34[26:37])
    defparam i18033_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 setpoint_23__I_0_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), 
            .I2(motor_state[14]), .I3(n22074), .O(\PID_CONTROLLER.err_23__N_3392 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18031_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n7163[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18031_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY setpoint_23__I_0_add_2_16 (.CI(n22074), .I0(setpoint[14]), 
            .I1(motor_state[14]), .CO(n22075));
    SB_LUT4 setpoint_23__I_0_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), 
            .I2(motor_state[13]), .I3(n22073), .O(\PID_CONTROLLER.err_23__N_3392 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_15 (.CI(n22073), .I0(setpoint[13]), 
            .I1(motor_state[13]), .CO(n22074));
    SB_CARRY add_563_11 (.CI(n22022), .I0(n2529[9]), .I1(n2554[9]), .CO(n22023));
    SB_LUT4 add_563_10_lut (.I0(GND_net), .I1(n2529[8]), .I2(n2554[8]), 
            .I3(n22021), .O(duty_23__N_3491[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 setpoint_23__I_0_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), 
            .I2(motor_state[12]), .I3(n22072), .O(\PID_CONTROLLER.err_23__N_3392 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_14 (.CI(n22072), .I0(setpoint[12]), 
            .I1(motor_state[12]), .CO(n22073));
    SB_CARRY add_563_10 (.CI(n22021), .I0(n2529[8]), .I1(n2554[8]), .CO(n22022));
    SB_LUT4 add_563_9_lut (.I0(GND_net), .I1(n2529[7]), .I2(n2554[7]), 
            .I3(n22020), .O(duty_23__N_3491[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_561_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256), 
            .I3(GND_net), .O(n2554[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3368[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 setpoint_23__I_0_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), 
            .I2(motor_state[11]), .I3(n22071), .O(\PID_CONTROLLER.err_23__N_3392 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3368[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3368[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3368[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3368[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3368[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3368[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3368[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3368[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3368[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3368[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3368[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3368[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3368[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3368[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3368[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3368[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3368[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3368[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3368[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3368[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3368[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3392 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_3930));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY setpoint_23__I_0_add_2_13 (.CI(n22071), .I0(setpoint[11]), 
            .I1(motor_state[11]), .CO(n22072));
    SB_CARRY add_563_9 (.CI(n22020), .I0(n2529[7]), .I1(n2554[7]), .CO(n22021));
    SB_LUT4 setpoint_23__I_0_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), 
            .I2(motor_state[10]), .I3(n22070), .O(\PID_CONTROLLER.err_23__N_3392 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_3929));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_561_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256), 
            .I3(GND_net), .O(n2554[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_563_8_lut (.I0(GND_net), .I1(n2529[6]), .I2(n2554[6]), 
            .I3(n22019), .O(duty_23__N_3491[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_3928));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3927));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_8 (.CI(n22019), .I0(n2529[6]), .I1(n2554[6]), .CO(n22020));
    SB_CARRY setpoint_23__I_0_add_2_12 (.CI(n22070), .I0(setpoint[10]), 
            .I1(motor_state[10]), .CO(n22071));
    SB_LUT4 setpoint_23__I_0_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), 
            .I2(motor_state[9]), .I3(n22069), .O(\PID_CONTROLLER.err_23__N_3392 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_7_lut (.I0(GND_net), .I1(n2529[5]), .I2(n2554[5]), 
            .I3(n22018), .O(duty_23__N_3491[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1_adj_4311[23]), 
            .I3(n22207), .O(n47_adj_4049)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY setpoint_23__I_0_add_2_11 (.CI(n22069), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n22070));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[22]), 
            .I3(n22206), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_7 (.CI(n22018), .I0(n2529[5]), .I1(n2554[5]), .CO(n22019));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n22206), .I0(GND_net), .I1(n1_adj_4311[22]), 
            .CO(n22207));
    SB_LUT4 mux_561_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256), 
            .I3(GND_net), .O(n2554[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 setpoint_23__I_0_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), 
            .I2(motor_state[8]), .I3(n22068), .O(\PID_CONTROLLER.err_23__N_3392 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_6_lut (.I0(GND_net), .I1(n2529[4]), .I2(n2554[4]), 
            .I3(n22017), .O(duty_23__N_3491[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_10 (.CI(n22068), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n22069));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[21]), 
            .I3(n22205), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 setpoint_23__I_0_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), 
            .I2(motor_state[7]), .I3(n22067), .O(\PID_CONTROLLER.err_23__N_3392 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_6 (.CI(n22017), .I0(n2529[4]), .I1(n2554[4]), .CO(n22018));
    SB_CARRY setpoint_23__I_0_add_2_9 (.CI(n22067), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n22068));
    SB_LUT4 add_563_5_lut (.I0(GND_net), .I1(n2529[3]), .I2(n2554[3]), 
            .I3(n22016), .O(duty_23__N_3491[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n22205), .I0(GND_net), .I1(n1_adj_4311[21]), 
            .CO(n22206));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[20]), 
            .I3(n22204), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_561_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256), 
            .I3(GND_net), .O(n2554[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_561_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_3993));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_563_5 (.CI(n22016), .I0(n2529[3]), .I1(n2554[3]), .CO(n22017));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n22204), .I0(GND_net), .I1(n1_adj_4311[20]), 
            .CO(n22205));
    SB_LUT4 setpoint_23__I_0_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), 
            .I2(motor_state[6]), .I3(n22066), .O(\PID_CONTROLLER.err_23__N_3392 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3397_9_lut (.I0(GND_net), .I1(n6826[6]), .I2(n627_adj_4278), 
            .I3(n22874), .O(n6815[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_8 (.CI(n22066), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n22067));
    SB_CARRY add_3397_9 (.CI(n22874), .I0(n6826[6]), .I1(n627_adj_4278), 
            .CO(n22875));
    SB_LUT4 add_563_4_lut (.I0(GND_net), .I1(n2529[2]), .I2(n2554[2]), 
            .I3(n22015), .O(duty_23__N_3491[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3397_8_lut (.I0(GND_net), .I1(n6826[5]), .I2(n554_adj_4277), 
            .I3(n22873), .O(n6815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3397_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3397_8 (.CI(n22873), .I0(n6826[5]), .I1(n554_adj_4277), 
            .CO(n22874));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[19]), 
            .I3(n22203), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n22203), .I0(GND_net), .I1(n1_adj_4311[19]), 
            .CO(n22204));
    SB_CARRY add_563_4 (.CI(n22015), .I0(n2529[2]), .I1(n2554[2]), .CO(n22016));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[18]), 
            .I3(n22202), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3491[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3515), .I3(GND_net), .O(duty_23__N_3368[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_563_3_lut (.I0(GND_net), .I1(n2529[1]), .I2(n2554[1]), 
            .I3(n22014), .O(duty_23__N_3491[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_563_3 (.CI(n22014), .I0(n2529[1]), .I1(n2554[1]), .CO(n22015));
    SB_LUT4 setpoint_23__I_0_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), 
            .I2(motor_state[5]), .I3(n22065), .O(\PID_CONTROLLER.err_23__N_3392 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_7 (.CI(n22065), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n22066));
    SB_LUT4 setpoint_23__I_0_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), 
            .I2(motor_state[4]), .I3(n22064), .O(\PID_CONTROLLER.err_23__N_3392 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_563_2_lut (.I0(GND_net), .I1(n2529[0]), .I2(n2554[0]), 
            .I3(GND_net), .O(duty_23__N_3491[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_6 (.CI(n22064), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n22065));
    SB_CARRY unary_minus_16_add_3_20 (.CI(n22202), .I0(GND_net), .I1(n1_adj_4311[18]), 
            .CO(n22203));
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_3977));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 setpoint_23__I_0_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), 
            .I2(motor_state[3]), .I3(n22063), .O(\PID_CONTROLLER.err_23__N_3392 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[17]), 
            .I3(n22201), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n22201), .I0(GND_net), .I1(n1_adj_4311[17]), 
            .CO(n22202));
    SB_CARRY add_563_2 (.CI(GND_net), .I0(n2529[0]), .I1(n2554[0]), .CO(n22014));
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY setpoint_23__I_0_add_2_5 (.CI(n22063), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n22064));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[16]), 
            .I3(n22200), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 setpoint_23__I_0_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), 
            .I2(motor_state[2]), .I3(n22062), .O(\PID_CONTROLLER.err_23__N_3392 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n22200), .I0(GND_net), .I1(n1_adj_4311[16]), 
            .CO(n22201));
    SB_CARRY setpoint_23__I_0_add_2_4 (.CI(n22062), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n22063));
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3926));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[15]), 
            .I3(n22199), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n22199), .I0(GND_net), .I1(n1_adj_4311[15]), 
            .CO(n22200));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n22424), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n22423), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_24  (.CI(n22423), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n22424));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n22422), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_23  (.CI(n22422), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n22423));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n22421), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_22  (.CI(n22421), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n22422));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n22420), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_21  (.CI(n22420), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n22421));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n22419), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_20  (.CI(n22419), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n22420));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n22418), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_19  (.CI(n22418), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n22419));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n22417), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3925));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_3924));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_3923));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_3973));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_18  (.CI(n22417), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n22418));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n22416), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_3963));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_4268));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24282_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n29372));
    defparam i24282_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_4266));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_4270));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24293_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n29383));
    defparam i24293_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_4263));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i18000_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n7157[0]));   // verilog/motorControl.v(34[26:37])
    defparam i18000_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_3922));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_17  (.CI(n22416), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n22417));
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_3921));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n22415), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_16  (.CI(n22415), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n22416));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n22414), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_15  (.CI(n22414), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n22415));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n22413), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 i17878_2_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\Kp[1] ), .I3(\PID_CONTROLLER.err [19]), .O(n6860[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17878_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24248_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n29338));
    defparam i24248_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_14  (.CI(n22413), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n22414));
    SB_LUT4 i24258_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n29348));
    defparam i24258_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n22412), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_13  (.CI(n22412), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n22413));
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[0]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 setpoint_23__I_0_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), 
            .I2(motor_state[1]), .I3(n22061), .O(\PID_CONTROLLER.err_23__N_3392 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[1]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n22411), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_12  (.CI(n22411), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n22412));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n22410), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_11  (.CI(n22410), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n22411));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n22409), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[2]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[14]), 
            .I3(n22198), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[3]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_10  (.CI(n22409), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n22410));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n22408), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_9  (.CI(n22408), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n22409));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n22407), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY setpoint_23__I_0_add_2_3 (.CI(n22061), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n22062));
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[4]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_8  (.CI(n22407), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n22408));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n22198), .I0(GND_net), .I1(n1_adj_4311[14]), 
            .CO(n22199));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n22406), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_7  (.CI(n22406), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n22407));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n22405), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 setpoint_23__I_0_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), 
            .I2(motor_state[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3392 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam setpoint_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_6  (.CI(n22405), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n22406));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[13]), 
            .I3(n22197), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n22404), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[5]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_5  (.CI(n22404), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n22405));
    SB_CARRY unary_minus_16_add_3_15 (.CI(n22197), .I0(GND_net), .I1(n1_adj_4311[13]), 
            .CO(n22198));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n22403), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_4  (.CI(n22403), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n22404));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n22402), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_3  (.CI(n22402), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n22403));
    SB_LUT4 \PID_CONTROLLER.integral_1128_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1128_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1128_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n22402));
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[6]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[7]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[8]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[9]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[10]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_3920));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[11]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_3962));   // verilog/motorControl.v(34[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[12]), 
            .I3(n22196), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n22196), .I0(GND_net), .I1(n1_adj_4311[12]), 
            .CO(n22197));
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE \PID_CONTROLLER.integral_1128__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[1]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[2]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[3]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[4]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[5]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[6]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[7]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[8]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[9]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[10]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[11]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[12]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[13]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[14]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[15]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[16]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[17]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[18]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[19]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[20]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[21]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[22]));   // verilog/motorControl.v(32[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1128__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3464 ), .D(n28[23]));   // verilog/motorControl.v(32[21:33])
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3913));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17860_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4309), .I3(n6860[1]), .O(n6_adj_4080));   // verilog/motorControl.v(34[17:23])
    defparam i17860_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[11]), 
            .I3(n22195), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1474 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n6860[1]), .I3(n4_adj_4309), .O(n6853[2]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1474.LUT_INIT = 16'h8778;
    SB_CARRY setpoint_23__I_0_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n22061));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n22195), .I0(GND_net), .I1(n1_adj_4311[11]), 
            .CO(n22196));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[10]), 
            .I3(n22194), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n6860[0]), .I3(n21643), .O(n6853[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h8778;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n22194), .I0(GND_net), .I1(n1_adj_4311[10]), 
            .CO(n22195));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[9]), 
            .I3(n22193), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n22193), .I0(GND_net), .I1(n1_adj_4311[9]), 
            .CO(n22194));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[8]), 
            .I3(n22192), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n22192), .I0(GND_net), .I1(n1_adj_4311[8]), 
            .CO(n22193));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[7]), 
            .I3(n22191), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n22191), .I0(GND_net), .I1(n1_adj_4311[7]), 
            .CO(n22192));
    SB_LUT4 i17852_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n21643), .I3(n6860[0]), .O(n4_adj_4309));   // verilog/motorControl.v(34[17:23])
    defparam i17852_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[6]), 
            .I3(n22190), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n22190), .I0(GND_net), .I1(n1_adj_4311[6]), 
            .CO(n22191));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[5]), 
            .I3(n22189), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17839_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n6853[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17839_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n22189), .I0(GND_net), .I1(n1_adj_4311[5]), 
            .CO(n22190));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[4]), 
            .I3(n22188), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n22188), .I0(GND_net), .I1(n1_adj_4311[4]), 
            .CO(n22189));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[3]), 
            .I3(n22187), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17841_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n21643));   // verilog/motorControl.v(34[17:23])
    defparam i17841_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n22187), .I0(GND_net), .I1(n1_adj_4311[3]), 
            .CO(n22188));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[2]), 
            .I3(n22186), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n22186), .I0(GND_net), .I1(n1_adj_4311[2]), 
            .CO(n22187));
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17922_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n21720), .I3(n6871[0]), .O(n4_adj_4091));   // verilog/motorControl.v(34[17:23])
    defparam i17922_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4311[1]), 
            .I3(n22185), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n6871[0]), .I3(n21720), .O(n6866[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h8778;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n22185), .I0(GND_net), .I1(n1_adj_4311[1]), 
            .CO(n22186));
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[12]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1_adj_4311[0]), 
            .I3(VCC_net), .O(n29248)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4311[0]), 
            .CO(n22185));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n22184), .O(\PID_CONTROLLER.integral_23__N_3467 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[13]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1477 (.I0(n62), .I1(n131), .I2(n6866[0]), 
            .I3(n204), .O(n6860[1]));   // verilog/motorControl.v(34[17:23])
    defparam i2_3_lut_4_lut_adj_1477.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n22183), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4311[14]));   // verilog/motorControl.v(39[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n22183), .I0(GND_net), .I1(n1[22]), 
            .CO(n22184));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n22182), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17891_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n6866[0]), 
            .O(n4_adj_4085));   // verilog/motorControl.v(34[17:23])
    defparam i17891_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i17911_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n21720));   // verilog/motorControl.v(34[17:23])
    defparam i17911_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i17909_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n6866[0]));   // verilog/motorControl.v(34[17:23])
    defparam i17909_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i14877_2_lut_2_lut (.I0(n256), .I1(n5022[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2529[23]));   // verilog/motorControl.v(38[19:35])
    defparam i14877_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n22182), .I0(GND_net), .I1(n1[21]), 
            .CO(n22183));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n22181), .O(n41_adj_3918)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n22181), .I0(GND_net), .I1(n1[20]), 
            .CO(n22182));
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_out_frame[19] , n15009, \data_in[1] , clk32MHz, GND_net, 
            \data_out_frame[15] , \data_out_frame[17] , \data_out_frame[20] , 
            \data_out_frame[14] , \data_out_frame[16] , setpoint, n15008, 
            \data_in_frame[3] , \data_out_frame[24] , \data_out_frame[23] , 
            \data_out_frame[11] , \data_out_frame[9] , \data_out_frame[7] , 
            \data_out_frame[13] , n15007, n4167, n10927, \data_out_frame[6] , 
            \data_out_frame[10] , \data_out_frame[12] , \data_out_frame[5] , 
            n4169, \data_out_frame[18] , \data_out_frame[8] , rx_data, 
            n15006, \data_in_frame[1] , n15005, \data_in_frame[2] , 
            n15004, n15003, n15002, \data_in[0] , \data_in_frame[6] , 
            n15001, n15000, n14999, rx_data_ready, n14998, n14997, 
            \data_in_frame[9] , \data_in_frame[10] , n14996, \data_in_frame[5] , 
            \data_out_frame[25] , n123, n63, n13620, \data_in_frame[4] , 
            \data_in_frame[13] , n3303, \FRAME_MATCHER.state_31__N_2508[1] , 
            n52, n7480, \FRAME_MATCHER.state_31__N_2380[2] , \FRAME_MATCHER.state_31__N_2540[2] , 
            \data_in[3] , \data_in[2] , \data_in_frame[12] , \data_in_frame[8] , 
            n63_adj_3, \data_in_frame[11] , n13615, n26676, n13618, 
            n6, n14994, IntegralLimit, n14993, tx_active, n14992, 
            DE_c, LED_c, n14991, n14990, n14989, n14988, n14987, 
            n14986, n14985, n14984, n14983, n14982, n14981, n14980, 
            n14979, n14978, n14977, n14976, n14975, n14974, n14973, 
            n14972, n7330, n30906, n30907, n15436, PWMLimit, n15435, 
            n15434, n15433, n15432, n15431, n15430, n15429, n15428, 
            n15427, n15426, n15425, n15424, n15423, n15422, n15421, 
            n15420, n15419, n15418, n15417, n15416, n15415, n15414, 
            n15413, control_mode, n15412, n15411, n15410, n15409, 
            n15408, n15407, n15231, neopxl_color, n15230, n15229, 
            n15228, n15227, n15226, n15225, n15224, n15223, n15222, 
            n15221, n15220, n15219, n15218, n15217, n15216, n15215, 
            n15214, n15213, n15212, n15211, n15210, n15209, n15208, 
            n15207, n15206, n15205, n15204, n15203, n15202, n15201, 
            n15200, n15199, n15198, n15197, n15196, n15195, n15194, 
            n15193, n15192, n15191, n15190, n15189, n15188, n15187, 
            n15186, n15185, n15184, n15183, n15182, n15181, n15180, 
            n15179, n15178, n15177, n15176, n15175, n15174, n15173, 
            n15172, n15171, n15170, n15169, n15168, n15167, n15166, 
            n15165, n15164, n15163, n15162, n15161, n15160, n15159, 
            n15158, n15157, n15156, n15155, n15154, n15153, n15152, 
            n15151, n15150, n15149, n15148, n15147, n15146, n15145, 
            n15144, n15143, n15142, n15141, n15140, n15139, n15138, 
            n15137, n15136, n15135, n15134, n15133, n15132, n15131, 
            n15130, n15129, n15128, n15127, n15126, n15125, n15124, 
            n15123, n15122, n15121, n15120, n15119, n15118, n15117, 
            n15116, n15115, n15114, n15113, n15112, n15111, n15110, 
            n15109, n15108, n15107, n15106, n15105, n15104, n15103, 
            n14953, n14952, n14950, n15102, n15101, n15100, n15099, 
            n15098, n15097, n15096, n14949, \Ki[0] , n14948, \Kp[0] , 
            n14947, n15095, n15094, n15093, n15092, n15091, n15090, 
            n15089, n15088, n15087, n15086, n15085, n15084, n15083, 
            n15082, n15081, n15080, n15079, n15078, n15077, n15076, 
            n15075, n15074, n15073, n15072, n15071, n15070, n15069, 
            n15068, n15067, n15066, n14941, n15065, n15064, n15063, 
            n15062, n15061, n15060, n15059, n15058, n15057, n15056, 
            \Ki[15] , n15055, \Ki[14] , n15054, \Ki[13] , n15053, 
            \Ki[12] , n15052, \Ki[11] , n15051, \Ki[10] , n15050, 
            \Ki[9] , n15049, \Ki[8] , n15048, \Ki[7] , n15047, \Ki[6] , 
            n15046, \Ki[5] , n15045, \Ki[4] , n15044, \Ki[3] , n15043, 
            \Ki[2] , n15042, \Ki[1] , n15041, \Kp[15] , n15040, 
            \Kp[14] , n15039, \Kp[13] , n15038, \Kp[12] , n15037, 
            \Kp[11] , n15036, \Kp[10] , n15035, \Kp[9] , n15034, 
            \Kp[8] , n15033, \Kp[7] , n15032, \Kp[6] , n15031, \Kp[5] , 
            n15030, \Kp[4] , n15029, \Kp[3] , n15028, \Kp[2] , n15027, 
            \Kp[1] , n15026, n15025, n15024, n15023, n15022, n15021, 
            n15020, n15019, n15018, n15017, n15016, n15015, n15014, 
            n15013, n15012, n15011, n15010, n26810, n26830, \r_Bit_Index[0] , 
            r_SM_Main, tx_o, \r_SM_Main_2__N_3333[1] , VCC_net, n14961, 
            n4, n14955, n30923, n7410, tx_enable, n14794, n14921, 
            r_SM_Main_adj_11, r_Rx_Data, RX_N_2, n14995, \r_SM_Main_2__N_3262[2] , 
            \r_Bit_Index[0]_adj_7 , n13657, n4_adj_8, n4_adj_9, n13652, 
            n4_adj_10, n25972, n14971, n14970, n14969, n14968, n14957, 
            n14964, n25630, n18503, n14946, n14945) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_out_frame[19] ;
    input n15009;
    output [7:0]\data_in[1] ;
    input clk32MHz;
    input GND_net;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[16] ;
    output [23:0]setpoint;
    input n15008;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[13] ;
    input n15007;
    output n4167;
    output n10927;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[5] ;
    output n4169;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]rx_data;
    input n15006;
    output [7:0]\data_in_frame[1] ;
    input n15005;
    output [7:0]\data_in_frame[2] ;
    input n15004;
    input n15003;
    input n15002;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in_frame[6] ;
    input n15001;
    input n15000;
    input n14999;
    output rx_data_ready;
    input n14998;
    input n14997;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[10] ;
    input n14996;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_out_frame[25] ;
    output n123;
    output n63;
    output n13620;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[13] ;
    output n3303;
    output \FRAME_MATCHER.state_31__N_2508[1] ;
    output n52;
    output n7480;
    output \FRAME_MATCHER.state_31__N_2380[2] ;
    output \FRAME_MATCHER.state_31__N_2540[2] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[8] ;
    output n63_adj_3;
    output [7:0]\data_in_frame[11] ;
    output n13615;
    output n26676;
    output n13618;
    output n6;
    input n14994;
    output [23:0]IntegralLimit;
    input n14993;
    output tx_active;
    input n14992;
    output DE_c;
    output LED_c;
    input n14991;
    input n14990;
    input n14989;
    input n14988;
    input n14987;
    input n14986;
    input n14985;
    input n14984;
    input n14983;
    input n14982;
    input n14981;
    input n14980;
    input n14979;
    input n14978;
    input n14977;
    input n14976;
    input n14975;
    input n14974;
    input n14973;
    input n14972;
    output n7330;
    input n30906;
    input n30907;
    input n15436;
    output [23:0]PWMLimit;
    input n15435;
    input n15434;
    input n15433;
    input n15432;
    input n15431;
    input n15430;
    input n15429;
    input n15428;
    input n15427;
    input n15426;
    input n15425;
    input n15424;
    input n15423;
    input n15422;
    input n15421;
    input n15420;
    input n15419;
    input n15418;
    input n15417;
    input n15416;
    input n15415;
    input n15414;
    input n15413;
    output [7:0]control_mode;
    input n15412;
    input n15411;
    input n15410;
    input n15409;
    input n15408;
    input n15407;
    input n15231;
    output [23:0]neopxl_color;
    input n15230;
    input n15229;
    input n15228;
    input n15227;
    input n15226;
    input n15225;
    input n15224;
    input n15223;
    input n15222;
    input n15221;
    input n15220;
    input n15219;
    input n15218;
    input n15217;
    input n15216;
    input n15215;
    input n15214;
    input n15213;
    input n15212;
    input n15211;
    input n15210;
    input n15209;
    input n15208;
    input n15207;
    input n15206;
    input n15205;
    input n15204;
    input n15203;
    input n15202;
    input n15201;
    input n15200;
    input n15199;
    input n15198;
    input n15197;
    input n15196;
    input n15195;
    input n15194;
    input n15193;
    input n15192;
    input n15191;
    input n15190;
    input n15189;
    input n15188;
    input n15187;
    input n15186;
    input n15185;
    input n15184;
    input n15183;
    input n15182;
    input n15181;
    input n15180;
    input n15179;
    input n15178;
    input n15177;
    input n15176;
    input n15175;
    input n15174;
    input n15173;
    input n15172;
    input n15171;
    input n15170;
    input n15169;
    input n15168;
    input n15167;
    input n15166;
    input n15165;
    input n15164;
    input n15163;
    input n15162;
    input n15161;
    input n15160;
    input n15159;
    input n15158;
    input n15157;
    input n15156;
    input n15155;
    input n15154;
    input n15153;
    input n15152;
    input n15151;
    input n15150;
    input n15149;
    input n15148;
    input n15147;
    input n15146;
    input n15145;
    input n15144;
    input n15143;
    input n15142;
    input n15141;
    input n15140;
    input n15139;
    input n15138;
    input n15137;
    input n15136;
    input n15135;
    input n15134;
    input n15133;
    input n15132;
    input n15131;
    input n15130;
    input n15129;
    input n15128;
    input n15127;
    input n15126;
    input n15125;
    input n15124;
    input n15123;
    input n15122;
    input n15121;
    input n15120;
    input n15119;
    input n15118;
    input n15117;
    input n15116;
    input n15115;
    input n15114;
    input n15113;
    input n15112;
    input n15111;
    input n15110;
    input n15109;
    input n15108;
    input n15107;
    input n15106;
    input n15105;
    input n15104;
    input n15103;
    input n14953;
    input n14952;
    input n14950;
    input n15102;
    input n15101;
    input n15100;
    input n15099;
    input n15098;
    input n15097;
    input n15096;
    input n14949;
    output \Ki[0] ;
    input n14948;
    output \Kp[0] ;
    input n14947;
    input n15095;
    input n15094;
    input n15093;
    input n15092;
    input n15091;
    input n15090;
    input n15089;
    input n15088;
    input n15087;
    input n15086;
    input n15085;
    input n15084;
    input n15083;
    input n15082;
    input n15081;
    input n15080;
    input n15079;
    input n15078;
    input n15077;
    input n15076;
    input n15075;
    input n15074;
    input n15073;
    input n15072;
    input n15071;
    input n15070;
    input n15069;
    input n15068;
    input n15067;
    input n15066;
    input n14941;
    input n15065;
    input n15064;
    input n15063;
    input n15062;
    input n15061;
    input n15060;
    input n15059;
    input n15058;
    input n15057;
    input n15056;
    output \Ki[15] ;
    input n15055;
    output \Ki[14] ;
    input n15054;
    output \Ki[13] ;
    input n15053;
    output \Ki[12] ;
    input n15052;
    output \Ki[11] ;
    input n15051;
    output \Ki[10] ;
    input n15050;
    output \Ki[9] ;
    input n15049;
    output \Ki[8] ;
    input n15048;
    output \Ki[7] ;
    input n15047;
    output \Ki[6] ;
    input n15046;
    output \Ki[5] ;
    input n15045;
    output \Ki[4] ;
    input n15044;
    output \Ki[3] ;
    input n15043;
    output \Ki[2] ;
    input n15042;
    output \Ki[1] ;
    input n15041;
    output \Kp[15] ;
    input n15040;
    output \Kp[14] ;
    input n15039;
    output \Kp[13] ;
    input n15038;
    output \Kp[12] ;
    input n15037;
    output \Kp[11] ;
    input n15036;
    output \Kp[10] ;
    input n15035;
    output \Kp[9] ;
    input n15034;
    output \Kp[8] ;
    input n15033;
    output \Kp[7] ;
    input n15032;
    output \Kp[6] ;
    input n15031;
    output \Kp[5] ;
    input n15030;
    output \Kp[4] ;
    input n15029;
    output \Kp[3] ;
    input n15028;
    output \Kp[2] ;
    input n15027;
    output \Kp[1] ;
    input n15026;
    input n15025;
    input n15024;
    input n15023;
    input n15022;
    input n15021;
    input n15020;
    input n15019;
    input n15018;
    input n15017;
    input n15016;
    input n15015;
    input n15014;
    input n15013;
    input n15012;
    input n15011;
    input n15010;
    output n26810;
    output n26830;
    output \r_Bit_Index[0] ;
    output [2:0]r_SM_Main;
    output tx_o;
    output \r_SM_Main_2__N_3333[1] ;
    input VCC_net;
    input n14961;
    output n4;
    input n14955;
    input n30923;
    output n7410;
    output tx_enable;
    output n14794;
    output n14921;
    output [2:0]r_SM_Main_adj_11;
    output r_Rx_Data;
    input RX_N_2;
    input n14995;
    output \r_SM_Main_2__N_3262[2] ;
    output \r_Bit_Index[0]_adj_7 ;
    output n13657;
    output n4_adj_8;
    output n4_adj_9;
    output n13652;
    output n4_adj_10;
    input n25972;
    input n14971;
    input n14970;
    input n14969;
    input n14968;
    input n14957;
    input n14964;
    input n25630;
    output n18503;
    input n14946;
    input n14945;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n15, n20, n24669, n28011, n26271, n26272, n13844, n1445, 
        n6_c, n24594, n26326, n21941;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n21942, n2, n21940, n1656, n4_c, n26245, n3964, n14715, 
        n2_adj_3581, n3;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n3963, n3965, n24639, n26417, n12, n26545, n27697, n26214, 
        n26123, n29, n27, n23, n24, n30, n13779, n26490, n11797, 
        n16, n14211, n26602, n26542, n17;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n28321, n13814, n13, n25896, n23731, n26378, n13611, 
        n26050, n14243, n26511, n24649, n6_adj_3582, n13703, n24641, 
        n21466;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    wire [31:0]\FRAME_MATCHER.state_31__N_2444 ;
    
    wire n6_adj_3583, n26396, n26999, n26608, n26161, n13347, n10, 
        n26650, n26242, n26475, n14412, n22, n26144, n26435, n20_adj_3584, 
        n13828, n16_adj_3585, n26599, n24_adj_3586, n23741, n26632, 
        n26313, n14, n10_adj_3587, n14111, n24531, n24609, n26300, 
        n24600, n14216, n26348, n26478, n26141, n6_adj_3588, n11807, 
        n26104, n13610, n1, n26158, n26469, n14668, n12_adj_3589, 
        n14453, n26596, n26100, n23785, n24582, n7, n24607, n26307, 
        n24550, n14056, n26340, n13308, n6_adj_3590, n28156, n13294, 
        n10_adj_3591, n26180, n26536, n26487, n2_adj_3592, n21939, 
        n26623, n12033, n26508, Kp_23__N_1053, n14_adj_3593, n14527, 
        n21969;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n21970, n2_adj_3594, n21938, n26037, n14511, n18, n13756, 
        n16_adj_3595, n20_adj_3596;
    wire [7:0]n8825;
    
    wire n21968, n26151, n21967, n14034, n16_adj_3597, n13707, n1427, 
        n17_adj_3598, n2_adj_3599, Kp_23__N_1030, n10_adj_3600, n3_adj_3601, 
        n24618, n14237, n18_adj_3602, n23759, n26186, n20_adj_3603, 
        n16_adj_3604, n26481, n14219, n23749, n14185, n6_adj_3605, 
        n8, n26126, n26107, n14_adj_3606, n26113, n15_adj_3607, 
        n23733, n26197, n18978, n25997;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n15293, n14680, n26472, n6_adj_3608, n26647, n6_adj_3609, 
        n1180, n26364, n15294, n26611, n1265, n26575, n26148, 
        n24584, n1563, n26438, n26096, n14314, n26046, n13906, 
        n12_adj_3610, n14116, n26084, n26463, n26590, n6_adj_3611, 
        n26070, n18565, n14763, n14737, n13651, n14863;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n3987, n3986, n3985, n3984, n3983, n3982, n3981, n3980;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n3979, n3978, n3977, n3976, n3975, n3974, n3973, n3972, 
        n3971, n3970, n3969, n3968, n3967, n3966, n6_adj_3612, 
        n5, n29161, n7_adj_3613, n30487, n30475, n14_adj_3614, n30511, 
        n29218, n16_adj_3615, n17_adj_3616, n29223, n29222, n16_adj_3617, 
        n17_adj_3618, n29220, n29219, n6_adj_3619, n5_adj_3620, n7_adj_3621, 
        n8_adj_3622, n15279, n2_adj_3623, n21937, n30469, n30457, 
        n14_adj_3624, n30517, n29221, n6_adj_3625, n5_adj_3626, n7_adj_3627, 
        n30463, n30499, n14_adj_3628, n30277, n29224, n15280, n15281, 
        n13892, n26074, n6_adj_3629, n15282, n15283, n15284, n15285, 
        n6_adj_3630, n5_adj_3631, n7_adj_3632, n30451, n30349, n14_adj_3633, 
        n30283, n29227, n29573, n5_adj_3634, n7_adj_3635, n30445, 
        n30547, n14_adj_3636, n30289, n29230, n2_adj_3637, n21936;
    wire [0:0]n2813;
    wire [2:0]r_SM_Main_2__N_3336;
    
    wire n26785, tx_transmit_N_3233, n29567, n5_adj_3638, n7_adj_3639, 
        n30439, n30565, n14_adj_3640, n30325, n29233, n15286, n6_adj_3641, 
        \FRAME_MATCHER.rx_data_ready_prev , n25396, n25624, n5_adj_3642, 
        n7_adj_3643, n30433, n30415, n14_adj_3644, n30331, n29237, 
        n6_adj_3645, n5_adj_3646, n7_adj_3647, n161, n30493, n30403, 
        n14_adj_3648, n30343, n29240, n14082, n27069, n23743, n26202, 
        n26040, n13937, n10_adj_3649, n28341, n26557, n26167, n26131, 
        n13972, n13_adj_3650, n11166, n7_adj_3651, n8_adj_3652, n27074, 
        n26220, n6_adj_3653, Kp_23__N_810, n14491, n26408, n26566, 
        n26563, n26280, n13665, n8_adj_3654, n15271, n14_adj_3655, 
        n26429, n26411, n24656, n26189, n26502, n15_adj_3656, n26384, 
        n15272, n13369, n13747, n26304, n13919, n23804, n2406, 
        n27864, n2400, n27830, n62, n53, n8634, n2_adj_3657, n21966, 
        n11123, n3_adj_3658, n25434, n25432, n25430, n2_adj_3659, 
        n21965, n15273, n15274, n2_adj_3660, n21964, n25428, n26484, 
        n6_adj_3661, n14297, n15275, n7_adj_3662, n25426, n15276, 
        n7_adj_3663, n25424, n25382, n25388, n15277, n2_adj_3664, 
        n21963, n18428, n7_adj_3665, n7_adj_3666, n15278, n7_adj_3667, 
        n7_adj_3668, n2_adj_3669, n21962, n25422, n25420, n2_adj_3670, 
        n21961, n8_adj_3671, n15263, n25418, n25416, n2_adj_3672, 
        n21960, n25414, n15264, n25412, n25408, n18424, n18426, 
        n7_adj_3673, n15265, n7_adj_3674, n18422, n2_adj_3675, n21959, 
        n8_adj_3676, n25404, n184, n44, n25264, n18938, n8_adj_3677, 
        n18936, n2_adj_3678, n21958, n18934, n15266, n15267;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n26211, n25894, n19125, n25892, n6_adj_3679, n18435, n25990, 
        n15268, n15269, n16455, n2_adj_3680, n21957, n15270, n13686, 
        n14075, n8_adj_3681, n26514, n26881, n24654, n2_adj_3682, 
        n21956, n8_adj_3683, n15255, n15256, n15257, n10_adj_3684, 
        n25438, n25478, n25480, n15258, n25442, n25482, n25484, 
        n25486, n25508, n15259, n25384, n771, n4452, n25490, n25492, 
        n25494, n15260, n25496, n15261, n25498, n25500, n25502, 
        n26605, n14_adj_3685, n9, n13606, n10_adj_3686, n15262, 
        n26587, n13867, n26620, n13641, n18_adj_3687, n16_adj_3688, 
        n20_adj_3689, n13496, n28377, n9_adj_3690, n13628, n16_adj_3691, 
        n28383, n16_adj_3692, n17_adj_3693, n28365, n4040, n21, 
        n20_adj_3694, n24_adj_3695, n5_adj_3696, n14328, n17_adj_3697, 
        n21_adj_3698, n26498, n13852, n26034, n14_adj_3699, n8_adj_3700, 
        n28118, n14420, n20_adj_3701, n23686, n24_adj_3702, n23717, 
        n10_adj_3703, Kp_23__N_698, n27195, n26370, Kp_23__N_708, 
        n13621, n10_adj_3705, n18939, n2254;
    wire [31:0]\FRAME_MATCHER.state_31__N_2380 ;
    
    wire n14017, n13808, n13988, n26629, n6_adj_3706, n26333, n26028, 
        n26059, n23761, n8_adj_3707, n13625, n44_adj_3708, n42, 
        n43, n41, n40, n39, n13508, n26155, n2_adj_3709, n21955, 
        n50, n45, n13505, n26134, n14396, n8_adj_3710, n10_adj_3711, 
        n13794, n12_adj_3712, n8_adj_3713, n26297, n26120, n16_adj_3714, 
        n28307, n5_adj_3715, n11, n13616, n8_adj_3716, n15247, n26678, 
        n27507, n28267, n15248, Kp_23__N_888, n14153, n26387, n10_adj_3717, 
        n13950, n26223, n26505, n23702, n26402, n13_adj_3718, n14380, 
        n26205, n2_adj_3720, n21954, n26283, n15249, Kp_23__N_656, 
        n6_adj_3721, n26087, n12058;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n26457, n26361, n26554, n26584, n26323, n26031, n26432, 
        n10_adj_3722, n26656, n26208, n26581, n14308, n23700, n26274, 
        n26653, Kp_23__N_713, n12_adj_3723, Kp_23__N_1041, Kp_23__N_1256, 
        n12_adj_3724;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n26117, n26183, n24689, n10_adj_3725, n13877, n23768, n26056, 
        n24652, n10_adj_3726, n26420, n26016, n19121, n6_adj_3727, 
        n806, n15250, n18966, n2_adj_3728, n21953, n26688, n26217, 
        n7_adj_3729, n6_adj_3730, n18983, n8_adj_3731, n15251, n15252, 
        n15253, n15254, n26093, n2_adj_3732, n21952, n6_adj_3733, 
        n16_adj_3734, n17_adj_3735, n29242, n29241, n16_adj_3736, 
        n17_adj_3737, n29239, n29238, n16_adj_3738, n17_adj_3739, 
        n29236, n10_adj_3740, n29235, n24696, n14_adj_3741, n16_adj_3742, 
        n26043, n14_adj_3743, n17_adj_3744, n18_adj_3745, n10_adj_3746, 
        n26110, n29232, n24_adj_3747, n29231, n23692, n22_adj_3748, 
        n16_adj_3749, n17_adj_3750, n29229, n26, n26239, n29228, 
        n25, n13675, n26494, n26527, n10_adj_3751, n6_adj_3752, 
        n24523, n7_adj_3753, n26286, n24578, n10_adj_3754, n14383, 
        n13377, n26330, n24533, n12137, n26336, n6_adj_3755, n24249, 
        n14677, n12_adj_3756, n26289, n13964, n10_adj_3757, n8_adj_3758, 
        n14005, n12_adj_3759, n13788, n26172, n24560, n26175, n26284, 
        n21_adj_3760, n20_adj_3761, n18_adj_3762, n26641, n24_adj_3763, 
        n24566, n18_adj_3764, n30_adj_3765, n28, Kp_23__N_1237, n8_adj_3766, 
        n15239, n29_adj_3767, n27_adj_3768, n20_adj_3769, n26533, 
        n19, n26077, n13391, n21_adj_3770, n14665, n10_adj_3771, 
        n26426, n26460, n23747, n15240, n61, n26659, n26626, n60, 
        n68, n55, n26081, n66, n13723, n26635, n64, n26447, 
        n26441, n65, n26090, n63_adj_3772, n46, n70, Kp_23__N_1218, 
        n69, n73, n75, n26399, n26539, n23770, n26252, n14599, 
        n13873, n6_adj_3773, n26423, n26381, n14130, n30562, n8_adj_3774, 
        n26560, n23706, n30295, n30550, n4_adj_3775;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n30544, n30301, n30538, n30307, n30532, n30313, n30526, 
        n8_adj_3776, n30319, n30520;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n30514, n30508, n30496, n26569, n30490, n26064, n30484, 
        n26053, n12_adj_3777, n14205, n30472, n30466, n30460, n26067, 
        n18_adj_3778, n30454, n10_adj_3779, n30448;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n12_adj_3780, n30442, n16_adj_3781, n30436;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n10_adj_3782, n30430, n26524, n27617, n6_adj_3783, n8_adj_3784, 
        n30412, n27118, n28121, n30400, n30955, n26319, n9_adj_3785, 
        n38, n6_adj_3786, n27002, n30337, n30376, n11_adj_3787, 
        n30361, n30370, n14_adj_3788, n30364, n29670, n12_adj_3789, 
        n18_adj_3790, n30358, n4_adj_3791, n30352, n28125, n30346, 
        n8_adj_3792, n30340, n3_adj_3793, n13751, n2122, n3_adj_3794, 
        n3_adj_3795, n15241, n24544, n24554, n24251, n3_adj_3796, 
        n3_adj_3797, n3_adj_3798, n23772, n3_adj_3799, n15242, n15243, 
        n3_adj_3800, n3_adj_3801, n3_adj_3802, n3_adj_3803, n27514, 
        n3_adj_3804, n3_adj_3805, n3_adj_3806, n3_adj_3807, n10_adj_3808, 
        n3_adj_3809, n3_adj_3810, n3_adj_3811, n3_adj_3812, n3_adj_3813, 
        n3_adj_3814, n3_adj_3815, n3_adj_3816, n3_adj_3817, n2_adj_3818, 
        n3_adj_3819, n2_adj_3820, n3_adj_3821, n2_adj_3822, n3_adj_3823, 
        n2_adj_3824, n3_adj_3825, n2_adj_3826, n3_adj_3827, n2_adj_3828, 
        n3_adj_3829, n2_adj_3830, n3_adj_3831, n2_adj_3832, n2_adj_3833, 
        n2_adj_3834, n27684, n26852, n27278, n26391, n26392, n11578, 
        n26890, n27205, n26972, n25400, n8_adj_3835, n8_adj_3836, 
        n8_adj_3837, n8_adj_3838, n8_adj_3839, n8_adj_3840, n8_adj_3841, 
        n25378, n15244, n15245, n15246, n15399, n15400, n16_adj_3842, 
        n17_adj_3843, n21951, n15401, n29226, n26572, n29225, n15522, 
        n26794, n15402, n15403, n15404, n15405, n15406, n14853, 
        n13_adj_3844, n27660, n21950, n21949, n15391, n15392, n15393, 
        n15394, n15395, n15396, n15397, n15398, n21948, n21947, 
        n15383, n15384, n15385, n15386, n30334, n15387, n15388, 
        n21944, n21945, n15389, n15390, n14951, n15375, n15376, 
        n15377, n21946, n15378, n15379, n15380, n15381, n15382, 
        n15367, n15368, n12_adj_3845, n15232, n15369, n15233, n61_adj_3846, 
        n15370, n26779, n51, n15234, n15235, n15371, n15372, n15_adj_3847, 
        n15373, n15236, n15374, n15359, n15360, n15361, n28339, 
        n15237, n15362, n15363, n15364, n15238, n15365, n30328, 
        n20_adj_3848, n30322, n19_adj_3849, n30316, n27779, n30310, 
        n28357, n30304, n6_adj_3850, n30298, n27142, n30292, n26310, 
        n20_adj_3851, n15366, n25981, n15351, n15352, n15353, n15354, 
        n15355, n15356, n15357, n15358, n18_adj_3852, n21973, n21972, 
        n21943, n15343, n15344, n15345, n194, n15346, n21971, 
        n26638, n15350, n15349, n15348, n15347, n15342, n15341, 
        n15340, n15339, n15338, n15337, n15336, n15335, n15334, 
        n15333, n15332, n15331, n15330, n15329, n15328, n15327, 
        n15326, n15325, n15324, n15323, n15322, n15321, n15320, 
        n15319, n15318, n15317, n15316, n15315, n15314, n15313, 
        n15312, n15311, n15310, n15309, n15308, n15307, n15306, 
        n15305, n15304, n15303, n15302, n15301, n15300, n15299, 
        n15298, n15297, n15296, n15295, n15292, n15291, n15290, 
        n15289, n15288, n15287, n19_adj_3853, n18_adj_3854, n30286, 
        n17_adj_3855, n30280, n30274, n11119, n11125, n13805, n28_adj_3856, 
        n18_adj_3857, n17_adj_3858, n19_adj_3859, n6_adj_3860, n26644, 
        n27904, n26265, n24558, n26393, n14487, n24046, n24615, 
        n26390, n26551, n26268, n14_adj_3861, n24598, n26351, n26343, 
        n6_adj_3862, n24180, n6_adj_3863, n26262, n11926, n26228, 
        n1927, n23696, n26248, n14_adj_3864, n9_adj_3865, n24546, 
        n26255, n26530, n26578, n18_adj_3866, n16_adj_3867, n20_adj_3868, 
        n27626, n23715, n25_adj_3869, n24574, n30_adj_3870, n26234, 
        n23989, n24580, n28_adj_3871, n26025, n29_adj_3872, n27_adj_3873, 
        n26259, n42_adj_3874, n40_adj_3875, n41_adj_3876, n14171, 
        n39_adj_3877, n43_adj_3878, n48, n47, n18_adj_3879, n26405, 
        n20_adj_3880, n13_adj_3881, n7_adj_3882, n14524, n13933, n14337, 
        n26989, n16_adj_3883, n13767, n17_adj_3884, n10_adj_3885, 
        n27058, n14_adj_3886, n4_adj_3887, n24142, n12_adj_3888, n26349, 
        n7_adj_3889, n21_adj_3890, n20_adj_3891, n24_adj_3892, n18_adj_3893;
    
    SB_LUT4 i10_4_lut (.I0(n15), .I1(n20), .I2(n24669), .I3(\data_out_frame[19] [6]), 
            .O(n28011));
    defparam i10_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n15009));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(n28011), .I1(n26271), .I2(GND_net), .I3(GND_net), 
            .O(n26272));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[15] [5]), .I1(n13844), .I2(n1445), 
            .I3(n6_c), .O(n24594));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_836 (.I0(\data_out_frame[17] [4]), .I1(n24594), 
            .I2(GND_net), .I3(GND_net), .O(n24669));
    defparam i1_2_lut_adj_836.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_837 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26326));
    defparam i1_2_lut_adj_837.LUT_INIT = 16'h6666;
    SB_CARRY add_43_8 (.CI(n21941), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n21942));
    SB_LUT4 add_43_7_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n21940), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[17] [1]), 
            .I2(n4_c), .I3(\data_out_frame[16] [7]), .O(n26245));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n14715), .D(n3964));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3581), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n15008));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_985_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n3963), .I3(GND_net), .O(n3965));
    defparam mux_985_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(n24639), .I1(n26417), .I2(\data_out_frame[24] [1]), 
            .I3(\data_out_frame[19] [7]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[24] [2]), .I1(n12), .I2(n26545), 
            .I3(\data_out_frame[23] [7]), .O(n27697));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[11] [2]), .I1(n26214), .I2(\data_out_frame[9] [0]), 
            .I3(\data_out_frame[7] [0]), .O(n26123));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n29), .I1(n27), .I2(n23), .I3(n24), .O(n30));
    defparam i15_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_838 (.I0(n13779), .I1(\data_out_frame[9] [1]), 
            .I2(n26490), .I3(n11797), .O(n16));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_838.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n14211), .I1(\data_out_frame[15] [4]), .I2(n26602), 
            .I3(n26542), .O(n17));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23234_2_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28321));
    defparam i23234_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n26123), .I2(n16), .I3(\data_out_frame[13] [3]), 
            .O(n13814));   // verilog/coms.v(85[17:28])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n15007));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_839 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [2]), .O(n13));
    defparam i5_4_lut_adj_839.LUT_INIT = 16'h0800;
    SB_LUT4 i7_4_lut_adj_840 (.I0(n13), .I1(\data_in_frame[0] [7]), .I2(n28321), 
            .I3(\data_in_frame[0] [3]), .O(n25896));
    defparam i7_4_lut_adj_840.LUT_INIT = 16'h0008;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[16] [6]), .I1(n23731), .I2(\data_out_frame[17] [0]), 
            .I3(GND_net), .O(n26378));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_841 (.I0(n30), .I1(n25896), .I2(n13611), .I3(GND_net), 
            .O(n4167));
    defparam i2_3_lut_adj_841.LUT_INIT = 16'h0808;
    SB_LUT4 i2_3_lut_adj_842 (.I0(n26050), .I1(\data_out_frame[19] [6]), 
            .I2(n14243), .I3(GND_net), .O(n26511));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_842.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[19] [2]), .I1(n24649), .I2(n6_adj_3582), 
            .I3(n13703), .O(n24641));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_843 (.I0(n21466), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state_31__N_2444 [3]), .I3(n6_adj_3583), 
            .O(n10927));
    defparam i4_4_lut_adj_843.LUT_INIT = 16'h1000;
    SB_LUT4 i3_4_lut_adj_844 (.I0(\data_out_frame[23] [6]), .I1(n26396), 
            .I2(\data_out_frame[24] [0]), .I3(\data_out_frame[24] [1]), 
            .O(n26999));
    defparam i3_4_lut_adj_844.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_845 (.I0(\data_out_frame[11] [1]), .I1(n26608), 
            .I2(n26161), .I3(n13347), .O(n10));
    defparam i4_4_lut_adj_845.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26542));
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_847 (.I0(n26650), .I1(n26242), .I2(n26475), .I3(n14412), 
            .O(n22));
    defparam i9_4_lut_adj_847.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n26144), .I1(n26435), .I2(\data_out_frame[15] [1]), 
            .I3(GND_net), .O(n20_adj_3584));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(n13828), .I1(n22), .I2(n16_adj_3585), .I3(n26599), 
            .O(n24_adj_3586));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[13] [0]), .I1(n24_adj_3586), 
            .I2(n20_adj_3584), .I3(\data_out_frame[14] [7]), .O(n23741));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_848 (.I0(n26632), .I1(\data_out_frame[10] [6]), 
            .I2(n26313), .I3(\data_out_frame[12] [7]), .O(n14));
    defparam i6_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_849 (.I0(\data_out_frame[15] [3]), .I1(n14), .I2(n10_adj_3587), 
            .I3(n14111), .O(n24531));
    defparam i7_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_850 (.I0(n24531), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26417));
    defparam i1_2_lut_adj_850.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_851 (.I0(\data_out_frame[17] [3]), .I1(n23741), 
            .I2(GND_net), .I3(GND_net), .O(n24609));
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_852 (.I0(\data_out_frame[14] [5]), .I1(n26300), 
            .I2(GND_net), .I3(GND_net), .O(n24600));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_853 (.I0(\data_out_frame[12] [4]), .I1(n14216), 
            .I2(GND_net), .I3(GND_net), .O(n26348));
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_854 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26478));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_855 (.I0(n14211), .I1(n26141), .I2(\data_out_frame[9] [1]), 
            .I3(\data_out_frame[7] [1]), .O(n1445));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_856 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[6] [6]), .I3(n6_adj_3588), .O(n11807));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_857 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26104));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n13844));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_859 (.I0(n13610), .I1(n25896), .I2(n1), .I3(GND_net), 
            .O(n4169));
    defparam i2_3_lut_adj_859.LUT_INIT = 16'h0404;
    SB_LUT4 i5_4_lut_adj_860 (.I0(n26158), .I1(n26469), .I2(n14668), .I3(n26144), 
            .O(n12_adj_3589));
    defparam i5_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_861 (.I0(n14453), .I1(n12_adj_3589), .I2(n26596), 
            .I3(n26100), .O(n23785));
    defparam i6_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_out_frame[16] [7]), .I1(n23785), 
            .I2(GND_net), .I3(GND_net), .O(n24582));
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_863 (.I0(n7), .I1(n24600), .I2(\data_out_frame[19] [1]), 
            .I3(n24607), .O(n26307));
    defparam i4_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_864 (.I0(n24550), .I1(n26307), .I2(n24582), .I3(GND_net), 
            .O(n14056));
    defparam i2_3_lut_adj_864.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_865 (.I0(\data_out_frame[24] [0]), .I1(n14056), 
            .I2(\data_out_frame[23] [7]), .I3(GND_net), .O(n26340));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_865.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_866 (.I0(\data_out_frame[23] [5]), .I1(\data_out_frame[19] [5]), 
            .I2(n13308), .I3(n6_adj_3590), .O(n28156));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_CARRY add_43_7 (.CI(n21940), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n21941));
    SB_LUT4 i1_2_lut_adj_867 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26214));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_868 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14453));
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_869 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n13779));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_870 (.I0(n13294), .I1(\data_out_frame[12] [5]), 
            .I2(n14111), .I3(\data_out_frame[12] [6]), .O(n10_adj_3591));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n26180), .I1(n10_adj_3591), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n26144));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_871 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n26632));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_871.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_872 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26536));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_872.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_873 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26487));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_6_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n21939), .O(n2_adj_3592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_874 (.I0(n26623), .I1(n12033), .I2(n26508), .I3(Kp_23__N_1053), 
            .O(n14_adj_3593));
    defparam i6_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_875 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14527));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_875.LUT_INIT = 16'h6666;
    SB_CARRY add_3971_5 (.CI(n21969), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n21970));
    SB_CARRY add_43_6 (.CI(n21939), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n21940));
    SB_LUT4 add_43_5_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n21938), .O(n2_adj_3594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_876 (.I0(n14527), .I1(\data_out_frame[8] [3]), 
            .I2(n26037), .I3(n14511), .O(n18));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_876.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[8] [4]), .I1(n13756), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_3595));   // verilog/coms.v(85[17:28])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_43_5 (.CI(n21938), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n21939));
    SB_LUT4 i9_4_lut_adj_877 (.I0(\data_out_frame[7] [7]), .I1(n18), .I2(\data_out_frame[8] [2]), 
            .I3(n26487), .O(n20_adj_3596));   // verilog/coms.v(85[17:28])
    defparam i9_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n21968), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_878 (.I0(n26151), .I1(n20_adj_3596), .I2(n16_adj_3595), 
            .I3(\data_out_frame[8] [6]), .O(n13347));   // verilog/coms.v(85[17:28])
    defparam i10_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_4 (.CI(n21968), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n21969));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n21967), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_879 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14034));
    defparam i1_2_lut_adj_879.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_880 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [1]), 
            .I2(n14034), .I3(n26608), .O(n16_adj_3597));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_881 (.I0(n13707), .I1(n1427), .I2(\data_out_frame[8] [5]), 
            .I3(n26536), .O(n17_adj_3598));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_882 (.I0(n17_adj_3598), .I1(\data_out_frame[9] [2]), 
            .I2(n16_adj_3597), .I3(\data_out_frame[9] [1]), .O(n26650));   // verilog/coms.v(85[17:28])
    defparam i9_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_8_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n21941), .O(n2_adj_3599)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_883 (.I0(Kp_23__N_1030), .I1(n14_adj_3593), .I2(n10_adj_3600), 
            .I3(n3_adj_3601), .O(n24618));
    defparam i7_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_884 (.I0(\data_out_frame[10] [4]), .I1(n14237), 
            .I2(n26602), .I3(\data_out_frame[11] [5]), .O(n18_adj_3602));
    defparam i7_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_885 (.I0(n23759), .I1(n18_adj_3602), .I2(n26186), 
            .I3(n26650), .O(n20_adj_3603));
    defparam i9_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_886 (.I0(n26632), .I1(n20_adj_3603), .I2(n16_adj_3604), 
            .I3(n26481), .O(n13294));
    defparam i10_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_887 (.I0(n14219), .I1(n26144), .I2(GND_net), 
            .I3(GND_net), .O(n23749));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_888 (.I0(\data_out_frame[12] [3]), .I1(n14185), 
            .I2(\data_out_frame[12] [0]), .I3(\data_out_frame[12] [7]), 
            .O(n26180));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_889 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(n26435), .I3(n6_adj_3605), .O(n14216));
    defparam i4_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_890 (.I0(\data_out_frame[15] [0]), .I1(n23749), 
            .I2(n8), .I3(n13294), .O(n23731));
    defparam i1_4_lut_adj_890.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26126));
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_892 (.I0(n14211), .I1(n11797), .I2(n26107), .I3(GND_net), 
            .O(n14_adj_3606));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_893 (.I0(n26475), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(n26113), .O(n15_adj_3607));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_893.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_3607), .I1(\data_out_frame[6] [1]), .I2(n14_adj_3606), 
            .I3(\data_out_frame[10] [5]), .O(n14243));   // verilog/coms.v(85[17:28])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_894 (.I0(n23733), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26197));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14237));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_LUT4 i639_2_lut (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1427));   // verilog/coms.v(71[16:27])
    defparam i639_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_896 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26151));
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_LUT4 i11462_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n15293));
    defparam i11462_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_897 (.I0(\data_out_frame[10] [3]), .I1(n14680), 
            .I2(n26472), .I3(n6_adj_3608), .O(n14219));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_out_frame[7] [4]), .I1(n26647), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3609));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_899 (.I0(\data_out_frame[12] [3]), .I1(n1180), 
            .I2(\data_out_frame[12] [2]), .I3(n6_adj_3609), .O(n26364));
    defparam i4_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26161));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i11463_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n15294));
    defparam i11463_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_901 (.I0(\data_out_frame[6] [2]), .I1(n26611), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n1265));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_901.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(n1265), .I3(\data_out_frame[6] [0]), .O(n14680));
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_903 (.I0(n14680), .I1(n13828), .I2(\data_out_frame[9] [7]), 
            .I3(n14511), .O(n26481));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_out_frame[10] [1]), .I1(n26481), 
            .I2(GND_net), .I3(GND_net), .O(n23759));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_out_frame[5] [2]), .I1(n26575), 
            .I2(GND_net), .I3(GND_net), .O(n26148));
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14185));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_907 (.I0(n14185), .I1(n26148), .I2(n23759), .I3(GND_net), 
            .O(n24584));
    defparam i2_3_lut_adj_907.LUT_INIT = 16'h9696;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(71[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_908 (.I0(n1563), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[12] [0]), .O(n26599));
    defparam i3_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\data_out_frame[7] [5]), .I1(n26599), 
            .I2(GND_net), .I3(GND_net), .O(n26438));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i392_2_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1180));   // verilog/coms.v(74[16:27])
    defparam i392_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_910 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n13828));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_911 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26096));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n15006));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_912 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14314));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_out_frame[9] [5]), .I1(n13828), 
            .I2(GND_net), .I3(GND_net), .O(n13707));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_914 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26046));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_915 (.I0(n13707), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[9] [6]), .I3(n14314), .O(n26575));
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_916 (.I0(\data_out_frame[12] [1]), .I1(n26575), 
            .I2(n13906), .I3(n26046), .O(n12_adj_3610));
    defparam i5_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_917 (.I0(n1180), .I1(n12_adj_3610), .I2(\data_out_frame[14] [2]), 
            .I3(n26438), .O(n14116));
    defparam i6_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_918 (.I0(n26300), .I1(n26364), .I2(GND_net), 
            .I3(GND_net), .O(n24649));
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_919 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26084));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n13703));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_921 (.I0(n26463), .I1(n26084), .I2(n26590), .I3(n6_adj_3611), 
            .O(n26070));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n18565), .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n14763));
    defparam i3_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i11032_2_lut (.I0(n14737), .I1(n13651), .I2(GND_net), .I3(GND_net), 
            .O(n14863));   // verilog/coms.v(127[12] 300[6])
    defparam i11032_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_985_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n3963), .I3(GND_net), .O(n3987));
    defparam mux_985_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n3963), .I3(GND_net), .O(n3986));
    defparam mux_985_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n3963), .I3(GND_net), .O(n3985));
    defparam mux_985_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n3963), .I3(GND_net), .O(n3984));
    defparam mux_985_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n3963), .I3(GND_net), .O(n3983));
    defparam mux_985_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n3963), .I3(GND_net), .O(n3982));
    defparam mux_985_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n3963), .I3(GND_net), .O(n3981));
    defparam mux_985_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n15005));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_985_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n3963), .I3(GND_net), .O(n3980));
    defparam mux_985_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n3963), .I3(GND_net), .O(n3979));
    defparam mux_985_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n3963), .I3(GND_net), .O(n3978));
    defparam mux_985_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n3963), .I3(GND_net), .O(n3977));
    defparam mux_985_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n3963), .I3(GND_net), .O(n3976));
    defparam mux_985_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n3963), .I3(GND_net), .O(n3975));
    defparam mux_985_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n3963), .I3(GND_net), .O(n3974));
    defparam mux_985_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n3963), .I3(GND_net), .O(n3973));
    defparam mux_985_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n3963), .I3(GND_net), .O(n3972));
    defparam mux_985_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n3963), .I3(GND_net), .O(n3971));
    defparam mux_985_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n3963), .I3(GND_net), .O(n3970));
    defparam mux_985_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n15004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n15003));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_985_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n3963), .I3(GND_net), .O(n3969));
    defparam mux_985_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n15002));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_985_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n3963), .I3(GND_net), .O(n3968));
    defparam mux_985_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n3963), .I3(GND_net), .O(n3967));
    defparam mux_985_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_985_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n3963), .I3(GND_net), .O(n3966));
    defparam mux_985_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i6_3_lut (.I0(\data_out_frame[5] [1]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3612));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut (.I0(n5), .I1(n6_adj_3612), 
            .I2(n29161), .I3(GND_net), .O(n7_adj_3613));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1536544_i1_3_lut (.I0(n30487), .I1(n30475), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3614));
    defparam i1536544_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24507_2_lut (.I0(n30511), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29218));
    defparam i24507_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3615));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3616));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24495_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29223));
    defparam i24495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24497_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29222));
    defparam i24497_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3617));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3618));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24499_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29220));
    defparam i24499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24502_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29219));
    defparam i24502_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3619));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3620));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_adj_3620), 
            .I1(n6_adj_3619), .I2(n29161), .I3(GND_net), .O(n7_adj_3621));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11448_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n15279));
    defparam i11448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_4_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n21937), .O(n2_adj_3623)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1537147_i1_3_lut (.I0(n30469), .I1(n30457), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3624));
    defparam i1537147_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24501_2_lut (.I0(n30517), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29221));
    defparam i24501_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3625));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3626));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_3626), 
            .I1(n6_adj_3625), .I2(n29161), .I3(GND_net), .O(n7_adj_3627));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1537750_i1_3_lut (.I0(n30463), .I1(n30499), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3628));
    defparam i1537750_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24496_2_lut (.I0(n30277), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29224));
    defparam i24496_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n15001));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11449_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n15280));
    defparam i11449_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11450_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n15281));
    defparam i11450_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_922 (.I0(n13892), .I1(n26074), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3629));
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h6666;
    SB_LUT4 i11451_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n15282));
    defparam i11451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11452_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n15283));
    defparam i11452_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11453_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n15284));
    defparam i11453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11454_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n15285));
    defparam i11454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n15000));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3630));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3631));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_3631), 
            .I1(n6_adj_3630), .I2(n29161), .I3(GND_net), .O(n7_adj_3632));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1538353_i1_3_lut (.I0(n30451), .I1(n30349), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3633));
    defparam i1538353_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24492_2_lut (.I0(n30283), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29227));
    defparam i24492_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n29573));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n14999));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3634));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_3634), 
            .I1(byte_transmit_counter[0]), .I2(n29161), .I3(n29573), .O(n7_adj_3635));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1538956_i1_3_lut (.I0(n30445), .I1(n30547), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3636));
    defparam i1538956_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24487_2_lut (.I0(n30289), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29230));
    defparam i24487_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_4 (.CI(n21937), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n21938));
    SB_CARRY add_3971_3 (.CI(n21967), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n21968));
    SB_LUT4 add_43_3_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n21936), .O(n2_adj_3637)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3336[0]), .C(clk32MHz), 
            .D(n2813[0]), .R(n26785));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3233), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_3 (.CI(n21936), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n21937));
    SB_LUT4 i24477_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29567));   // verilog/coms.v(106[34:55])
    defparam i24477_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3638));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_3638), 
            .I1(n29567), .I2(n29161), .I3(byte_transmit_counter[0]), .O(n7_adj_3639));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1539559_i1_3_lut (.I0(n30439), .I1(n30565), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3640));
    defparam i1539559_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24484_2_lut (.I0(n30325), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29233));
    defparam i24484_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11455_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n15286));
    defparam i11455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23449_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n29161));   // verilog/coms.v(106[34:55])
    defparam i23449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i6_3_lut (.I0(\data_out_frame[5] [7]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n6_adj_3641));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
            .D(n25396), .S(n25624));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3642));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut (.I0(n5_adj_3642), 
            .I1(n6_adj_3641), .I2(n29161), .I3(GND_net), .O(n7_adj_3643));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1540162_i1_3_lut (.I0(n30433), .I1(n30415), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3644));
    defparam i1540162_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24479_2_lut (.I0(n30331), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29237));
    defparam i24479_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n6_adj_3645));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hb0bc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3646));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n14998));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_4_lut (.I0(n5_adj_3646), 
            .I1(n6_adj_3645), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n7_adj_3647));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 add_43_2_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_3581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n21936));
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3233), 
            .CO(n21967));
    SB_LUT4 i1541368_i1_3_lut (.I0(n30493), .I1(n30403), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_3648));
    defparam i1541368_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24472_2_lut (.I0(n30343), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n29240));
    defparam i24472_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n14997));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_923 (.I0(\data_in_frame[9] [0]), .I1(n14082), .I2(n24618), 
            .I3(n6_adj_3629), .O(n27069));
    defparam i4_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_924 (.I0(n27069), .I1(n24618), .I2(GND_net), 
            .I3(GND_net), .O(n23743));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_925 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [1]), .I3(n26202), .O(n26074));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_926 (.I0(n26040), .I1(\data_in_frame[1] [7]), .I2(n13937), 
            .I3(\data_in_frame[0] [3]), .O(n10_adj_3649));   // verilog/coms.v(166[9:87])
    defparam i4_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_LUT4 i23253_2_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28341));
    defparam i23253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_927 (.I0(n26557), .I1(n26167), .I2(\data_in_frame[0] [4]), 
            .I3(n26131), .O(n13972));
    defparam i3_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_928 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [0]), .I3(\data_in_frame[0] [6]), .O(n13_adj_3650));
    defparam i5_4_lut_adj_928.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_929 (.I0(n13_adj_3650), .I1(\data_in_frame[0] [3]), 
            .I2(n28341), .I3(\data_in_frame[0] [2]), .O(n11166));
    defparam i7_4_lut_adj_929.LUT_INIT = 16'hefff;
    SB_LUT4 i2_4_lut_adj_930 (.I0(\data_in_frame[10] [7]), .I1(n14082), 
            .I2(n13972), .I3(n23743), .O(n7_adj_3651));
    defparam i2_4_lut_adj_930.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_931 (.I0(n7_adj_3651), .I1(n13972), .I2(n8_adj_3652), 
            .I3(n26074), .O(n27074));
    defparam i4_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n14996));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_932 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(n26220), .I3(n6_adj_3653), .O(Kp_23__N_810));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [3]), 
            .I2(n14491), .I3(n26408), .O(n15));   // verilog/coms.v(85[17:28])
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [3]), 
            .I2(n14491), .I3(\data_out_frame[18] [0]), .O(n26566));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[11] [4]), .I1(n11807), .I2(n26563), 
            .I3(\data_out_frame[13] [6]), .O(n26280));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n13665));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i11440_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n15271));
    defparam i11440_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_934 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[6] [7]), .I3(GND_net), .O(n14_adj_3655));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_adj_934.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[11] [4]), .I1(n11807), .I2(n14668), 
            .I3(GND_net), .O(n26429));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_935 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[18] [2]), .I3(n26411), .O(n24656));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_936 (.I0(n26189), .I1(\data_in_frame[6] [6]), .I2(\data_in_frame[2] [3]), 
            .I3(n26502), .O(n15_adj_3656));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_937 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n26384));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_LUT4 i11441_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n15272));
    defparam i11441_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_938 (.I0(n13369), .I1(n13747), .I2(\data_out_frame[18] [4]), 
            .I3(\data_out_frame[20] [5]), .O(n26304));
    defparam i2_3_lut_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_939 (.I0(n15_adj_3656), .I1(\data_in_frame[2] [2]), 
            .I2(n14_adj_3655), .I3(\data_in_frame[0] [1]), .O(n13919));   // verilog/coms.v(72[16:27])
    defparam i8_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_940 (.I0(\data_out_frame[25] [5]), .I1(n23804), 
            .I2(\data_out_frame[25] [6]), .I3(n2406), .O(n27864));
    defparam i2_3_lut_4_lut_adj_940.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_941 (.I0(\data_out_frame[25] [5]), .I1(n23804), 
            .I2(n2400), .I3(\data_out_frame[25] [4]), .O(n27830));
    defparam i2_3_lut_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_942 (.I0(n62), .I1(n53), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));
    defparam i1_2_lut_3_lut_adj_942.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_943 (.I0(n62), .I1(n53), .I2(n63), .I3(GND_net), 
            .O(n8634));
    defparam i1_2_lut_3_lut_adj_943.LUT_INIT = 16'h8080;
    SB_LUT4 add_43_33_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n21966), .O(n2_adj_3657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [30]), 
            .I3(n3_adj_3658), .O(n25434));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_944 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [29]), 
            .I3(n3_adj_3658), .O(n25432));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_944.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_945 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [28]), 
            .I3(n3_adj_3658), .O(n25430));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_945.LUT_INIT = 16'hf040;
    SB_LUT4 add_43_32_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n21965), .O(n2_adj_3659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n21965), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n21966));
    SB_LUT4 i11442_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n15273));
    defparam i11442_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11443_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n15274));
    defparam i11443_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_31_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n21964), .O(n2_adj_3660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_946 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [27]), 
            .I3(n3_adj_3658), .O(n25428));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_946.LUT_INIT = 16'hf040;
    SB_LUT4 i4_4_lut_adj_947 (.I0(n13665), .I1(n26484), .I2(Kp_23__N_810), 
            .I3(n6_adj_3661), .O(n14297));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i11444_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n15275));
    defparam i11444_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_948 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [26]), 
            .I3(n3_adj_3658), .O(n7_adj_3662));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_948.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_949 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [25]), 
            .I3(n3_adj_3658), .O(n25426));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_949.LUT_INIT = 16'hf040;
    SB_LUT4 i11445_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n15276));
    defparam i11445_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_950 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [24]), 
            .I3(n3_adj_3658), .O(n7_adj_3663));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_950.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_951 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [23]), 
            .I3(n3_adj_3658), .O(n25424));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_951.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_952 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [22]), 
            .I3(n3_adj_3658), .O(n25382));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_952.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_953 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [21]), 
            .I3(n3_adj_3658), .O(n25388));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_953.LUT_INIT = 16'hf040;
    SB_LUT4 i11446_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n15277));
    defparam i11446_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_31 (.CI(n21964), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n21965));
    SB_LUT4 add_43_30_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n21963), .O(n2_adj_3664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_954 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [20]), 
            .I3(n3_adj_3658), .O(n18428));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_954.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_955 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [19]), 
            .I3(n3_adj_3658), .O(n7_adj_3665));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_955.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_956 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [18]), 
            .I3(n3_adj_3658), .O(n7_adj_3666));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_956.LUT_INIT = 16'hf040;
    SB_LUT4 i11447_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n15278));
    defparam i11447_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_30 (.CI(n21963), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n21964));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_957 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [17]), 
            .I3(n3_adj_3658), .O(n7_adj_3667));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_957.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_958 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [16]), 
            .I3(n3_adj_3658), .O(n7_adj_3668));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_958.LUT_INIT = 16'hf040;
    SB_LUT4 add_43_29_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n21962), .O(n2_adj_3669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_959 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [15]), 
            .I3(n3_adj_3658), .O(n25422));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_959.LUT_INIT = 16'hf040;
    SB_CARRY add_43_29 (.CI(n21962), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n21963));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_960 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [14]), 
            .I3(n3_adj_3658), .O(n25420));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_960.LUT_INIT = 16'hf040;
    SB_LUT4 add_43_28_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n21961), .O(n2_adj_3670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11432_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n15263));
    defparam i11432_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_961 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [13]), 
            .I3(n3_adj_3658), .O(n25418));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_961.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_962 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [12]), 
            .I3(n3_adj_3658), .O(n25416));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_962.LUT_INIT = 16'hf040;
    SB_CARRY add_43_28 (.CI(n21961), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n21962));
    SB_LUT4 add_43_27_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n21960), .O(n2_adj_3672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_27 (.CI(n21960), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n21961));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_963 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [11]), 
            .I3(n3_adj_3658), .O(n25414));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_963.LUT_INIT = 16'hf040;
    SB_LUT4 i11433_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n15264));
    defparam i11433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_964 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [10]), 
            .I3(n3_adj_3658), .O(n25412));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_964.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_965 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [9]), 
            .I3(n3_adj_3658), .O(n25408));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_965.LUT_INIT = 16'hf040;
    SB_LUT4 i14604_2_lut_3_lut_4_lut (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [5]), 
            .I3(n3_adj_3658), .O(n18424));   // verilog/coms.v(254[5:25])
    defparam i14604_2_lut_3_lut_4_lut.LUT_INIT = 16'hf040;
    SB_LUT4 i14605_2_lut_3_lut_4_lut (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [7]), 
            .I3(n3_adj_3658), .O(n18426));   // verilog/coms.v(254[5:25])
    defparam i14605_2_lut_3_lut_4_lut.LUT_INIT = 16'hf040;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_966 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [8]), 
            .I3(n3_adj_3658), .O(n7_adj_3673));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_966.LUT_INIT = 16'hf040;
    SB_LUT4 i11434_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n15265));
    defparam i11434_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_967 (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [6]), 
            .I3(n3_adj_3658), .O(n7_adj_3674));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_967.LUT_INIT = 16'hf040;
    SB_LUT4 i14603_2_lut_3_lut_4_lut (.I0(n13620), .I1(n11123), .I2(\FRAME_MATCHER.state [4]), 
            .I3(n3_adj_3658), .O(n18422));   // verilog/coms.v(254[5:25])
    defparam i14603_2_lut_3_lut_4_lut.LUT_INIT = 16'hf040;
    SB_LUT4 add_43_26_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n21959), .O(n2_adj_3675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_3_lut_4_lut (.I0(n13620), .I1(n11123), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [3]), .O(n25404));   // verilog/coms.v(254[5:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_4_lut_adj_968 (.I0(n184), .I1(n44), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [8]), .O(n25264));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_968.LUT_INIT = 16'hfe00;
    SB_LUT4 i15110_2_lut_4_lut (.I0(n184), .I1(n44), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [7]), .O(n18938));   // verilog/coms.v(115[11:12])
    defparam i15110_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_CARRY add_43_26 (.CI(n21959), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n21960));
    SB_LUT4 i1_2_lut_4_lut_adj_969 (.I0(n184), .I1(n44), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [6]), .O(n8_adj_3677));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_969.LUT_INIT = 16'hfe00;
    SB_LUT4 i15109_2_lut_4_lut (.I0(n184), .I1(n44), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [5]), .O(n18936));   // verilog/coms.v(115[11:12])
    defparam i15109_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 add_43_25_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n21958), .O(n2_adj_3678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15108_2_lut_4_lut (.I0(n184), .I1(n44), .I2(n8_adj_3676), 
            .I3(\FRAME_MATCHER.state [4]), .O(n18934));   // verilog/coms.v(115[11:12])
    defparam i15108_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_970 (.I0(n14297), .I1(n13919), .I2(GND_net), 
            .I3(GND_net), .O(n26623));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i11435_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n15266));
    defparam i11435_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11436_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n15267));
    defparam i11436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_971 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n26211));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_971.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n25894), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n19125), .I3(n25892), .O(n6_adj_3679));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h0001;
    SB_LUT4 i3_4_lut_adj_973 (.I0(n18435), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n25990));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_973.LUT_INIT = 16'hffdf;
    SB_LUT4 i11437_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n15268));
    defparam i11437_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11438_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n15269));
    defparam i11438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_974 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n16455), .I3(n6_adj_3679), .O(n14715));
    defparam i4_4_lut_adj_974.LUT_INIT = 16'h4000;
    SB_CARRY add_43_25 (.CI(n21958), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n21959));
    SB_LUT4 add_43_24_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n21957), .O(n2_adj_3680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11439_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n15270));
    defparam i11439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(n13686), .I3(n14075), .O(n8_adj_3681));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(n26070), .I3(n26514), .O(n26881));
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(\data_out_frame[14] [3]), .I1(n24584), 
            .I2(\data_out_frame[14] [4]), .I3(n26364), .O(n24607));
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_977 (.I0(\data_out_frame[14] [3]), .I1(n24584), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n24654));
    defparam i1_2_lut_3_lut_adj_977.LUT_INIT = 16'h9696;
    SB_CARRY add_43_24 (.CI(n21957), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n21958));
    SB_LUT4 add_43_23_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n21956), .O(n2_adj_3682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11424_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n15255));
    defparam i11424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11425_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n15256));
    defparam i11425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n14737), .D(n8825[0]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11426_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n15257));
    defparam i11426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_978 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [31]), .O(n25438));
    defparam i1_2_lut_4_lut_adj_978.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_979 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [30]), .O(n25478));
    defparam i1_2_lut_4_lut_adj_979.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_980 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [29]), .O(n25480));
    defparam i1_2_lut_4_lut_adj_980.LUT_INIT = 16'hea00;
    SB_LUT4 i11427_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n15258));
    defparam i11427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_981 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [28]), .O(n25442));
    defparam i1_2_lut_4_lut_adj_981.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_982 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [27]), .O(n25482));
    defparam i1_2_lut_4_lut_adj_982.LUT_INIT = 16'hea00;
    SB_LUT4 i2_3_lut_adj_983 (.I0(n63), .I1(n3303), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2508[1] ));
    defparam i2_3_lut_adj_983.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_4_lut_adj_984 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [25]), .O(n25484));
    defparam i1_2_lut_4_lut_adj_984.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_985 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [23]), .O(n25486));
    defparam i1_2_lut_4_lut_adj_985.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_986 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [22]), .O(n25508));
    defparam i1_2_lut_4_lut_adj_986.LUT_INIT = 16'hea00;
    SB_LUT4 i11428_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n15259));
    defparam i11428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_987 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [21]), .O(n25384));
    defparam i1_2_lut_4_lut_adj_987.LUT_INIT = 16'hea00;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n53), .I2(n62), 
            .I3(GND_net), .O(n52));
    defparam i1_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i3731_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n7480));   // verilog/coms.v(157[6] 159[9])
    defparam i3731_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14627_2_lut (.I0(\FRAME_MATCHER.state_31__N_2380[2] ), .I1(n4452), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2540[2] ));   // verilog/coms.v(259[6] 261[9])
    defparam i14627_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_988 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [15]), .O(n25490));
    defparam i1_2_lut_4_lut_adj_988.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_989 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [14]), .O(n25492));
    defparam i1_2_lut_4_lut_adj_989.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_990 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [13]), .O(n25494));
    defparam i1_2_lut_4_lut_adj_990.LUT_INIT = 16'hea00;
    SB_LUT4 i11429_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n15260));
    defparam i11429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_991 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [12]), .O(n25496));
    defparam i1_2_lut_4_lut_adj_991.LUT_INIT = 16'hea00;
    SB_LUT4 i11430_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n15261));
    defparam i11430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_992 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [11]), .O(n25498));
    defparam i1_2_lut_4_lut_adj_992.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_993 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [10]), .O(n25500));
    defparam i1_2_lut_4_lut_adj_993.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_994 (.I0(n8_adj_3676), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n10_adj_3684), .I3(\FRAME_MATCHER.state [9]), .O(n25502));
    defparam i1_2_lut_4_lut_adj_994.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_995 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [1]), .I3(n26605), .O(n6_adj_3661));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_996 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3685));
    defparam i6_4_lut_adj_996.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\data_in[3] [3]), .I1(\data_in[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_998 (.I0(n9), .I1(n14_adj_3685), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [1]), .O(n13606));
    defparam i7_4_lut_adj_998.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut_adj_999 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3686));
    defparam i4_4_lut_adj_999.LUT_INIT = 16'hfdff;
    SB_LUT4 i11431_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n15262));
    defparam i11431_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1000 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[6] [3]), .O(n26587));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1001 (.I0(n13892), .I1(n13867), .I2(\data_in_frame[10] [5]), 
            .I3(\data_in_frame[12] [7]), .O(n26620));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1001.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1002 (.I0(\data_in[2] [7]), .I1(n10_adj_3686), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n13641));
    defparam i5_3_lut_adj_1002.LUT_INIT = 16'hdfdf;
    SB_LUT4 i7_4_lut_adj_1003 (.I0(\data_in[1] [3]), .I1(n13641), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n18_adj_3687));
    defparam i7_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut_adj_1004 (.I0(\data_in[3] [7]), .I1(\data_in[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3688));
    defparam i5_2_lut_adj_1004.LUT_INIT = 16'hdddd;
    SB_LUT4 i9_4_lut_adj_1005 (.I0(\data_in[0] [5]), .I1(n18_adj_3687), 
            .I2(\data_in[2] [5]), .I3(\data_in[2] [6]), .O(n20_adj_3689));
    defparam i9_4_lut_adj_1005.LUT_INIT = 16'hfeff;
    SB_LUT4 i10_4_lut_adj_1006 (.I0(\data_in[1] [6]), .I1(n20_adj_3689), 
            .I2(n16_adj_3688), .I3(\data_in[2] [0]), .O(n13496));
    defparam i10_4_lut_adj_1006.LUT_INIT = 16'hfffd;
    SB_LUT4 i23287_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [2]), .I2(\data_in[0] [3]), 
            .I3(\data_in[1] [0]), .O(n28377));
    defparam i23287_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3690));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1008 (.I0(n9_adj_3690), .I1(n28377), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n13628));
    defparam i7_4_lut_adj_1008.LUT_INIT = 16'hffbf;
    SB_LUT4 i6_4_lut_adj_1009 (.I0(n13628), .I1(\data_in[3] [6]), .I2(\data_in[0] [7]), 
            .I3(n13496), .O(n16_adj_3691));
    defparam i6_4_lut_adj_1009.LUT_INIT = 16'hfffe;
    SB_LUT4 i23293_4_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n28383));
    defparam i23293_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i9_4_lut_adj_1010 (.I0(n28383), .I1(\data_in[3] [1]), .I2(n16_adj_3691), 
            .I3(\data_in[3] [5]), .O(n62));
    defparam i9_4_lut_adj_1010.LUT_INIT = 16'hf7ff;
    SB_LUT4 i6_4_lut_adj_1011 (.I0(\data_in[3] [0]), .I1(n13606), .I2(n13496), 
            .I3(\data_in[2] [2]), .O(n16_adj_3692));
    defparam i6_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1012 (.I0(\data_out_frame[5] [2]), .I1(n26096), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[5] [1]), .O(n13756));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1013 (.I0(\data_in[2] [4]), .I1(\data_in[1] [0]), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n17_adj_3693));
    defparam i7_4_lut_adj_1013.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1014 (.I0(n17_adj_3693), .I1(\data_in[0] [6]), 
            .I2(n16_adj_3692), .I3(\data_in[1] [4]), .O(n53));
    defparam i9_4_lut_adj_1014.LUT_INIT = 16'hfbff;
    SB_LUT4 i23277_2_lut (.I0(\data_in[3] [2]), .I1(\data_in[1] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n28365));
    defparam i23277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25070_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4040));
    defparam i25070_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i8_4_lut_adj_1015 (.I0(\data_in[3] [7]), .I1(n13628), .I2(n13606), 
            .I3(n13641), .O(n21));
    defparam i8_4_lut_adj_1015.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1016 (.I0(\data_in[1] [3]), .I1(\data_in[2] [5]), 
            .I2(\data_in[1] [6]), .I3(GND_net), .O(n20_adj_3694));
    defparam i7_3_lut_adj_1016.LUT_INIT = 16'hf7f7;
    SB_LUT4 i11_4_lut_adj_1017 (.I0(n21), .I1(\data_in[2] [6]), .I2(n28365), 
            .I3(\data_in[0] [5]), .O(n24_adj_3695));
    defparam i11_4_lut_adj_1017.LUT_INIT = 16'hefff;
    SB_LUT4 i12_4_lut_adj_1018 (.I0(\data_in[0] [1]), .I1(n24_adj_3695), 
            .I2(n20_adj_3694), .I3(\data_in[2] [0]), .O(n63));
    defparam i12_4_lut_adj_1018.LUT_INIT = 16'hfdff;
    SB_LUT4 i4_4_lut_adj_1019 (.I0(n5_adj_3696), .I1(n8_adj_3652), .I2(n14328), 
            .I3(n13972), .O(n17_adj_3697));
    defparam i4_4_lut_adj_1019.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1020 (.I0(n13919), .I1(n13892), .I2(n13867), 
            .I3(n14082), .O(n21_adj_3698));
    defparam i8_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1021 (.I0(n26498), .I1(n13852), .I2(n26034), 
            .I3(\data_in_frame[8] [1]), .O(n14_adj_3699));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1022 (.I0(n8_adj_3700), .I1(n28118), .I2(n14420), 
            .I3(\data_in_frame[8] [0]), .O(n20_adj_3701));
    defparam i7_4_lut_adj_1022.LUT_INIT = 16'hfbfe;
    SB_LUT4 i11_4_lut_adj_1023 (.I0(n21_adj_3698), .I1(n17_adj_3697), .I2(n23686), 
            .I3(n3_adj_3601), .O(n24_adj_3702));
    defparam i11_4_lut_adj_1023.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1024 (.I0(n23717), .I1(n14_adj_3699), .I2(n10_adj_3703), 
            .I3(Kp_23__N_698), .O(n27195));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1025 (.I0(\data_out_frame[5] [2]), .I1(n26096), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[9] [4]), .O(n13906));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1026 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n26370));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1027 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(Kp_23__N_708), .I3(\data_in_frame[3] [0]), .O(n26167));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1028 (.I0(\FRAME_MATCHER.state [3]), .I1(n21466), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n4040), .O(n63_adj_3));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1028.LUT_INIT = 16'hfdff;
    SB_CARRY add_43_23 (.CI(n21956), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n21957));
    SB_LUT4 i4_4_lut_adj_1029 (.I0(n63_adj_3), .I1(n13621), .I2(n13610), 
            .I3(n13611), .O(n10_adj_3705));
    defparam i4_4_lut_adj_1029.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut_adj_1030 (.I0(n13651), .I1(n10_adj_3705), .I2(n18939), 
            .I3(GND_net), .O(n2254));
    defparam i5_3_lut_adj_1030.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut_adj_1031 (.I0(n63), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n53), .I3(n62), .O(\FRAME_MATCHER.state_31__N_2380 [0]));
    defparam i3_4_lut_adj_1031.LUT_INIT = 16'hdfff;
    SB_LUT4 i12_4_lut_adj_1032 (.I0(n27195), .I1(n24_adj_3702), .I2(n20_adj_3701), 
            .I3(n14297), .O(n1));
    defparam i12_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1033 (.I0(\data_in_frame[7] [6]), .I1(n14017), 
            .I2(n13808), .I3(GND_net), .O(n13988));
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n13937));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1035 (.I0(\data_in_frame[6] [7]), .I1(n26629), 
            .I2(\data_in_frame[6] [4]), .I3(GND_net), .O(n26034));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1035.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3706));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1037 (.I0(n26333), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(n6_adj_3706), .O(n26028));
    defparam i4_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_0__2__I_0_2_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_698));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_0__2__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1038 (.I0(\data_in_frame[9] [3]), .I1(Kp_23__N_1053), 
            .I2(n26059), .I3(\data_in_frame[11] [5]), .O(n23761));
    defparam i2_3_lut_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1039 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n26113));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1039.LUT_INIT = 16'h9696;
    SB_LUT4 i14691_4_lut (.I0(n8_adj_3707), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n13625), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i14691_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_3708));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1040 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1041 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(n13508), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n13651));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1041.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_3_lut_adj_1042 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n26155));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1042.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_22_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n21955), .O(n2_adj_3709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44_adj_3708), 
            .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_22 (.CI(n21955), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n21956));
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n13625));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\FRAME_MATCHER.i [4]), .I1(n13625), .I2(GND_net), 
            .I3(GND_net), .O(n13505));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1044 (.I0(\data_in_frame[5] [4]), .I1(n26370), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n13808));
    defparam i2_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1045 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[4] [3]), .O(n26040));   // verilog/coms.v(166[9:87])
    defparam i3_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26134));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(n14396), .I1(\data_in_frame[3] [5]), 
            .I2(n8_adj_3710), .I3(\data_in_frame[5] [3]), .O(n10_adj_3711));
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut (.I0(n13794), .I1(n26028), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_3712));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14563_4_lut (.I0(n8_adj_3713), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n13505), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i14563_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i7_4_lut_adj_1048 (.I0(n26134), .I1(n26297), .I2(n26120), 
            .I3(n10_adj_3711), .O(n16_adj_3714));
    defparam i7_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1049 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(n13508), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n13611));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1049.LUT_INIT = 16'hfffd;
    SB_LUT4 i2_2_lut_adj_1050 (.I0(\FRAME_MATCHER.state [0]), .I1(n28307), 
            .I2(GND_net), .I3(GND_net), .O(n13615));   // verilog/coms.v(222[5:21])
    defparam i2_2_lut_adj_1050.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1051 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(n13508), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n13610));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1051.LUT_INIT = 16'hffdf;
    SB_LUT4 i14632_4_lut (.I0(n5_adj_3715), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i14632_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i21601_2_lut (.I0(n13620), .I1(n4452), .I2(GND_net), .I3(GND_net), 
            .O(n26676));
    defparam i21601_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_in_frame[6] [0]), .I1(n26498), .I2(n26370), 
            .I3(GND_net), .O(n11));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\FRAME_MATCHER.state [0]), .I1(n13616), 
            .I2(GND_net), .I3(GND_net), .O(n13618));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'hdddd;
    SB_LUT4 i11416_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n15247));
    defparam i11416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1053 (.I0(n13618), .I1(n26676), .I2(n771), .I3(n26678), 
            .O(n27507));
    defparam i2_4_lut_adj_1053.LUT_INIT = 16'hc800;
    SB_LUT4 i3_4_lut_adj_1054 (.I0(\FRAME_MATCHER.state [3]), .I1(n21466), 
            .I2(n4040), .I3(\FRAME_MATCHER.state [0]), .O(n28267));
    defparam i3_4_lut_adj_1054.LUT_INIT = 16'h0020;
    SB_LUT4 i11417_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n15248));
    defparam i11417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1055 (.I0(n26040), .I1(n16_adj_3714), .I2(n12_adj_3712), 
            .I3(n13808), .O(n23717));
    defparam i8_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1056 (.I0(n14017), .I1(Kp_23__N_888), .I2(n14153), 
            .I3(n26387), .O(n10_adj_3717));
    defparam i4_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n13950));
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(n14396), .I1(\data_in_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26223));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1059 (.I0(n26505), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[10] [0]), .I3(GND_net), .O(n23702));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1059.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1060 (.I0(\data_in_frame[10] [2]), .I1(n26402), 
            .I2(n26223), .I3(n13950), .O(n13_adj_3718));
    defparam i5_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1061 (.I0(n13_adj_3718), .I1(n11), .I2(n28118), 
            .I3(\data_in_frame[7] [6]), .O(n14380));
    defparam i7_4_lut_adj_1061.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1062 (.I0(\data_in_frame[6] [0]), .I1(n26498), 
            .I2(n26205), .I3(GND_net), .O(n12033));
    defparam i1_2_lut_3_lut_adj_1062.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1063 (.I0(n28267), .I1(\FRAME_MATCHER.state_31__N_2380 [0]), 
            .I2(n27507), .I3(GND_net), .O(n25624));
    defparam i1_3_lut_adj_1063.LUT_INIT = 16'haeae;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\FRAME_MATCHER.state_31__N_2380 [0]), .I1(n6), 
            .I2(GND_net), .I3(GND_net), .O(n25396));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_21_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n21954), .O(n2_adj_3720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1065 (.I0(n14017), .I1(n14396), .I2(\data_in_frame[5] [5]), 
            .I3(n23717), .O(n26283));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1066 (.I0(n14017), .I1(n14396), .I2(\data_in_frame[5] [5]), 
            .I3(\data_in_frame[7] [7]), .O(n26205));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_CARRY add_43_21 (.CI(n21954), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n21955));
    SB_LUT4 i11418_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n15249));
    defparam i11418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[6] [2]), .I1(Kp_23__N_656), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3721));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [3]), 
            .I2(Kp_23__N_810), .I3(n6_adj_3721), .O(n13867));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1069 (.I0(n13867), .I1(n26087), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n12058));
    defparam i2_3_lut_adj_1069.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26457));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26361));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1072 (.I0(\data_in_frame[18] [6]), .I1(n26554), 
            .I2(n26584), .I3(n26361), .O(n26323));
    defparam i1_4_lut_adj_1072.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1073 (.I0(n26031), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[6] [5]), .I3(n26432), .O(n10_adj_3722));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1074 (.I0(\data_in_frame[2] [3]), .I1(n10_adj_3722), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n8_adj_3700));   // verilog/coms.v(73[16:42])
    defparam i5_3_lut_adj_1074.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26656));
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1076 (.I0(\data_in_frame[13] [1]), .I1(n26656), 
            .I2(\data_in_frame[11] [0]), .I3(n8_adj_3700), .O(n26208));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1077 (.I0(\data_in_frame[10] [5]), .I1(n26581), 
            .I2(n26208), .I3(\data_in_frame[12] [6]), .O(n14308));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1078 (.I0(n23700), .I1(\data_in_frame[17] [5]), 
            .I2(n14308), .I3(\data_in_frame[17] [4]), .O(n26274));
    defparam i1_4_lut_adj_1078.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26653));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1080 (.I0(\data_in_frame[4] [4]), .I1(n26653), 
            .I2(\data_in_frame[4] [2]), .I3(\data_in_frame[2] [0]), .O(n26031));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1081 (.I0(\data_in_frame[4] [3]), .I1(Kp_23__N_713), 
            .I2(\data_in_frame[8] [7]), .I3(n13852), .O(n12_adj_3723));   // verilog/coms.v(73[16:42])
    defparam i5_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1082 (.I0(\data_in_frame[6] [6]), .I1(n12_adj_3723), 
            .I2(n26031), .I3(\data_in_frame[4] [5]), .O(Kp_23__N_1030));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1083 (.I0(n13919), .I1(n8_adj_3652), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1041));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1084 (.I0(Kp_23__N_1041), .I1(Kp_23__N_1030), .I2(\data_in_frame[13] [5]), 
            .I3(Kp_23__N_1256), .O(n12_adj_3724));
    defparam i5_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1085 (.I0(\data_in_frame[16] [0]), .I1(n12_adj_3724), 
            .I2(\data_in_frame[16] [1]), .I3(\data_in_frame[14] [0]), .O(n26117));
    defparam i6_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26183));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(\data_in_frame[18] [2]), .I1(n26183), 
            .I2(n24689), .I3(\data_in_frame[15] [6]), .O(n10_adj_3725));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1088 (.I0(n26117), .I1(n10_adj_3725), .I2(n13877), 
            .I3(GND_net), .O(n23768));
    defparam i5_3_lut_adj_1088.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1256));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1089 (.I0(\data_in_frame[16] [2]), .I1(n26056), 
            .I2(n24652), .I3(Kp_23__N_1256), .O(n10_adj_3726));
    defparam i4_4_lut_adj_1089.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26220));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1091 (.I0(n14017), .I1(n26420), .I2(n26220), 
            .I3(\data_in_frame[5] [6]), .O(n13794));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n14994));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26016));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i25140_2_lut (.I0(n19121), .I1(n6_adj_3727), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3233));
    defparam i25140_2_lut.LUT_INIT = 16'h1111;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n14993));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1093 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n14017));
    defparam i1_2_lut_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i14594_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3336[0]), .I2(GND_net), 
            .I3(GND_net), .O(n806));
    defparam i14594_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n14715), .D(n3965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1094 (.I0(n23741), .I1(\data_out_frame[14] [5]), 
            .I2(n26300), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i11419_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n15250));
    defparam i11419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15138_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n18966));
    defparam i15138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1095 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n18966), .I3(byte_transmit_counter[2]), .O(n19121));
    defparam i2_4_lut_adj_1095.LUT_INIT = 16'h8880;
    SB_LUT4 i2_3_lut_adj_1096 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n6_adj_3727));
    defparam i2_3_lut_adj_1096.LUT_INIT = 16'hfefe;
    SB_LUT4 add_43_20_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n21953), .O(n2_adj_3728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i21707_3_lut (.I0(n21466), .I1(n26688), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n26785));
    defparam i21707_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26420));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26217));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1099 (.I0(n19121), .I1(n806), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_3729));
    defparam i2_2_lut_adj_1099.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1100 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(n26205), .I3(GND_net), .O(n6_adj_3730));
    defparam i1_2_lut_3_lut_adj_1100.LUT_INIT = 16'h9696;
    SB_LUT4 mux_712_i1_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n7_adj_3729), 
            .I2(n18983), .I3(n8_adj_3731), .O(n2813[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_712_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i2_3_lut_4_lut_adj_1101 (.I0(\data_in_frame[3] [5]), .I1(n26420), 
            .I2(n26297), .I3(\data_in_frame[1] [6]), .O(Kp_23__N_656));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1102 (.I0(\data_in_frame[3] [5]), .I1(n26420), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[3] [6]), .O(n26498));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1103 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n6_adj_3727), .I3(\FRAME_MATCHER.state [2]), .O(n8_adj_3731));
    defparam i3_3_lut_4_lut_adj_1103.LUT_INIT = 16'hf7ff;
    SB_LUT4 i11420_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n15251));
    defparam i11420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11421_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n15252));
    defparam i11421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1104 (.I0(n12033), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[8] [1]), .I3(GND_net), .O(n26087));
    defparam i2_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1105 (.I0(\data_in_frame[8] [2]), .I1(n26016), 
            .I2(n13794), .I3(Kp_23__N_656), .O(n3_adj_3601));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n13877));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i11422_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n15253));
    defparam i11422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11423_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n15254));
    defparam i11423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14740_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n21466), .I3(GND_net), .O(n18565));
    defparam i14740_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n6_adj_3583));
    defparam i1_4_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i21611_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n26688));
    defparam i21611_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1107 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(n26490), .I3(GND_net), .O(n26611));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1108 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [7]), .O(n26297));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(n10_adj_3717), .I3(n23717), .O(n28118));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1109 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[9] [0]), .I3(n13347), .O(n26608));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 mux_985_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n3963), .I3(GND_net), .O(n3964));
    defparam mux_985_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1110 (.I0(\data_out_frame[12] [4]), .I1(n26093), 
            .I2(n14219), .I3(GND_net), .O(n26300));
    defparam i1_2_lut_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_CARRY add_43_20 (.CI(n21953), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n21954));
    SB_LUT4 add_43_19_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n21952), .O(n2_adj_3732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1111 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n6_adj_3733));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3734));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3735));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1112 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(n3_adj_3601), .I3(\data_in_frame[10] [4]), .O(n26581));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i24457_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29242));
    defparam i24457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24459_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29241));
    defparam i24459_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3736));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3737));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24471_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29239));
    defparam i24471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24473_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29238));
    defparam i24473_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3738));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3739));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24476_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29236));
    defparam i24476_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1113 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3740));
    defparam i2_2_lut_adj_1113.LUT_INIT = 16'heeee;
    SB_LUT4 i24465_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29235));
    defparam i24465_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[11] [1]), .I1(n27074), 
            .I2(GND_net), .I3(GND_net), .O(n24696));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1115 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(\FRAME_MATCHER.state [8]), 
            .O(n14_adj_3741));
    defparam i6_4_lut_adj_1115.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1116 (.I0(\FRAME_MATCHER.state [10]), .I1(n14_adj_3741), 
            .I2(n10_adj_3740), .I3(\FRAME_MATCHER.state [15]), .O(n25892));
    defparam i7_4_lut_adj_1116.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3742));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1117 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[10] [6]), .I3(n26043), .O(n14_adj_3743));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3744));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3745));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1118 (.I0(\data_in_frame[10] [7]), .I1(n14_adj_3743), 
            .I2(n10_adj_3746), .I3(n26623), .O(n26110));   // verilog/coms.v(85[17:70])
    defparam i7_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i24482_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29232));
    defparam i24482_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10_4_lut_adj_1119 (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [22]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n24_adj_3747));
    defparam i10_4_lut_adj_1119.LUT_INIT = 16'hfffe;
    SB_LUT4 i24485_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29231));
    defparam i24485_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(n24696), .I1(n26620), .I2(n26211), 
            .I3(\data_in_frame[10] [6]), .O(n23692));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1121 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [16]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n22_adj_3748));
    defparam i8_4_lut_adj_1121.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3749));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3750));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24486_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29229));
    defparam i24486_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1122 (.I0(\FRAME_MATCHER.state [17]), .I1(n24_adj_3747), 
            .I2(n18_adj_3745), .I3(\FRAME_MATCHER.state [28]), .O(n26));
    defparam i12_4_lut_adj_1122.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26239));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i24488_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29228));
    defparam i24488_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11_3_lut (.I0(\FRAME_MATCHER.state [23]), .I1(n22_adj_3748), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n25));
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut_4_lut_adj_1124 (.I0(\data_in_frame[4] [1]), .I1(n13675), 
            .I2(n26494), .I3(n26502), .O(n8_adj_3710));   // verilog/coms.v(78[16:27])
    defparam i3_3_lut_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1125 (.I0(n26494), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[7] [2]), .I3(n26527), .O(n10_adj_3751));
    defparam i4_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1126 (.I0(n25), .I1(\FRAME_MATCHER.state [18]), 
            .I2(n26), .I3(\FRAME_MATCHER.state [20]), .O(n19125));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1127 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [7]), .I3(\data_in_frame[9] [4]), .O(n26202));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_in_frame[11] [7]), .I1(n26202), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3752));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1129 (.I0(n23686), .I1(n13892), .I2(n13877), 
            .I3(n6_adj_3752), .O(n24523));
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1130 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3753));
    defparam i2_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(n7_adj_3753), .I1(\data_in_frame[14] [3]), 
            .I2(n24523), .I3(n27069), .O(n26286));
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1132 (.I0(n24618), .I1(n24578), .I2(\data_in_frame[16] [4]), 
            .I3(n26286), .O(n10_adj_3754));
    defparam i4_4_lut_adj_1132.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1133 (.I0(n14383), .I1(n10_adj_3754), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n13377));
    defparam i5_3_lut_adj_1133.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1134 (.I0(n13377), .I1(n26330), .I2(n24533), 
            .I3(GND_net), .O(n12137));
    defparam i2_3_lut_adj_1134.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1135 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [5]), 
            .I2(n26336), .I3(\data_in_frame[19] [4]), .O(n6_adj_3755));
    defparam i2_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1136 (.I0(\data_in_frame[19] [1]), .I1(n6_adj_3755), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [3]), .O(n24249));
    defparam i3_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1137 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [6]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n25894));
    defparam i3_4_lut_adj_1137.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1138 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[7] [1]), .I3(n14677), .O(n12_adj_3756));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1139 (.I0(n25894), .I1(n19125), .I2(n25892), 
            .I3(GND_net), .O(n21466));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_1139.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1140 (.I0(\data_in_frame[2] [6]), .I1(n12_adj_3756), 
            .I2(n26239), .I3(n14153), .O(n14328));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n14328), .I1(n14420), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1053));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\FRAME_MATCHER.state [3]), .I1(n21466), 
            .I2(GND_net), .I3(GND_net), .O(n13508));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1143 (.I0(n26056), .I1(n26289), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n13964));
    defparam i2_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_LUT4 i23248_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n28307), .I2(n13508), 
            .I3(\FRAME_MATCHER.state [2]), .O(n18939));
    defparam i23248_4_lut.LUT_INIT = 16'hddd5;
    SB_LUT4 i4_4_lut_adj_1144 (.I0(n24696), .I1(n26289), .I2(\data_in_frame[15] [5]), 
            .I3(\data_in_frame[13] [4]), .O(n10_adj_3757));
    defparam i4_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i15112_1_lut (.I0(n18939), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1656));
    defparam i15112_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(n26286), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3758));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1146 (.I0(n24618), .I1(n14005), .I2(\data_in_frame[16] [5]), 
            .I3(\data_in_frame[14] [5]), .O(n12_adj_3759));
    defparam i5_4_lut_adj_1146.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1147 (.I0(\data_in_frame[18] [7]), .I1(n13788), 
            .I2(n12_adj_3759), .I3(n8_adj_3758), .O(n26172));
    defparam i1_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_in_frame[16] [5]), .I1(n24560), 
            .I2(GND_net), .I3(GND_net), .O(n26584));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26333));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n13675));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1151 (.I0(\data_in_frame[5] [0]), .I1(n26167), 
            .I2(\data_in_frame[4] [6]), .I3(GND_net), .O(n26494));
    defparam i2_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26175));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26432));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(Kp_23__N_888), .I1(n26283), .I2(GND_net), 
            .I3(GND_net), .O(n26284));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1155 (.I0(\data_in_frame[7] [7]), .I1(n13950), 
            .I2(n26653), .I3(\data_in_frame[9] [2]), .O(n21_adj_3760));
    defparam i8_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_adj_1156 (.I0(\data_in_frame[7] [0]), .I1(n26587), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n20_adj_3761));
    defparam i7_3_lut_adj_1156.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1157 (.I0(n21_adj_3760), .I1(n27069), .I2(n18_adj_3762), 
            .I3(n26641), .O(n24_adj_3763));
    defparam i11_4_lut_adj_1157.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1158 (.I0(\data_in_frame[8] [7]), .I1(n24_adj_3763), 
            .I2(n20_adj_3761), .I3(n13675), .O(n24566));
    defparam i12_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1159 (.I0(n26151), .I1(n26155), .I2(n14237), 
            .I3(n1427), .O(n26647));
    defparam i2_3_lut_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n24523), .I1(n23743), .I2(n23702), .I3(n18_adj_3764), 
            .O(n30_adj_3765));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1160 (.I0(n24566), .I1(n26557), .I2(n26284), 
            .I3(n26432), .O(n28));
    defparam i11_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_15__7__I_0_3897_2_lut (.I0(\data_in_frame[15] [7]), 
            .I1(\data_in_frame[15] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1237));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_15__7__I_0_3897_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_63_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3766));
    defparam equal_63_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[14] [2]), .I3(GND_net), .O(n26596));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1162 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[14] [7]), 
            .I2(n26180), .I3(n14216), .O(n8));   // verilog/coms.v(85[17:28])
    defparam i3_3_lut_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i11408_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n15239));
    defparam i11408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1163 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[4] [3]), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[11] [7]), .O(n29_adj_3767));
    defparam i12_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1164 (.I0(n26175), .I1(n26494), .I2(\data_in_frame[12] [0]), 
            .I3(\data_in_frame[4] [7]), .O(n27_adj_3768));
    defparam i10_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1165 (.I0(n27_adj_3768), .I1(n29_adj_3767), .I2(n28), 
            .I3(n30_adj_3765), .O(n24560));
    defparam i16_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 equal_64_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3713));
    defparam equal_64_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1166 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[4] [6]), .I3(\data_in_frame[0] [3]), .O(n26189));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_in_frame[11] [6]), .I1(n24652), 
            .I2(GND_net), .I3(GND_net), .O(n24689));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1168 (.I0(n26016), .I1(n26629), .I2(\data_in_frame[11] [5]), 
            .I3(n26283), .O(n20_adj_3769));
    defparam i8_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1169 (.I0(n26189), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[13] [7]), .I3(n26533), .O(n19));
    defparam i7_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1170 (.I0(n26077), .I1(n13391), .I2(n13852), 
            .I3(n24566), .O(n21_adj_3770));
    defparam i9_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1171 (.I0(n21_adj_3770), .I1(n19), .I2(n20_adj_3769), 
            .I3(GND_net), .O(n24578));
    defparam i11_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1172 (.I0(n24578), .I1(\data_in_frame[16] [1]), 
            .I2(n23761), .I3(n14665), .O(n10_adj_3771));
    defparam i4_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3622));
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2_3_lut_adj_1173 (.I0(n24560), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[16] [3]), .I3(GND_net), .O(n26426));
    defparam i2_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1174 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[6] [4]), .I3(\data_in_frame[4] [3]), .O(n26077));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(\data_in_frame[8] [5]), .I1(n26077), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n26460));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26533));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26641));
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_713));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1178 (.I0(n23686), .I1(\data_in_frame[9] [5]), 
            .I2(n13972), .I3(GND_net), .O(n23747));
    defparam i2_3_lut_adj_1178.LUT_INIT = 16'h9696;
    SB_LUT4 i11409_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n15240));
    defparam i11409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15150_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n18978));
    defparam i15150_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1363_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_3707));
    defparam i1363_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_4_lut_adj_1179 (.I0(n13508), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n13621));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1179.LUT_INIT = 16'hffef;
    SB_LUT4 i22_4_lut (.I0(n26361), .I1(n27074), .I2(n26043), .I3(\data_in_frame[18] [7]), 
            .O(n61));
    defparam i22_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut (.I0(n26659), .I1(Kp_23__N_1237), .I2(n26211), .I3(n26626), 
            .O(n60));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[15] [4]), .I3(\data_in_frame[18] [5]), .O(n68));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n55));
    defparam i16_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i27_4_lut (.I0(n23768), .I1(n26117), .I2(n26274), .I3(n26081), 
            .O(n66));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1180 (.I0(\data_in_frame[18] [1]), .I1(n26656), 
            .I2(n13723), .I3(n26635), .O(n64));
    defparam i25_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n26605), .I1(n26447), .I2(n26508), .I3(n26441), 
            .O(n65));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1181 (.I0(n26090), .I1(n23747), .I2(Kp_23__N_713), 
            .I3(n23761), .O(n63_adj_3772));
    defparam i24_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n61), .I1(n26641), .I2(n46), .I3(n26533), 
            .O(n70));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(Kp_23__N_1218), .I1(n60), .I2(\data_in_frame[8] [1]), 
            .I3(n26460), .O(n69));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34_4_lut (.I0(n55), .I1(n68), .I2(\data_in_frame[9] [1]), 
            .I3(n23743), .O(n73));
    defparam i34_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i36_4_lut (.I0(n63_adj_3772), .I1(n65), .I2(n64), .I3(n66), 
            .O(n75));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i38_4_lut (.I0(n75), .I1(n73), .I2(n69), .I3(n70), .O(n24533));
    defparam i38_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1182 (.I0(n26426), .I1(n26399), .I2(n26539), 
            .I3(n23770), .O(n26330));
    defparam i2_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1183 (.I0(\data_in_frame[2] [7]), .I1(Kp_23__N_708), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n26252));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1184 (.I0(n26252), .I1(\data_in_frame[5] [1]), 
            .I2(n26131), .I3(GND_net), .O(n26527));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1185 (.I0(Kp_23__N_708), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[3] [1]), .I3(GND_net), .O(n14599));
    defparam i2_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1186 (.I0(n14599), .I1(n26527), .I2(n26239), 
            .I3(\data_in_frame[5] [2]), .O(n26120));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n14677));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(n23686), .I1(n14420), .I2(GND_net), 
            .I3(GND_net), .O(n13391));
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[11] [4]), .I1(n26059), 
            .I2(GND_net), .I3(GND_net), .O(n26447));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_in_frame[9] [2]), .I1(n14328), 
            .I2(GND_net), .I3(GND_net), .O(n26090));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1191 (.I0(\data_in_frame[11] [5]), .I1(n13873), 
            .I2(\data_in_frame[16] [0]), .I3(n6_adj_3773), .O(n23770));
    defparam i4_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1218));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1192 (.I0(n26423), .I1(\data_in_frame[18] [1]), 
            .I2(n23770), .I3(GND_net), .O(n26381));
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1193 (.I0(\data_in_frame[0] [5]), .I1(n26252), 
            .I2(\data_in_frame[5] [3]), .I3(GND_net), .O(n14130));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1193.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1194 (.I0(\data_in_frame[1] [4]), .I1(n26484), 
            .I2(n26217), .I3(\data_in_frame[1] [3]), .O(Kp_23__N_708));   // verilog/coms.v(73[16:34])
    defparam i3_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26131));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1196 (.I0(\data_in_frame[5] [2]), .I1(n26370), 
            .I2(n14130), .I3(\data_in_frame[7] [4]), .O(n26557));
    defparam i3_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30562));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30562_bdd_4_lut (.I0(n30562), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30565));
    defparam n30562_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1197 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[11] [3]), 
            .I2(n8_adj_3774), .I3(n13873), .O(n26560));
    defparam i1_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(n23692), .I1(n26110), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n23706));
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n30295), .I2(n29240), .I3(byte_transmit_counter[4]), .O(n30550));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1199 (.I0(n13508), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n4_adj_3775));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1199.LUT_INIT = 16'h1000;
    SB_LUT4 n30550_bdd_4_lut (.I0(n30550), .I1(n14_adj_3648), .I2(n7_adj_3647), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n30550_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(n23706), .I1(n26560), .I2(Kp_23__N_1237), 
            .I3(GND_net), .O(n26399));
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25420 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30544));
    defparam byte_transmit_counter_0__bdd_4_lut_25420.LUT_INIT = 16'he4aa;
    SB_LUT4 n30544_bdd_4_lut (.I0(n30544), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30547));
    defparam n30544_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1201 (.I0(\data_in_frame[17] [7]), .I1(n14665), 
            .I2(n23700), .I3(GND_net), .O(n26423));
    defparam i2_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25411 (.I0(byte_transmit_counter[3]), 
            .I1(n30301), .I2(n29237), .I3(byte_transmit_counter[4]), .O(n30538));
    defparam byte_transmit_counter_3__bdd_4_lut_25411.LUT_INIT = 16'he4aa;
    SB_LUT4 n30538_bdd_4_lut (.I0(n30538), .I1(n14_adj_3644), .I2(n7_adj_3643), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n30538_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26387));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25401 (.I0(byte_transmit_counter[3]), 
            .I1(n30307), .I2(n29233), .I3(byte_transmit_counter[4]), .O(n30532));
    defparam byte_transmit_counter_3__bdd_4_lut_25401.LUT_INIT = 16'he4aa;
    SB_LUT4 n30532_bdd_4_lut (.I0(n30532), .I1(n14_adj_3640), .I2(n7_adj_3639), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n30532_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1203 (.I0(\data_in_frame[7] [5]), .I1(n26223), 
            .I2(n14599), .I3(n14130), .O(n14082));
    defparam i3_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25396 (.I0(byte_transmit_counter[3]), 
            .I1(n30313), .I2(n29230), .I3(byte_transmit_counter[4]), .O(n30526));
    defparam byte_transmit_counter_3__bdd_4_lut_25396.LUT_INIT = 16'he4aa;
    SB_LUT4 n30526_bdd_4_lut (.I0(n30526), .I1(n14_adj_3636), .I2(n7_adj_3635), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n30526_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_4_lut_adj_1204 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [5]), .O(n8_adj_3776));   // verilog/coms.v(74[16:27])
    defparam i3_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25391 (.I0(byte_transmit_counter[3]), 
            .I1(n30319), .I2(n29227), .I3(byte_transmit_counter[4]), .O(n30520));
    defparam byte_transmit_counter_3__bdd_4_lut_25391.LUT_INIT = 16'he4aa;
    SB_LUT4 n30520_bdd_4_lut (.I0(n30520), .I1(n14_adj_3633), .I2(n7_adj_3632), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n30520_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1205 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[8] [0]), 
            .I2(n26387), .I3(n6_adj_3730), .O(n26081));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25406 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30514));
    defparam byte_transmit_counter_0__bdd_4_lut_25406.LUT_INIT = 16'he4aa;
    SB_LUT4 n30514_bdd_4_lut (.I0(n30514), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30517));
    defparam n30514_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n13788));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25381 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30508));
    defparam byte_transmit_counter_0__bdd_4_lut_25381.LUT_INIT = 16'he4aa;
    SB_LUT4 n30508_bdd_4_lut (.I0(n30508), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30511));
    defparam n30508_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26441));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1208 (.I0(n13508), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n13620));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1208.LUT_INIT = 16'hefff;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_in_frame[10] [1]), .I1(n26081), 
            .I2(\data_in_frame[9] [7]), .I3(n14082), .O(n14383));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25376 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30496));
    defparam byte_transmit_counter_0__bdd_4_lut_25376.LUT_INIT = 16'he4aa;
    SB_LUT4 n30496_bdd_4_lut (.I0(n30496), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30499));
    defparam n30496_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1210 (.I0(\data_out_frame[16] [3]), .I1(n26569), 
            .I2(n14116), .I3(n26429), .O(n13369));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25366 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30490));
    defparam byte_transmit_counter_0__bdd_4_lut_25366.LUT_INIT = 16'he4aa;
    SB_LUT4 n30490_bdd_4_lut (.I0(n30490), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30493));
    defparam n30490_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1211 (.I0(\data_in_frame[17] [3]), .I1(n14308), 
            .I2(n26064), .I3(n6_adj_3733), .O(n13723));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25361 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30484));
    defparam byte_transmit_counter_0__bdd_4_lut_25361.LUT_INIT = 16'he4aa;
    SB_LUT4 n30484_bdd_4_lut (.I0(n30484), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30487));
    defparam n30484_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1212 (.I0(\data_in_frame[10] [5]), .I1(n26053), 
            .I2(\data_in_frame[14] [7]), .I3(\data_in_frame[12] [5]), .O(n12_adj_3777));
    defparam i5_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1213 (.I0(n14383), .I1(n12_adj_3777), .I2(n26441), 
            .I3(n13788), .O(n14205));
    defparam i6_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25356 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n30472));
    defparam byte_transmit_counter_0__bdd_4_lut_25356.LUT_INIT = 16'he4aa;
    SB_LUT4 n30472_bdd_4_lut (.I0(n30472), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n30475));
    defparam n30472_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1214 (.I0(n26460), .I1(n26587), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n13892));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25346 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30466));
    defparam byte_transmit_counter_0__bdd_4_lut_25346.LUT_INIT = 16'he4aa;
    SB_LUT4 n30466_bdd_4_lut (.I0(n30466), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30469));
    defparam n30466_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1215 (.I0(n14380), .I1(n23702), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[12] [3]), .O(n26554));
    defparam i3_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25341 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30460));
    defparam byte_transmit_counter_0__bdd_4_lut_25341.LUT_INIT = 16'he4aa;
    SB_LUT4 n30460_bdd_4_lut (.I0(n30460), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30463));
    defparam n30460_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1216 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[12] [5]), 
            .I2(n26067), .I3(\data_in_frame[16] [7]), .O(n18_adj_3778));   // verilog/coms.v(76[16:43])
    defparam i7_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25336 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n30454));
    defparam byte_transmit_counter_0__bdd_4_lut_25336.LUT_INIT = 16'he4aa;
    SB_LUT4 n30454_bdd_4_lut (.I0(n30454), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n30457));
    defparam n30454_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[17] [2]), .I1(n26208), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3779));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25331 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30448));
    defparam byte_transmit_counter_0__bdd_4_lut_25331.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1218 (.I0(n13972), .I1(n13988), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n26505));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_CARRY add_43_19 (.CI(n21952), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n21953));
    SB_LUT4 i2_3_lut_4_lut_adj_1219 (.I0(n13972), .I1(n13988), .I2(n28118), 
            .I3(n23686), .O(n26508));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1219.LUT_INIT = 16'h9669;
    SB_LUT4 n30448_bdd_4_lut (.I0(n30448), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30451));
    defparam n30448_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_adj_1220 (.I0(\data_in_frame[21] [6]), .I1(\data_in_frame[19] [5]), 
            .I2(\data_in_frame[19] [4]), .I3(GND_net), .O(n12_adj_3780));
    defparam i3_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25326 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30442));
    defparam byte_transmit_counter_0__bdd_4_lut_25326.LUT_INIT = 16'he4aa;
    SB_LUT4 n30442_bdd_4_lut (.I0(n30442), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30445));
    defparam n30442_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1221 (.I0(n26067), .I1(\data_in_frame[17] [4]), 
            .I2(n23692), .I3(n10_adj_3779), .O(n16_adj_3781));
    defparam i7_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25321 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30436));
    defparam byte_transmit_counter_0__bdd_4_lut_25321.LUT_INIT = 16'he4aa;
    SB_LUT4 n30436_bdd_4_lut (.I0(n30436), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30439));
    defparam n30436_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1222 (.I0(n13377), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[18] [4]), .I3(\data_in_frame[18] [5]), .O(n10_adj_3782));
    defparam i4_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25316 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30430));
    defparam byte_transmit_counter_0__bdd_4_lut_25316.LUT_INIT = 16'he4aa;
    SB_LUT4 n30430_bdd_4_lut (.I0(n30430), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30433));
    defparam n30430_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1223 (.I0(n26524), .I1(n16_adj_3781), .I2(n12_adj_3780), 
            .I3(n26064), .O(n27617));
    defparam i8_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[21] [3]), .I1(n26172), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3783));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1225 (.I0(\data_in_frame[20] [4]), .I1(n23768), 
            .I2(n26539), .I3(GND_net), .O(n8_adj_3784));
    defparam i3_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25311 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30412));
    defparam byte_transmit_counter_0__bdd_4_lut_25311.LUT_INIT = 16'he4aa;
    SB_LUT4 n30412_bdd_4_lut (.I0(n30412), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30415));
    defparam n30412_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1226 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[19] [2]), 
            .I2(n14205), .I3(n6_adj_3783), .O(n27118));
    defparam i4_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(\data_in_frame[19] [5]), .I1(n26336), 
            .I2(\data_in_frame[21] [7]), .I3(n13723), .O(n28121));
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25296 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30400));
    defparam byte_transmit_counter_0__bdd_4_lut_25296.LUT_INIT = 16'he4aa;
    SB_LUT4 n30400_bdd_4_lut (.I0(n30400), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30403));
    defparam n30400_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_rep_15_2_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30955));
    defparam i1_rep_15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1228 (.I0(tx_transmit_N_3233), .I1(n806), 
            .I2(n13651), .I3(n2254), .O(n6));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut_adj_1228.LUT_INIT = 16'hff0e;
    SB_LUT4 i1_3_lut_4_lut_adj_1229 (.I0(tx_transmit_N_3233), .I1(n806), 
            .I2(n8634), .I3(n13651), .O(n3_adj_3658));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut_adj_1229.LUT_INIT = 16'h00e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1230 (.I0(n24654), .I1(n26319), .I2(\data_out_frame[16] [3]), 
            .I3(n26384), .O(n9_adj_3785));
    defparam i1_2_lut_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_out_frame[24] [1]), .I1(n26514), 
            .I2(n23733), .I3(\data_out_frame[19] [4]), .O(n38));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1231 (.I0(\data_in_frame[19] [0]), .I1(n12137), 
            .I2(n24249), .I3(GND_net), .O(n6_adj_3786));
    defparam i2_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1232 (.I0(n26426), .I1(n30955), .I2(n26539), 
            .I3(\data_in_frame[20] [5]), .O(n27002));
    defparam i2_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25386 (.I0(byte_transmit_counter[3]), 
            .I1(n30337), .I2(n29224), .I3(byte_transmit_counter[4]), .O(n30376));
    defparam byte_transmit_counter_3__bdd_4_lut_25386.LUT_INIT = 16'he4aa;
    SB_LUT4 n30376_bdd_4_lut (.I0(n30376), .I1(n14_adj_3628), .I2(n7_adj_3627), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n30376_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_adj_1233 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n11_adj_3787));
    defparam i1_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25269 (.I0(byte_transmit_counter[3]), 
            .I1(n30361), .I2(n29221), .I3(byte_transmit_counter[4]), .O(n30370));
    defparam byte_transmit_counter_3__bdd_4_lut_25269.LUT_INIT = 16'he4aa;
    SB_LUT4 n30370_bdd_4_lut (.I0(n30370), .I1(n14_adj_3624), .I2(n7_adj_3621), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n30370_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_3_lut (.I0(n26581), .I1(\data_in_frame[17] [2]), .I2(n26457), 
            .I3(GND_net), .O(n14_adj_3788));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n29219), .I2(n29220), .I3(byte_transmit_counter[2]), .O(n30364));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30364_bdd_4_lut (.I0(n30364), .I1(n17_adj_3618), .I2(n16_adj_3617), 
            .I3(byte_transmit_counter[2]), .O(n29670));
    defparam n30364_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1234 (.I0(\data_in_frame[12] [7]), .I1(n11_adj_3787), 
            .I2(\data_in_frame[12] [2]), .I3(n12_adj_3789), .O(n18_adj_3790));
    defparam i8_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25259 (.I0(byte_transmit_counter[1]), 
            .I1(n29222), .I2(n29223), .I3(byte_transmit_counter[2]), .O(n30358));
    defparam byte_transmit_counter_1__bdd_4_lut_25259.LUT_INIT = 16'he4aa;
    SB_LUT4 n30358_bdd_4_lut (.I0(n30358), .I1(n17_adj_3616), .I2(n16_adj_3615), 
            .I3(byte_transmit_counter[2]), .O(n30361));
    defparam n30358_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1235 (.I0(n26330), .I1(\data_in_frame[18] [5]), 
            .I2(n24533), .I3(\data_in_frame[20] [7]), .O(n4_adj_3791));
    defparam i1_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_25264 (.I0(byte_transmit_counter[3]), 
            .I1(n29670), .I2(n29218), .I3(byte_transmit_counter[4]), .O(n30352));
    defparam byte_transmit_counter_3__bdd_4_lut_25264.LUT_INIT = 16'he4aa;
    SB_LUT4 n30352_bdd_4_lut (.I0(n30352), .I1(n14_adj_3614), .I2(n7_adj_3613), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n30352_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1236 (.I0(n26554), .I1(n18_adj_3790), .I2(n14_adj_3788), 
            .I3(n13892), .O(n28125));
    defparam i9_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25286 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30346));
    defparam byte_transmit_counter_0__bdd_4_lut_25286.LUT_INIT = 16'he4aa;
    SB_LUT4 n30346_bdd_4_lut (.I0(n30346), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30349));
    defparam n30346_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_adj_1237 (.I0(n14205), .I1(n13723), .I2(\data_in_frame[21] [5]), 
            .I3(GND_net), .O(n8_adj_3792));
    defparam i3_3_lut_adj_1237.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25245 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n30340));
    defparam byte_transmit_counter_0__bdd_4_lut_25245.LUT_INIT = 16'he4aa;
    SB_LUT4 n30340_bdd_4_lut (.I0(n30340), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n30343));
    defparam n30340_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_292_Select_31_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_3793));
    defparam select_292_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_4_lut_adj_1238 (.I0(\data_out_frame[23] [2]), .I1(n13751), 
            .I2(n2122), .I3(\data_out_frame[23] [3]), .O(n2400));
    defparam i1_2_lut_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 select_292_Select_30_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_3794));
    defparam select_292_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_29_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_3795));
    defparam select_292_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i11410_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n15241));
    defparam i11410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1239 (.I0(n24544), .I1(n26070), .I2(n24554), 
            .I3(n24251), .O(n13751));
    defparam i1_2_lut_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 select_292_Select_28_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_3796));
    defparam select_292_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_27_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_3797));
    defparam select_292_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n14715), .D(n3966));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n14715), .D(n3967));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n14715), .D(n3968));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n14715), .D(n3969));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n14715), .D(n3970));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n14715), .D(n3971));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n14715), .D(n3972));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n14715), .D(n3973));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n14715), 
            .D(n3974));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n14715), 
            .D(n3975));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n14715), 
            .D(n3976));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n14715), 
            .D(n3977));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n14715), 
            .D(n3978));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n14715), 
            .D(n3979));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n14715), 
            .D(n3980));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n14715), 
            .D(n3981));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n14715), 
            .D(n3982));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n14715), 
            .D(n3983));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n14715), 
            .D(n3984));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n14715), 
            .D(n3985));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n14715), 
            .D(n3986));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n14715), 
            .D(n3987));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3637), .S(n3_adj_3798));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1240 (.I0(n24251), .I1(n26304), .I2(n24554), 
            .I3(n24544), .O(n23772));
    defparam i2_3_lut_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 select_292_Select_26_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_3799));
    defparam select_292_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i11411_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n15242));
    defparam i11411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11412_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n15243));
    defparam i11412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_292_Select_25_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_3800));
    defparam select_292_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_24_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_3801));
    defparam select_292_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_23_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_3802));
    defparam select_292_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_22_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_3803));
    defparam select_292_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i3_4_lut_adj_1241 (.I0(\data_in_frame[19] [7]), .I1(n26423), 
            .I2(n26399), .I3(\data_in_frame[20] [1]), .O(n27514));
    defparam i3_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 select_292_Select_21_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_3804));
    defparam select_292_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_20_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_3805));
    defparam select_292_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_19_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_3806));
    defparam select_292_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_18_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_3807));
    defparam select_292_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n14992));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[23] [0]), .I1(n23772), .I2(n24544), 
            .I3(GND_net), .O(n10_adj_3808));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_292_Select_17_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_3809));
    defparam select_292_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_4_lut_adj_1242 (.I0(\FRAME_MATCHER.state [0]), .I1(n13616), 
            .I2(n771), .I3(n8634), .O(n184));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_4_lut_adj_1242.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_4_lut_adj_1243 (.I0(\FRAME_MATCHER.state [0]), .I1(n28307), 
            .I2(n8634), .I3(n3303), .O(n44));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_1243.LUT_INIT = 16'h0020;
    SB_LUT4 select_292_Select_16_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_3810));
    defparam select_292_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_15_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_3811));
    defparam select_292_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_14_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_3812));
    defparam select_292_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3623), .S(n3_adj_3813));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3594), .S(n3_adj_3814));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3592), .S(n3_adj_3815));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3816));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3599), .S(n3_adj_3817));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3818), .S(n3_adj_3819));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3820), .S(n3_adj_3821));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3822), .S(n3_adj_3823));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3824), .S(n3_adj_3825));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3826), .S(n3_adj_3827));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3828), .S(n3_adj_3829));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3830), .S(n3_adj_3831));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3832), .S(n3_adj_3812));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3833), .S(n3_adj_3811));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3834), .S(n3_adj_3810));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3732), .S(n3_adj_3809));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3728), .S(n3_adj_3807));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3720), .S(n3_adj_3806));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3709), .S(n3_adj_3805));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3682), .S(n3_adj_3804));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3680), .S(n3_adj_3803));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3678), .S(n3_adj_3802));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3675), .S(n3_adj_3801));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3672), .S(n3_adj_3800));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3670), .S(n3_adj_3799));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3669), .S(n3_adj_3797));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3664), .S(n3_adj_3796));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3660), .S(n3_adj_3795));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3659), .S(n3_adj_3794));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3657), .S(n3_adj_3793));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_13_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_3831));
    defparam select_292_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_12_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_3829));
    defparam select_292_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_11_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_3827));
    defparam select_292_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n14763), .D(n26881));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_10_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_3825));
    defparam select_292_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_9_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_3823));
    defparam select_292_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n14763), .D(n28156));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n14763), .D(n26999));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n14763), .D(n27697));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n14763), .D(n26272));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n14763), .D(n27684));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n14763), .D(n26852));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n14763), .D(n27278));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n14763), .D(n26391));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n14763), .D(n26392));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n14763), .D(n11578));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n14763), .D(n26890));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n14763), .D(n27205));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n14763), .D(n26972));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n14763), .D(n27830));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n14763), .D(n27864));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n14737), .D(n8825[7]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_8_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_3821));
    defparam select_292_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_7_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_3819));
    defparam select_292_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n25404), .S(n25400));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n18422), .S(n18934));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n18424), .S(n18936));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n7_adj_3674), .S(n8_adj_3677));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n18426), .S(n18938));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n7_adj_3673), .S(n25264));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n25408), .S(n25502));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n25412), .S(n25500));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n25414), .S(n25498));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n25416), .S(n25496));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n25418), .S(n25494));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n25420), .S(n25492));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n25422), .S(n25490));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n7_adj_3668), .S(n8_adj_3835));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n7_adj_3667), .S(n8_adj_3836));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_3666), .S(n8_adj_3837));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n7_adj_3665), .S(n8_adj_3838));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n18428), .S(n8_adj_3839));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n25388), .S(n25384));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n25382), .S(n25508));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n25424), .S(n25486));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n7_adj_3663), .S(n8_adj_3840));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n25426), .S(n25484));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n7_adj_3662), .S(n8_adj_3841));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n25428), .S(n25482));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n25430), .S(n25442));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n25432), .S(n25480));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n25434), .S(n25478));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n25378), .S(n25438));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_292_Select_6_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_3817));
    defparam select_292_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_5_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_3816));
    defparam select_292_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_4_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_3815));
    defparam select_292_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_3_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_3814));
    defparam select_292_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i11413_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n15244));
    defparam i11413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11414_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n15245));
    defparam i11414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_292_Select_2_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_3813));
    defparam select_292_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_1_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_3798));
    defparam select_292_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_292_Select_0_i3_2_lut_4_lut (.I0(n18939), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n13616), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_292_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i11415_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n15246));
    defparam i11415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11568_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n15399));
    defparam i11568_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1244 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n26186));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_LUT4 i11569_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n15400));
    defparam i11569_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3842));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_3843));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_18_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n21951), .O(n2_adj_3834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11570_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n15401));
    defparam i11570_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24491_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29226));
    defparam i24491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1245 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[12] [5]), .I3(n26472), .O(n26572));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i24493_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n29225));
    defparam i24493_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n15522), 
            .D(n4040), .R(n26794));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11571_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n15402));
    defparam i11571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11572_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n15403));
    defparam i11572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11573_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n15404));
    defparam i11573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11574_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n15405));
    defparam i11574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11575_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n15406));
    defparam i11575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n13_adj_3844), .D(n14853), 
            .R(n27660));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_75_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3654));   // verilog/coms.v(154[7:23])
    defparam equal_75_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_CARRY add_43_18 (.CI(n21951), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n21952));
    SB_LUT4 equal_76_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3671));   // verilog/coms.v(154[7:23])
    defparam equal_76_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 add_43_17_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n21950), .O(n2_adj_3833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_17 (.CI(n21950), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n21951));
    SB_LUT4 add_43_16_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n21949), .O(n2_adj_3832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n21949), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n21950));
    SB_LUT4 i25128_2_lut_3_lut (.I0(n26785), .I1(n18983), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n26794));
    defparam i25128_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i11560_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n15391));
    defparam i11560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11561_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n15392));
    defparam i11561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11562_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n15393));
    defparam i11562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n14737), .D(n8825[6]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11563_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n15394));
    defparam i11563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11564_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n15395));
    defparam i11564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11565_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n15396));
    defparam i11565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n26605));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i11566_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n15397));
    defparam i11566_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11567_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n15398));
    defparam i11567_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i25157_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n14853));
    defparam i25157_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 add_43_15_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n21948), .O(n2_adj_3830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_15 (.CI(n21948), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n21949));
    SB_LUT4 add_43_14_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n21947), .O(n2_adj_3828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[21] [4]), .I1(n26524), .I2(n26626), 
            .I3(n13867), .O(n12_adj_3789));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1247 (.I0(Kp_23__N_1030), .I1(\data_in_frame[9] [0]), 
            .I2(\data_in_frame[11] [2]), .I3(\data_in_frame[13] [4]), .O(n8_adj_3774));   // verilog/coms.v(73[16:42])
    defparam i3_3_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(\data_in_frame[11] [4]), .I1(n26059), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n6_adj_3773));
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1249 (.I0(n13919), .I1(\data_in_frame[9] [2]), 
            .I2(n14328), .I3(GND_net), .O(n13873));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1249.LUT_INIT = 16'h9696;
    SB_LUT4 i11552_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n15383));
    defparam i11552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11553_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n15384));
    defparam i11553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11554_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n15385));
    defparam i11554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11555_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n15386));
    defparam i11555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_14 (.CI(n21947), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n21948));
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25254 (.I0(byte_transmit_counter[1]), 
            .I1(n29225), .I2(n29226), .I3(byte_transmit_counter[2]), .O(n30334));
    defparam byte_transmit_counter_1__bdd_4_lut_25254.LUT_INIT = 16'he4aa;
    SB_LUT4 i11556_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n15387));
    defparam i11556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n30334_bdd_4_lut (.I0(n30334), .I1(n17_adj_3843), .I2(n16_adj_3842), 
            .I3(byte_transmit_counter[2]), .O(n30337));
    defparam n30334_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11557_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n15388));
    defparam i11557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_11 (.CI(n21944), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n21945));
    SB_LUT4 i11558_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n15389));
    defparam i11558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11559_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n15390));
    defparam i11559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11120_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n14951));
    defparam i11120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n14737), .D(n8825[5]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1250 (.I0(\data_in_frame[9] [4]), .I1(n23686), 
            .I2(n14420), .I3(GND_net), .O(n26059));
    defparam i1_2_lut_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_LUT4 equal_69_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3683));   // verilog/coms.v(154[7:23])
    defparam equal_69_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n14991));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n14737), .D(n8825[4]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_78_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3716));   // verilog/coms.v(154[7:23])
    defparam equal_78_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i11544_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n15375));
    defparam i11544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n14737), .D(n8825[3]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11545_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n15376));
    defparam i11545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11546_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n15377));
    defparam i11546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_13_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n21946), .O(n2_adj_3826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11547_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n15378));
    defparam i11547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n14990));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1251 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [5]), .I3(n26120), .O(n23686));
    defparam i1_3_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_CARRY add_43_13 (.CI(n21946), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n21947));
    SB_LUT4 add_43_12_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n21945), .O(n2_adj_3824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n14989));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11548_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n15379));
    defparam i11548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11549_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n15380));
    defparam i11549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n14988));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11550_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n15381));
    defparam i11550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11551_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n15382));
    defparam i11551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11536_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n15367));
    defparam i11536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11537_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n15368));
    defparam i11537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1252 (.I0(n26110), .I1(n26381), .I2(Kp_23__N_1218), 
            .I3(n13964), .O(n12_adj_3845));
    defparam i5_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n14987));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11401_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n15232));
    defparam i11401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11538_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n15369));
    defparam i11538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11402_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n15233));
    defparam i11402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1253 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n18565), .I3(GND_net), .O(n61_adj_3846));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut_adj_1253.LUT_INIT = 16'hecec;
    SB_LUT4 i11539_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n15370));
    defparam i11539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21610_4_lut (.I0(n26785), .I1(n61_adj_3846), .I2(n26779), 
            .I3(\FRAME_MATCHER.state [0]), .O(n51));
    defparam i21610_4_lut.LUT_INIT = 16'h0545;
    SB_LUT4 i11403_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n15234));
    defparam i11403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(n26323), .I2(\data_in_frame[16] [6]), 
            .I3(\data_in_frame[17] [0]), .O(n46));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11404_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n15235));
    defparam i11404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1254 (.I0(n51), .I1(n18983), .I2(GND_net), .I3(GND_net), 
            .O(n27660));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut_adj_1254.LUT_INIT = 16'h2222;
    SB_LUT4 i11540_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n15371));
    defparam i11540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11541_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n15372));
    defparam i11541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(n16455), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2444 [3]), 
            .O(n15_adj_3847));
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h4474;
    SB_LUT4 i2_3_lut_adj_1256 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n26635));
    defparam i2_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_LUT4 i25057_4_lut (.I0(n51), .I1(n15_adj_3847), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n18983), .O(n13_adj_3844));
    defparam i25057_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 i11542_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n15373));
    defparam i11542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1257 (.I0(\data_in_frame[11] [6]), .I1(n24652), 
            .I2(n10_adj_3771), .I3(\data_in_frame[13] [7]), .O(n26539));
    defparam i5_3_lut_4_lut_adj_1257.LUT_INIT = 16'h9669;
    SB_LUT4 i11405_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n15236));
    defparam i11405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11543_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n15374));
    defparam i11543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11528_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n15359));
    defparam i11528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11529_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n15360));
    defparam i11529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1258 (.I0(n23686), .I1(\data_in_frame[9] [5]), 
            .I2(n13972), .I3(n26059), .O(n24652));
    defparam i1_2_lut_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i11530_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n15361));
    defparam i11530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21701_2_lut (.I0(n18983), .I1(\FRAME_MATCHER.state [3]), .I2(GND_net), 
            .I3(GND_net), .O(n26779));
    defparam i21701_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26043));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1260 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(n26155), .I3(\data_out_frame[10] [2]), .O(n26435));
    defparam i1_2_lut_3_lut_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i23251_2_lut (.I0(n26785), .I1(\FRAME_MATCHER.state [1]), .I2(GND_net), 
            .I3(GND_net), .O(n28339));
    defparam i23251_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1261 (.I0(n26056), .I1(n26289), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[15] [7]), .O(n14665));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26659));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1263 (.I0(\FRAME_MATCHER.state [2]), .I1(n26794), 
            .I2(n28339), .I3(n18565), .O(n15522));
    defparam i1_4_lut_adj_1263.LUT_INIT = 16'hcdcc;
    SB_LUT4 i2_3_lut_adj_1264 (.I0(n14380), .I1(n26659), .I2(n14005), 
            .I3(GND_net), .O(n26067));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1264.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1265 (.I0(n26620), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[15] [1]), .I3(n12058), .O(n26064));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i11406_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n15237));
    defparam i11406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26626));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[15] [0]), .I1(n14297), 
            .I2(GND_net), .I3(GND_net), .O(n26524));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(n26524), .I1(n26626), .I2(n13867), 
            .I3(GND_net), .O(n26053));
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n14986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n14985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n14984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n14983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n14982));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n14981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n14980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n14979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n14978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n14977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n14976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n14975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n14974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n14973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n14972));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11531_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n15362));
    defparam i11531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11532_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n15363));
    defparam i11532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1269 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[9] [3]), .I3(\data_in_frame[9] [5]), .O(n18_adj_3764));
    defparam i1_2_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i11533_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n15364));
    defparam i11533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11407_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25997), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n15238));
    defparam i11407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11534_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n15365));
    defparam i11534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1270 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n26475));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25240 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n30328));
    defparam byte_transmit_counter_0__bdd_4_lut_25240.LUT_INIT = 16'he4aa;
    SB_LUT4 n30328_bdd_4_lut (.I0(n30328), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n30331));
    defparam n30328_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1271 (.I0(\data_in_frame[19] [0]), .I1(n18_adj_3778), 
            .I2(\data_in_frame[18] [6]), .I3(n26584), .O(n20_adj_3848));   // verilog/coms.v(76[16:43])
    defparam i9_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25230 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n30322));
    defparam byte_transmit_counter_0__bdd_4_lut_25230.LUT_INIT = 16'he4aa;
    SB_LUT4 n30322_bdd_4_lut (.I0(n30322), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n30325));
    defparam n30322_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1272 (.I0(n26457), .I1(n12058), .I2(\data_in_frame[16] [4]), 
            .I3(\data_in_frame[21] [2]), .O(n19_adj_3849));   // verilog/coms.v(76[16:43])
    defparam i8_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25235 (.I0(byte_transmit_counter[1]), 
            .I1(n29228), .I2(n29229), .I3(byte_transmit_counter[2]), .O(n30316));
    defparam byte_transmit_counter_1__bdd_4_lut_25235.LUT_INIT = 16'he4aa;
    SB_LUT4 n30316_bdd_4_lut (.I0(n30316), .I1(n17_adj_3750), .I2(n16_adj_3749), 
            .I3(byte_transmit_counter[2]), .O(n30319));
    defparam n30316_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1273 (.I0(\data_in_frame[20] [2]), .I1(n12_adj_3845), 
            .I2(n26560), .I3(\data_in_frame[15] [6]), .O(n27779));
    defparam i6_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25220 (.I0(byte_transmit_counter[1]), 
            .I1(n29231), .I2(n29232), .I3(byte_transmit_counter[2]), .O(n30310));
    defparam byte_transmit_counter_1__bdd_4_lut_25220.LUT_INIT = 16'he4aa;
    SB_LUT4 n30310_bdd_4_lut (.I0(n30310), .I1(n17_adj_3744), .I2(n16_adj_3742), 
            .I3(byte_transmit_counter[2]), .O(n30313));
    defparam n30310_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i23269_4_lut (.I0(\data_in_frame[19] [3]), .I1(n27514), .I2(n8_adj_3792), 
            .I3(\data_in_frame[19] [4]), .O(n28357));
    defparam i23269_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25215 (.I0(byte_transmit_counter[1]), 
            .I1(n29235), .I2(n29236), .I3(byte_transmit_counter[2]), .O(n30304));
    defparam byte_transmit_counter_1__bdd_4_lut_25215.LUT_INIT = 16'he4aa;
    SB_LUT4 n30304_bdd_4_lut (.I0(n30304), .I1(n17_adj_3739), .I2(n16_adj_3738), 
            .I3(byte_transmit_counter[2]), .O(n30307));
    defparam n30304_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1274 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n26336), .I3(GND_net), .O(n6_adj_3850));
    defparam i2_3_lut_adj_1274.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25210 (.I0(byte_transmit_counter[1]), 
            .I1(n29238), .I2(n29239), .I3(byte_transmit_counter[2]), .O(n30298));
    defparam byte_transmit_counter_1__bdd_4_lut_25210.LUT_INIT = 16'he4aa;
    SB_LUT4 n30298_bdd_4_lut (.I0(n30298), .I1(n17_adj_3737), .I2(n16_adj_3736), 
            .I3(byte_transmit_counter[2]), .O(n30301));
    defparam n30298_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1275 (.I0(\data_in_frame[21] [1]), .I1(n26172), 
            .I2(n24249), .I3(n12137), .O(n27142));
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_25205 (.I0(byte_transmit_counter[1]), 
            .I1(n29241), .I2(n29242), .I3(byte_transmit_counter[2]), .O(n30292));
    defparam byte_transmit_counter_1__bdd_4_lut_25205.LUT_INIT = 16'he4aa;
    SB_LUT4 n30292_bdd_4_lut (.I0(n30292), .I1(n17_adj_3735), .I2(n16_adj_3734), 
            .I3(byte_transmit_counter[2]), .O(n30295));
    defparam n30292_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n26310), .I1(n27617), .I2(n10_adj_3782), 
            .I3(n26426), .O(n20_adj_3851));
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h4884;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n14737), .D(n8825[2]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11535_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25990), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n15366));
    defparam i11535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1277 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n26602));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i5_2_lut_4_lut (.I0(n13972), .I1(n13988), .I2(\data_in_frame[9] [7]), 
            .I3(n13877), .O(n18_adj_3762));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1278 (.I0(n11166), .I1(n30), .I2(n13611), 
            .I3(GND_net), .O(n7330));   // verilog/coms.v(238[12:32])
    defparam i1_2_lut_3_lut_adj_1278.LUT_INIT = 16'h0404;
    SB_LUT4 i12625_3_lut_4_lut_4_lut (.I0(n11166), .I1(n30), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n1), .O(n16455));   // verilog/coms.v(238[12:32])
    defparam i12625_3_lut_4_lut_4_lut.LUT_INIT = 16'h0454;
    SB_LUT4 i1_2_lut_3_lut_adj_1279 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n13852));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i11520_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n15351));
    defparam i11520_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1280 (.I0(n23692), .I1(n26110), .I2(\data_in_frame[17] [5]), 
            .I3(\data_in_frame[19] [6]), .O(n26336));
    defparam i1_2_lut_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i11521_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n15352));
    defparam i11521_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1281 (.I0(\FRAME_MATCHER.state [31]), .I1(n11123), 
            .I2(n3_adj_3658), .I3(n4_adj_3775), .O(n25378));
    defparam i1_4_lut_adj_1281.LUT_INIT = 16'ha8a0;
    SB_LUT4 i11522_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n15353));
    defparam i11522_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11523_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n15354));
    defparam i11523_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut_4_lut_adj_1282 (.I0(n13919), .I1(n26090), .I2(n10_adj_3757), 
            .I3(\data_in_frame[13] [3]), .O(n23700));
    defparam i5_3_lut_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_CARRY add_43_12 (.CI(n21945), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n21946));
    SB_LUT4 i11524_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n15355));
    defparam i11524_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1283 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[4] [0]), .O(n6_adj_3653));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i11525_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n15356));
    defparam i11525_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11526_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n15357));
    defparam i11526_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11527_3_lut_4_lut (.I0(n18978), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n15358));
    defparam i11527_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1284 (.I0(\data_in_frame[11] [3]), .I1(n13919), 
            .I2(n8_adj_3652), .I3(\data_in_frame[9] [1]), .O(n26289));
    defparam i2_3_lut_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1285 (.I0(\data_in_frame[2] [4]), .I1(n26333), 
            .I2(n10_adj_3751), .I3(n14677), .O(n14420));
    defparam i5_3_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1286 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [0]), .I3(GND_net), .O(n10_adj_3746));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1287 (.I0(\data_in_frame[18] [3]), .I1(n27118), 
            .I2(n8_adj_3784), .I3(n26310), .O(n18_adj_3852));
    defparam i2_4_lut_adj_1287.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1288 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18435), .O(n25997));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1288.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1289 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n18435), .O(n25981));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1289.LUT_INIT = 16'hefff;
    SB_LUT4 add_43_11_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n21944), .O(n2_adj_3822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(n11166), .I1(n1), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n3963));
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h1010;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n21973), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n21972), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_9 (.CI(n21942), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n21943));
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[12] [4]), .I1(n26093), 
            .I2(\data_out_frame[12] [2]), .I3(\data_out_frame[12] [1]), 
            .O(n16_adj_3585));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11512_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n15343));
    defparam i11512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(n3_adj_3601), .I1(n12033), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[8] [1]), .O(n14005));
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_8 (.CI(n21972), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n21973));
    SB_LUT4 i11513_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n15344));
    defparam i11513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n30906));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_10_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n21943), .O(n2_adj_3820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n30907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n15436));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n15435));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n15434));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11514_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n15345));
    defparam i11514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n15433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n15432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n15431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n15430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n15429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n15428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n15427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n15426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n15425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n15424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n15423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n15422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n15421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n15420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n15419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n15418));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n15417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n15416));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i215_2_lut (.I0(\FRAME_MATCHER.state [26]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3841));
    defparam i215_2_lut.LUT_INIT = 16'h8888;
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n15415));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11515_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n15346));
    defparam i11515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n15414));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(\data_out_frame[17] [5]), .I1(n13814), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n26050));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1293 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [3]), .O(n14396));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n15413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n15412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n15411));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n21971), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n15410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n15409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n15408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n15407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n15406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n15405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n15404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n15403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n15402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n15401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n15400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n15399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n15398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n15397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n15396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n15395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n15394));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1294 (.I0(\data_out_frame[17] [5]), .I1(n13814), 
            .I2(n24531), .I3(GND_net), .O(n26638));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n15393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n15392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n15391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n15390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n15389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n15388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n15387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n15386));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i204_2_lut (.I0(\FRAME_MATCHER.state [24]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3840));
    defparam i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15155_2_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n21466), .O(n18983));
    defparam i15155_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n15385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n15384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n15383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n15382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n15381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n15380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n15379));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n15378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n15377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n15376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n15375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n15374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n15373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n15372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n15371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n15370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n15369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n15368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n15367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n15366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n15365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n15364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n15363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n15362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n15361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n15360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n15359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n15358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n15357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n15356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n15355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n15354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n15353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n15352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n15351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n15350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n15349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n15348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n15347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n15346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n15345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n15344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n15343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n15342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n15341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n15340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n15339));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n15338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n15337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n15336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n15335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n15334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n15333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n15332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n15331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n15330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n15329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n15328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n15327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n15326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n15325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n15324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n15323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n15322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n15321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n15320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n15319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n15318));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n15317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n15316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n15315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n15314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n15313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n15312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n15311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n15310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n15309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n15308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n15307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n15306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n15305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n15304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n15303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n15302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n15301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n15300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n15299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n15298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n15297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n15296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n15295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n15294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n15293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n15292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n15291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n15290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n15289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n15288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n15287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n15286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n15285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n15284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n15283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n15282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n15281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n15280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n15279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n15278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n15277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n15276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n15275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n15274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n15273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n15272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n15271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n15270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n15269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n15268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n15267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n15266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n15265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n15264));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n15263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n15262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n15261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n15260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n15259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n15258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n15257));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n15256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n15255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n15254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n15253));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n15252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n15251));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n15250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n15249));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n15248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n15247));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1295 (.I0(n13919), .I1(n26090), .I2(n10_adj_3726), 
            .I3(\data_in_frame[11] [6]), .O(n26310));
    defparam i5_3_lut_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i11516_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n15347));
    defparam i11516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(n14153), .I1(Kp_23__N_888), .I2(n26283), 
            .I3(GND_net), .O(n26402));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[6] [1]), 
            .I2(n26034), .I3(GND_net), .O(Kp_23__N_888));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1298 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n13625), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_3715));
    defparam i1_3_lut_4_lut_adj_1298.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(n28121), .I1(n23768), .I2(n26381), 
            .I3(\data_in_frame[20] [3]), .O(n19_adj_3853));
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'h8228;
    SB_LUT4 i201_2_lut (.I0(\FRAME_MATCHER.state [20]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3839));
    defparam i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21603_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n28307), 
            .I2(n3303), .I3(GND_net), .O(n26678));
    defparam i21603_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i220_2_lut (.I0(\FRAME_MATCHER.state [19]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3838));
    defparam i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23223_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n21466), .I3(\FRAME_MATCHER.state [1]), .O(n28307));   // verilog/coms.v(212[5:16])
    defparam i23223_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i223_2_lut (.I0(\FRAME_MATCHER.state [18]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3837));
    defparam i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11517_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n15348));
    defparam i11517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1300 (.I0(\data_in_frame[9] [3]), .I1(n14328), 
            .I2(n14420), .I3(\data_in_frame[11] [4]), .O(n26056));
    defparam i1_2_lut_3_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i11518_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n15349));
    defparam i11518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i212_2_lut (.I0(\FRAME_MATCHER.state [17]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3836));
    defparam i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11519_3_lut_4_lut (.I0(n8_adj_3622), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n15350));
    defparam i11519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[7] [5]), .I3(n26599), .O(n18_adj_3854));   // verilog/coms.v(73[16:27])
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17713_4_lut (.I0(n184), .I1(n26678), .I2(n8634), .I3(n2254), 
            .O(n194));
    defparam i17713_4_lut.LUT_INIT = 16'hfaba;
    SB_LUT4 i11504_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n15335));
    defparam i11504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11505_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n15336));
    defparam i11505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11506_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n15337));
    defparam i11506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11507_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n15338));
    defparam i11507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11508_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n15339));
    defparam i11508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25225 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n30286));
    defparam byte_transmit_counter_0__bdd_4_lut_25225.LUT_INIT = 16'he4aa;
    SB_LUT4 i207_2_lut (.I0(\FRAME_MATCHER.state [16]), .I1(n194), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3835));
    defparam i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1301 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[6] [5]), .O(n26629));
    defparam i1_2_lut_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 n30286_bdd_4_lut (.I0(n30286), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n30289));
    defparam n30286_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1302 (.I0(n27142), .I1(\data_in_frame[20] [0]), 
            .I2(n6_adj_3850), .I3(n26274), .O(n17_adj_3855));
    defparam i1_4_lut_adj_1302.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25196 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n30280));
    defparam byte_transmit_counter_0__bdd_4_lut_25196.LUT_INIT = 16'he4aa;
    SB_LUT4 n30280_bdd_4_lut (.I0(n30280), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n30283));
    defparam n30280_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14613_2_lut_2_lut_3_lut (.I0(n18939), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n18435));
    defparam i14613_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_2_lut_3_lut_adj_1303 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[4] [5]), 
            .I2(\data_in_frame[6] [1]), .I3(GND_net), .O(n10_adj_3703));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n15246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n15245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n15244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n15243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n15242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n15241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n15240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n15239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n15238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n15237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n15236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n15235));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n15234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n15233));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n15232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n15231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n15230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n15229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n15228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n15227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n15226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n15225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n15224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n15223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n15222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n15221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n15220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n15219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n15218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n15217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n15216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n15215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n15214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n15213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n15212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n15211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n15210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n15209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n15208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n15207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n15206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n15205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n15204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n15203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n15202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n15201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n15200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n15199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n15198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n15197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n15196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n15195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n15194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n15193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n15192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n15191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n15190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n15189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n15188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n15187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n15186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n15185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n15184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n15183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n15182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n15181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n15180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n15179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n15178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n15177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n15176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n15175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n15174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n15173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n15172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n15171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n15170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n15169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n15168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n15167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n15166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n15165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n15164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n15163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n15162));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1304 (.I0(n13988), .I1(\data_in_frame[7] [7]), 
            .I2(n14153), .I3(n26284), .O(n5_adj_3696));
    defparam i1_3_lut_4_lut_adj_1304.LUT_INIT = 16'h7dd7;
    SB_LUT4 i8_4_lut_adj_1305 (.I0(\data_in_frame[21] [0]), .I1(n27002), 
            .I2(n6_adj_3786), .I3(n26323), .O(n24));
    defparam i8_4_lut_adj_1305.LUT_INIT = 16'h4884;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_25191 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n30274));
    defparam byte_transmit_counter_0__bdd_4_lut_25191.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1306 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n21466), .O(n13616));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1306.LUT_INIT = 16'hfffe;
    SB_LUT4 n30274_bdd_4_lut (.I0(n30274), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n30277));
    defparam n30274_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1307 (.I0(n28125), .I1(\data_in_frame[19] [0]), 
            .I2(n4_adj_3791), .I3(n24249), .O(n23));
    defparam i7_4_lut_adj_1307.LUT_INIT = 16'h2882;
    SB_LUT4 i11509_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n15340));
    defparam i11509_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11510_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n15341));
    defparam i11510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n13892), .I1(n13867), .I2(\data_in_frame[8] [0]), 
            .I3(\data_in_frame[8] [1]), .O(n10_adj_3600));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1308 (.I0(n63), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n53), .I3(n62), .O(\FRAME_MATCHER.state_31__N_2380[2] ));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_4_lut_adj_1308.LUT_INIT = 16'h8a0a;
    SB_LUT4 i11511_3_lut_4_lut (.I0(n8_adj_3654), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n15342));
    defparam i11511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1309 (.I0(n11119), .I1(n11125), .I2(n28307), 
            .I3(n13616), .O(n10_adj_3684));
    defparam i1_4_lut_adj_1309.LUT_INIT = 16'h0ace;
    SB_LUT4 i1_2_lut_3_lut_adj_1310 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n26484));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1311 (.I0(\data_in_frame[8] [7]), .I1(n10_adj_3649), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[4] [5]), .O(n8_adj_3652));   // verilog/coms.v(166[9:87])
    defparam i5_3_lut_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i11496_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n15327));
    defparam i11496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n14737), .D(n8825[1]), .R(n14863));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i25154_3_lut_4_lut (.I0(n63_adj_3), .I1(tx_active), .I2(r_SM_Main_2__N_3336[0]), 
            .I3(n13651), .O(n14737));
    defparam i25154_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_CARRY add_43_10 (.CI(n21943), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n21944));
    SB_LUT4 i2_3_lut_4_lut_adj_1312 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[23] [4]), 
            .I2(n23733), .I3(\data_out_frame[19] [4]), .O(n26514));
    defparam i2_3_lut_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(n771), .I1(n8634), .I2(GND_net), .I3(GND_net), 
            .O(n11125));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h4444;
    SB_LUT4 i11497_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n15328));
    defparam i11497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(n4452), .I1(n8634), .I2(GND_net), .I3(GND_net), 
            .O(n11123));   // verilog/coms.v(259[6] 261[9])
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h4444;
    SB_LUT4 i11498_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n15329));
    defparam i11498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1315 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[14] [5]), .I3(GND_net), .O(n6_adj_3611));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n15161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n15160));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1316 (.I0(n8634), .I1(n2254), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_3676));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n15159));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\data_in_frame[0] [5]), .I1(n26028), 
            .I2(GND_net), .I3(GND_net), .O(n13805));
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_LUT4 i39_4_lut (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[1] [7]), .I3(n13805), .O(n28_adj_3856));
    defparam i39_4_lut.LUT_INIT = 16'h1008;
    SB_LUT4 i11499_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n15330));
    defparam i11499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n15158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n15157));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1318 (.I0(n13852), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[2] [3]), .I3(n28_adj_3856), .O(n18_adj_3857));
    defparam i7_4_lut_adj_1318.LUT_INIT = 16'h0100;
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(n25896), .I3(GND_net), .O(n17_adj_3858));
    defparam i6_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i11500_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n15331));
    defparam i11500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1319 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [6]), .O(n19_adj_3859));
    defparam i8_4_lut_adj_1319.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_1320 (.I0(\data_in_frame[1] [2]), .I1(n19_adj_3859), 
            .I2(n17_adj_3858), .I3(n18_adj_3857), .O(n6_adj_3860));
    defparam i1_4_lut_adj_1320.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut_adj_1321 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n6_adj_3860), .O(\FRAME_MATCHER.state_31__N_2444 [3]));
    defparam i4_4_lut_adj_1321.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_adj_1322 (.I0(n14116), .I1(\data_out_frame[14] [3]), 
            .I2(n24584), .I3(\data_out_frame[16] [4]), .O(n26463));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut_adj_1322.LUT_INIT = 16'h9669;
    SB_LUT4 i11501_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n15332));
    defparam i11501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(\data_out_frame[16] [6]), .I1(n26300), 
            .I2(n26364), .I3(GND_net), .O(n26590));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(n8634), .I1(n3303), .I2(GND_net), .I3(GND_net), 
            .O(n11119));   // verilog/coms.v(142[7:84])
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h2222;
    SB_LUT4 i11502_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n15333));
    defparam i11502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11503_3_lut_4_lut (.I0(n8_adj_3671), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n15334));
    defparam i11503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1325 (.I0(n26245), .I1(n26348), .I2(\data_out_frame[17] [2]), 
            .I3(n23733), .O(n26644));
    defparam i1_2_lut_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1326 (.I0(\data_out_frame[6] [2]), .I1(n26611), 
            .I2(\data_out_frame[6] [1]), .I3(n26155), .O(n14511));
    defparam i1_2_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1327 (.I0(n26245), .I1(n26348), .I2(\data_out_frame[17] [2]), 
            .I3(\data_out_frame[19] [3]), .O(n24639));
    defparam i1_2_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1328 (.I0(n184), .I1(n3_adj_3658), .I2(n44), 
            .I3(GND_net), .O(n27904));
    defparam i2_3_lut_adj_1328.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1329 (.I0(\FRAME_MATCHER.state_31__N_2444 [3]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n13621), .I3(n27904), .O(n25400));
    defparam i1_4_lut_adj_1329.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26490));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i11488_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n15319));
    defparam i11488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11489_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n15320));
    defparam i11489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(n26611), .I3(GND_net), .O(n6_adj_3608));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i11490_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n15321));
    defparam i11490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1332 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[10] [1]), 
            .I2(n26481), .I3(GND_net), .O(n26093));
    defparam i1_2_lut_3_lut_adj_1332.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1333 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [6]), .I3(\data_out_frame[8] [2]), .O(n26472));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1334 (.I0(n13686), .I1(n26265), .I2(\data_out_frame[23] [1]), 
            .I3(n23772), .O(n26972));
    defparam i3_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1335 (.I0(n28357), .I1(n27779), .I2(n19_adj_3849), 
            .I3(n20_adj_3848), .O(n27));
    defparam i11_4_lut_adj_1335.LUT_INIT = 16'h4004;
    SB_LUT4 i2_3_lut_adj_1336 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(n24558), .I3(GND_net), .O(n27205));
    defparam i2_3_lut_adj_1336.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1337 (.I0(n14075), .I1(n26393), .I2(n13751), 
            .I3(n14487), .O(n26890));
    defparam i3_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_out_frame[25] [1]), .I1(n24046), 
            .I2(GND_net), .I3(GND_net), .O(n11578));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(n24615), .I1(n26390), .I2(GND_net), 
            .I3(GND_net), .O(n26392));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1340 (.I0(n26551), .I1(n13747), .I2(n26268), 
            .I3(n24554), .O(n14_adj_3861));
    defparam i6_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1341 (.I0(\data_out_frame[24] [7]), .I1(n14_adj_3861), 
            .I2(n10_adj_3808), .I3(\data_out_frame[18] [1]), .O(n24615));
    defparam i7_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(n24615), .I1(n24598), .I2(GND_net), 
            .I3(GND_net), .O(n26393));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(n14056), .I1(n26070), .I2(GND_net), 
            .I3(GND_net), .O(n2122));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i11491_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n15322));
    defparam i11491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11492_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n15323));
    defparam i11492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1344 (.I0(n14243), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[17] [2]), .I3(n23731), .O(n23733));
    defparam i2_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i11493_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n15324));
    defparam i11493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1345 (.I0(n13747), .I1(n26304), .I2(\data_out_frame[20] [4]), 
            .I3(n24656), .O(n24598));
    defparam i3_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 i11494_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n15325));
    defparam i11494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[23] [0]), .I1(n23772), 
            .I2(GND_net), .I3(GND_net), .O(n26351));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1347 (.I0(\data_out_frame[23] [2]), .I1(n26351), 
            .I2(n24598), .I3(n13751), .O(n24558));
    defparam i3_4_lut_adj_1347.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[23] [4]), .I1(n26343), 
            .I2(GND_net), .I3(GND_net), .O(n23804));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1349 (.I0(\data_out_frame[23] [5]), .I1(n24639), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3862));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1349.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1350 (.I0(n2122), .I1(\data_out_frame[23] [4]), 
            .I2(n24641), .I3(n6_adj_3862), .O(n2406));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1350.LUT_INIT = 16'h9669;
    SB_LUT4 i11495_3_lut_4_lut (.I0(n8_adj_3683), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n15326));
    defparam i11495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(n2406), .I1(n24180), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3863));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(n23804), .I1(n2400), .I2(n24558), .I3(n6_adj_3863), 
            .O(n26390));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1353 (.I0(\data_out_frame[25] [0]), .I1(n26393), 
            .I2(n26262), .I3(n11926), .O(n24046));
    defparam i3_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i11480_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n15311));
    defparam i11480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1354 (.I0(n24046), .I1(n26390), .I2(GND_net), 
            .I3(GND_net), .O(n26391));
    defparam i1_2_lut_adj_1354.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n13686));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n14075));
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26262));
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1358 (.I0(\data_out_frame[20] [6]), .I1(n26228), 
            .I2(n1927), .I3(n13369), .O(n24251));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1359 (.I0(n26070), .I1(n24554), .I2(n24251), 
            .I3(GND_net), .O(n23696));
    defparam i2_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1360 (.I0(n26396), .I1(n24550), .I2(n26248), 
            .I3(\data_out_frame[19] [3]), .O(n14_adj_3864));
    defparam i6_4_lut_adj_1360.LUT_INIT = 16'h9669;
    SB_LUT4 i11481_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n15312));
    defparam i11481_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1361 (.I0(n13308), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3865));
    defparam i1_2_lut_adj_1361.LUT_INIT = 16'h6666;
    SB_LUT4 i11482_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n15313));
    defparam i11482_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1362 (.I0(n9_adj_3865), .I1(n14_adj_3864), .I2(n26307), 
            .I3(n24582), .O(n24546));
    defparam i7_4_lut_adj_1362.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1363 (.I0(n26255), .I1(n26638), .I2(GND_net), 
            .I3(GND_net), .O(n26530));
    defparam i1_2_lut_adj_1363.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(n13751), .I1(n14056), .I2(n26070), 
            .I3(\data_out_frame[23] [3]), .O(n26265));
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(n26572), .I3(GND_net), .O(n6_adj_3605));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1366 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [4]), 
            .I2(n26578), .I3(n24546), .O(n18_adj_3866));
    defparam i7_4_lut_adj_1366.LUT_INIT = 16'h9669;
    SB_LUT4 i11483_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n15314));
    defparam i11483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_2_lut_adj_1367 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3867));
    defparam i5_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1368 (.I0(\data_out_frame[19] [0]), .I1(n18_adj_3866), 
            .I2(n24584), .I3(n26644), .O(n20_adj_3868));
    defparam i9_4_lut_adj_1368.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1369 (.I0(n26590), .I1(n20_adj_3868), .I2(n16_adj_3867), 
            .I3(n26530), .O(n24544));
    defparam i10_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1370 (.I0(n24607), .I1(n26530), .I2(\data_out_frame[16] [5]), 
            .I3(GND_net), .O(n27626));
    defparam i2_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 i11484_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n15315));
    defparam i11484_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1371 (.I0(\data_out_frame[20] [7]), .I1(n26644), 
            .I2(n24546), .I3(n27626), .O(n24554));
    defparam i3_4_lut_adj_1371.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(n24554), .I1(n24544), .I2(GND_net), 
            .I3(GND_net), .O(n23715));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n15156));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11485_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n15316));
    defparam i11485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26268));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1374 (.I0(\data_out_frame[23] [3]), .I1(n24641), 
            .I2(n14056), .I3(n23715), .O(n26343));
    defparam i1_4_lut_adj_1374.LUT_INIT = 16'h9669;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n16_adj_3604));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11486_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n15317));
    defparam i11486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11487_3_lut_4_lut (.I0(n8_adj_3716), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n15318));
    defparam i11487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_2_lut (.I0(n13814), .I1(\data_out_frame[16] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3869));
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1375 (.I0(n25_adj_3869), .I1(\data_out_frame[14] [7]), 
            .I2(n24574), .I3(n26566), .O(n30_adj_3870));
    defparam i13_4_lut_adj_1375.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n15155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n15154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n15153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n15152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n15151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n15150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n15149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n15148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n15147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n15146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n15145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n15144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n15143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n15142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n15141));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n15140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n15139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n15138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n15137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n15136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n15135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n15134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n15133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n15132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n15131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n15130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n15129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n15128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n15127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n15126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n15125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n15124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n15123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n15122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n15121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n15120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n15119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n15118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n15117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n15116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n15115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n15114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n15113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n15112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n15111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n15110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n15109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n15108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n15107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n15106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n15105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n15104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n15103));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11472_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n15303));
    defparam i11472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n14953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n14952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n14951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n14950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n15102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n15101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n15100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n15099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n15098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n15097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n15096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n14949));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11473_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n15304));
    defparam i11473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n14948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n14947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n15095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n15094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n15093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n15092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n15091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n15090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n15089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n15088));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1376 (.I0(n26234), .I1(n23989), .I2(n24580), 
            .I3(n26563), .O(n28_adj_3871));
    defparam i11_4_lut_adj_1376.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n15087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n15086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n15085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n15084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n15083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n15082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n15081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n15080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n15079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n15078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n15077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n15076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n15075));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1377 (.I0(n26378), .I1(n26126), .I2(n26245), 
            .I3(n26025), .O(n29_adj_3872));
    defparam i12_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1378 (.I0(n26104), .I1(\data_out_frame[14] [6]), 
            .I2(n26319), .I3(n26384), .O(n27_adj_3873));
    defparam i10_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1379 (.I0(n27_adj_3873), .I1(n29_adj_3872), .I2(n28_adj_3871), 
            .I3(n30_adj_3870), .O(n26255));
    defparam i16_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i11474_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n15305));
    defparam i11474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_out_frame[23] [0]), .I1(\data_out_frame[23] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14487));
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 i11475_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n15306));
    defparam i11475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11476_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n15307));
    defparam i11476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut_adj_1381 (.I0(n26343), .I1(n26259), .I2(n26268), 
            .I3(n26248), .O(n42_adj_3874));
    defparam i17_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n26037));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1383 (.I0(n24609), .I1(n26271), .I2(n14487), 
            .I3(n26255), .O(n40_adj_3875));
    defparam i15_4_lut_adj_1383.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_1384 (.I0(n23696), .I1(\data_out_frame[18] [6]), 
            .I2(n24251), .I3(\data_out_frame[23] [2]), .O(n41_adj_3876));
    defparam i16_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1385 (.I0(n26340), .I1(n14171), .I2(n26463), 
            .I3(n26262), .O(n39_adj_3877));
    defparam i14_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1386 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(n13852), .I3(n26175), .O(n14153));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1387 (.I0(n26050), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[20] [0]), .I3(\data_out_frame[20] [5]), 
            .O(n43_adj_3878));
    defparam i18_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i11477_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n15308));
    defparam i11477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23_4_lut (.I0(n39_adj_3877), .I1(n41_adj_3876), .I2(n40_adj_3875), 
            .I3(n42_adj_3874), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11478_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n15309));
    defparam i11478_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(n26186), .I3(\data_out_frame[10] [5]), .O(n14111));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1389 (.I0(n43_adj_3878), .I1(n24544), .I2(n38), 
            .I3(\data_out_frame[20] [6]), .O(n47));
    defparam i22_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1390 (.I0(n47), .I1(n8_adj_3681), .I2(\data_out_frame[25] [5]), 
            .I3(n48), .O(n24180));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1391 (.I0(n24639), .I1(\data_out_frame[25] [0]), 
            .I2(n14056), .I3(n24180), .O(n18_adj_3879));
    defparam i7_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1392 (.I0(\data_out_frame[23] [5]), .I1(n18_adj_3879), 
            .I2(\data_out_frame[20] [3]), .I3(n26405), .O(n20_adj_3880));
    defparam i9_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1393 (.I0(n13_adj_3881), .I1(n20_adj_3880), .I2(n24656), 
            .I3(\data_out_frame[24] [5]), .O(n27278));
    defparam i10_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n14211));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'h9696;
    SB_LUT4 i11479_3_lut_4_lut (.I0(n8_adj_3766), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n15310));
    defparam i11479_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n15074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n15073));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26259));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h6666;
    SB_CARRY add_3971_7 (.CI(n21971), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n21972));
    SB_LUT4 i2_2_lut_adj_1396 (.I0(\data_out_frame[20] [3]), .I1(n13814), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3882));
    defparam i2_2_lut_adj_1396.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1397 (.I0(n7_adj_3882), .I1(n14524), .I2(n24656), 
            .I3(\data_out_frame[20] [2]), .O(n11926));
    defparam i4_4_lut_adj_1397.LUT_INIT = 16'h9669;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n21970), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_43_9_lut (.I0(n1656), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n21942), .O(n2_adj_3818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n15072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n15071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n15070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n15069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n15068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n15067));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_6 (.CI(n21970), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n21971));
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n15066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n14941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n15065));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1398 (.I0(n11926), .I1(n26259), .I2(n28011), 
            .I3(GND_net), .O(n26852));
    defparam i2_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n21969), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1399 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26248));
    defparam i1_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1400 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[8] [7]), .O(n11797));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n26107));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(\data_out_frame[18] [3]), .I1(n26408), 
            .I2(GND_net), .I3(GND_net), .O(n13747));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1403 (.I0(\data_out_frame[17] [7]), .I1(n13933), 
            .I2(\data_out_frame[17] [6]), .I3(GND_net), .O(n26234));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_1404 (.I0(n17_adj_3855), .I1(n19_adj_3853), .I2(n18_adj_3852), 
            .I3(n20_adj_3851), .O(n29));
    defparam i13_4_lut_adj_1404.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[24] [0]), 
            .I2(n14056), .I3(\data_out_frame[23] [7]), .O(n6_adj_3590));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1406 (.I0(\data_out_frame[15] [6]), .I1(n26234), 
            .I2(n14337), .I3(\data_out_frame[18] [0]), .O(n14524));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(\data_out_frame[17] [3]), .I1(n23741), 
            .I2(n24531), .I3(\data_out_frame[17] [4]), .O(n13308));
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n14171));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1409 (.I0(\data_out_frame[24] [4]), .I1(n14171), 
            .I2(n26989), .I3(n26545), .O(n16_adj_3883));
    defparam i6_4_lut_adj_1409.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1410 (.I0(n26405), .I1(n14524), .I2(n13767), 
            .I3(\data_out_frame[24] [3]), .O(n17_adj_3884));
    defparam i7_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1411 (.I0(n17_adj_3884), .I1(n24609), .I2(n16_adj_3883), 
            .I3(n26248), .O(n27684));
    defparam i9_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(n14412), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26563));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(n23785), .I3(n26348), .O(n24550));
    defparam i2_3_lut_4_lut_adj_1413.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1414 (.I0(n11807), .I1(n1445), .I2(\data_out_frame[11] [3]), 
            .I3(\data_out_frame[11] [4]), .O(n26158));
    defparam i2_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[13] [3]), .I3(GND_net), .O(n26469));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1416 (.I0(n24654), .I1(n26319), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n1927));
    defparam i2_3_lut_adj_1416.LUT_INIT = 16'h9696;
    SB_LUT4 i11464_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n15295));
    defparam i11464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11465_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n15296));
    defparam i11465_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1417 (.I0(n26123), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[13] [4]), .I3(n26478), .O(n10_adj_3885));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1418 (.I0(\data_out_frame[8] [7]), .I1(n10_adj_3885), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n13933));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1419 (.I0(n26280), .I1(n27058), .I2(n13933), 
            .I3(GND_net), .O(n26411));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1419.LUT_INIT = 16'h6969;
    SB_LUT4 i11466_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n15297));
    defparam i11466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1420 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[14] [0]), .I3(GND_net), .O(n14668));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1420.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [0]), 
            .I2(n26141), .I3(GND_net), .O(n6_adj_3588));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n15064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n15063));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1422 (.I0(n26638), .I1(\data_out_frame[14] [3]), 
            .I2(n26411), .I3(n14116), .O(n14_adj_3886));
    defparam i6_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1423 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(n13852), .I3(\data_in_frame[4] [4]), .O(n26502));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n15062));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1424 (.I0(n9_adj_3785), .I1(n14_adj_3886), .I2(n26566), 
            .I3(n24584), .O(n26989));
    defparam i7_4_lut_adj_1424.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n15061));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1425 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n26141));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1425.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n15060));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1426 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [5]), 
            .I2(\data_out_frame[14] [3]), .I3(\data_out_frame[14] [1]), 
            .O(n26100));
    defparam i2_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n15059));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\data_out_frame[13] [5]), .I1(n26158), 
            .I2(GND_net), .I3(GND_net), .O(n14337));
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n15058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n15057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n15056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n15055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n15054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n15053));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11467_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n15298));
    defparam i11467_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1428 (.I0(\data_out_frame[16] [3]), .I1(n26569), 
            .I2(n14116), .I3(GND_net), .O(n26025));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1429 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n10_adj_3587));
    defparam i2_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(n13756), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[6] [7]), .O(n26242));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1431 (.I0(n13369), .I1(\data_out_frame[18] [3]), 
            .I2(n26408), .I3(n14491), .O(n26405));
    defparam i1_2_lut_3_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(n26280), .I1(n24594), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3887));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i11468_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n15299));
    defparam i11468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11469_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n15300));
    defparam i11469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11470_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n15301));
    defparam i11470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1433 (.I0(n14337), .I1(\data_out_frame[17] [7]), 
            .I2(n4_adj_3887), .I3(\data_out_frame[15] [7]), .O(n26551));
    defparam i2_4_lut_adj_1433.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1434 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[19] [7]), 
            .I2(n26989), .I3(GND_net), .O(n13_adj_3881));
    defparam i2_3_lut_adj_1434.LUT_INIT = 16'h6969;
    SB_LUT4 i11471_3_lut_4_lut (.I0(n8_adj_3713), .I1(n25981), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n15302));
    defparam i11471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1435 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26228));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1435.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1436 (.I0(\data_out_frame[12] [0]), .I1(n26148), 
            .I2(\data_out_frame[13] [7]), .I3(n14412), .O(n24142));
    defparam i3_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n15052));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1437 (.I0(n24142), .I1(n26100), .I2(GND_net), 
            .I3(GND_net), .O(n26578));
    defparam i1_2_lut_adj_1437.LUT_INIT = 16'h6666;
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n15051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n15050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n15049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n15048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n15047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n15046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n15045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n15044));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1438 (.I0(n26107), .I1(n26469), .I2(n23749), 
            .I3(\data_out_frame[13] [6]), .O(n12_adj_3888));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n15043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n15042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n15041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n15040));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1439 (.I0(\data_out_frame[13] [7]), .I1(n12_adj_3888), 
            .I2(n26572), .I3(\data_out_frame[13] [5]), .O(n23989));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n15039));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(\data_out_frame[11] [5]), .I1(n13756), 
            .I2(n26536), .I3(\data_out_frame[6] [7]), .O(n14412));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n15038));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1441 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(n10), .I3(\data_out_frame[10] [7]), .O(n26313));
    defparam i5_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(n23785), .I1(\data_out_frame[12] [4]), 
            .I2(n14216), .I3(GND_net), .O(n26349));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1443 (.I0(n24641), .I1(n26050), .I2(\data_out_frame[19] [6]), 
            .I3(n14243), .O(n26396));
    defparam i1_2_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1444 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3889));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_adj_1445 (.I0(\data_out_frame[16] [6]), .I1(n23731), 
            .I2(\data_out_frame[17] [0]), .I3(\data_out_frame[17] [1]), 
            .O(n6_adj_3582));
    defparam i2_2_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1446 (.I0(n13906), .I1(\data_out_frame[16] [2]), 
            .I2(n7_adj_3889), .I3(n8_adj_3776), .O(n26569));
    defparam i2_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1447 (.I0(n24142), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26319));
    defparam i1_2_lut_adj_1447.LUT_INIT = 16'h6666;
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n15037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n15036));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [4]), 
            .I2(n24594), .I3(n26326), .O(n26545));
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'h9669;
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n15035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n15034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n15033));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_1449 (.I0(\data_out_frame[15] [7]), .I1(n26596), 
            .I2(n26093), .I3(n26300), .O(n21_adj_3890));
    defparam i8_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n15032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n15031));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_3_lut_adj_1450 (.I0(n23989), .I1(\data_out_frame[16] [1]), 
            .I2(n26578), .I3(GND_net), .O(n20_adj_3891));
    defparam i7_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n15030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n15029));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[17] [4]), 
            .I2(n24594), .I3(GND_net), .O(n24574));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h6969;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n15028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n15027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n15026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n15025));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1452 (.I0(n21_adj_3890), .I1(n26349), .I2(n18_adj_3854), 
            .I3(n26647), .O(n24_adj_3892));
    defparam i11_4_lut_adj_1452.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n15024));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11456_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n15287));
    defparam i11456_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12_4_lut_adj_1453 (.I0(n26096), .I1(n24_adj_3892), .I2(n20_adj_3891), 
            .I3(n26037), .O(n27058));
    defparam i12_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1454 (.I0(n26084), .I1(n26228), .I2(\data_out_frame[18] [2]), 
            .I3(GND_net), .O(n14491));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n15023));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1455 (.I0(n27058), .I1(n26319), .I2(n26569), 
            .I3(n26429), .O(n26408));
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h9669;
    SB_LUT4 i11457_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n15288));
    defparam i11457_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11458_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n15289));
    defparam i11458_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1456 (.I0(\data_out_frame[19] [7]), .I1(n13814), 
            .I2(GND_net), .I3(GND_net), .O(n13767));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1457 (.I0(n14243), .I1(n24531), .I2(GND_net), 
            .I3(GND_net), .O(n24580));
    defparam i1_2_lut_adj_1457.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n15022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n15021));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1458 (.I0(\data_out_frame[24] [3]), .I1(n26197), 
            .I2(\data_out_frame[24] [2]), .I3(n26511), .O(n26271));
    defparam i3_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n15020));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11459_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n15290));
    defparam i11459_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n15019));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_3_lut_adj_1459 (.I0(n13_adj_3881), .I1(n26551), .I2(n13369), 
            .I3(GND_net), .O(n18_adj_3893));
    defparam i7_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n15018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n15017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n15016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n15015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n15014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n15013));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i9_4_lut_adj_1460 (.I0(n24580), .I1(n18_adj_3893), .I2(n26326), 
            .I3(n13767), .O(n20));
    defparam i9_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n15012));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11460_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n15291));
    defparam i11460_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n15011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n15010));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11461_3_lut_4_lut (.I0(n18978), .I1(n25997), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n15292));
    defparam i11461_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1461 (.I0(\data_out_frame[11] [3]), .I1(n26487), 
            .I2(n10), .I3(\data_out_frame[10] [7]), .O(n6_c));
    defparam i1_2_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    uart_tx tx (.clk32MHz(clk32MHz), .n26810(n26810), .n26830(n26830), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .GND_net(GND_net), .r_SM_Main({r_SM_Main}), 
            .tx_o(tx_o), .tx_data({tx_data}), .\r_SM_Main_2__N_3336[0] (r_SM_Main_2__N_3336[0]), 
            .\r_SM_Main_2__N_3333[1] (\r_SM_Main_2__N_3333[1] ), .VCC_net(VCC_net), 
            .n14961(n14961), .n4(n4), .n14955(n14955), .tx_active(tx_active), 
            .n30923(n30923), .n7410(n7410), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n14794(n14794), .n14921(n14921), 
            .r_SM_Main({r_SM_Main_adj_11}), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
            .n14995(n14995), .rx_data({rx_data}), .\r_SM_Main_2__N_3262[2] (\r_SM_Main_2__N_3262[2] ), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_7 ), .n13657(n13657), 
            .GND_net(GND_net), .n4(n4_adj_8), .n4_adj_1(n4_adj_9), .n13652(n13652), 
            .n4_adj_2(n4_adj_10), .n25972(n25972), .n14971(n14971), .n14970(n14970), 
            .n14969(n14969), .n14968(n14968), .n14957(n14957), .n14964(n14964), 
            .n25630(n25630), .rx_data_ready(rx_data_ready), .VCC_net(VCC_net), 
            .n18503(n18503), .n14946(n14946), .n14945(n14945)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, n26810, n26830, \r_Bit_Index[0] , GND_net, 
            r_SM_Main, tx_o, tx_data, \r_SM_Main_2__N_3336[0] , \r_SM_Main_2__N_3333[1] , 
            VCC_net, n14961, n4, n14955, tx_active, n30923, n7410, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output n26810;
    output n26830;
    output \r_Bit_Index[0] ;
    input GND_net;
    output [2:0]r_SM_Main;
    output tx_o;
    input [7:0]tx_data;
    input \r_SM_Main_2__N_3336[0] ;
    output \r_SM_Main_2__N_3333[1] ;
    input VCC_net;
    input n14961;
    output n4;
    input n14955;
    output tx_active;
    input n30923;
    output n7410;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n4091;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n14873;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n18899, n3, n10918;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n8779, n8778, n30505, n30397, o_Tx_Serial_N_3364, n10, 
        n28053, n3_adj_3580, n30502, n30394, n22439, n22438, n22437, 
        n22436, n22435, n22434, n22433, n22432;
    
    SB_DFFESR r_Clock_Count_1132__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n4091), .D(n41[3]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1132__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n4091), .D(n41[2]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1132__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n4091), .D(n41[1]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n26810), 
            .D(n307[2]), .R(n26830));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n26810), 
            .D(n307[1]), .R(n26830));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1132__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n4091), .D(n41[0]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1215_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1215_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n18899));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i25135_3_lut (.I0(n26810), .I1(n18899), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n26830));
    defparam i25135_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1222_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1222_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n4091), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n8779), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1132__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n4091), .D(n41[4]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i5021_4_lut (.I0(\r_SM_Main_2__N_3336[0] ), .I1(n18899), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3333[1] ), .O(n8778));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5021_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i5022_3_lut (.I0(n8778), .I1(\r_SM_Main_2__N_3333[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n8779));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5022_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1540765_i1_3_lut (.I0(n30505), .I1(n30397), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3364));
    defparam i1540765_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3364), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[3]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[4]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n28053));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6956_2_lut_3_lut (.I0(\r_SM_Main_2__N_3333[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3580));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6956_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i3_4_lut (.I0(n28053), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3333[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25064_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3333[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n14873));
    defparam i25064_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1059_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n4091));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1059_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n30502));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n30502_bdd_4_lut (.I0(n30502), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n30505));
    defparam n30502_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_25371 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n30394));
    defparam r_Bit_Index_0__bdd_4_lut_25371.LUT_INIT = 16'he4aa;
    SB_LUT4 n30394_bdd_4_lut (.I0(n30394), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n30397));
    defparam n30394_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_1132__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n4091), .D(n41[8]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1132__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n4091), .D(n41[7]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1132__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n4091), .D(n41[6]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1132__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n4091), .D(n41[5]), .R(n14873));   // verilog/uart_tx.v(118[34:51])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n10918), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3580), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1132_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n22439), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1132_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22438), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_9 (.CI(n22438), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n22439));
    SB_LUT4 r_Clock_Count_1132_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22437), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_8 (.CI(n22437), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22438));
    SB_LUT4 r_Clock_Count_1132_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22436), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_7 (.CI(n22436), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22437));
    SB_LUT4 r_Clock_Count_1132_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22435), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_6 (.CI(n22435), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22436));
    SB_LUT4 r_Clock_Count_1132_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22434), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_5 (.CI(n22434), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22435));
    SB_LUT4 r_Clock_Count_1132_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22433), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_4 (.CI(n22433), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22434));
    SB_LUT4 r_Clock_Count_1132_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22432), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_3 (.CI(n22432), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22433));
    SB_LUT4 r_Clock_Count_1132_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1132_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1132_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22432));
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n14961));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3333[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3336[0] ), 
            .I3(r_SM_Main[1]), .O(n10918));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i25144_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3333[1] ), .O(n26810));
    defparam i25144_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n14955));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n30923));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3663_2_lut (.I0(\r_SM_Main_2__N_3336[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n7410));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i3663_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n14794, n14921, r_SM_Main, r_Rx_Data, RX_N_2, 
            n14995, rx_data, \r_SM_Main_2__N_3262[2] , \r_Bit_Index[0] , 
            n13657, GND_net, n4, n4_adj_1, n13652, n4_adj_2, n25972, 
            n14971, n14970, n14969, n14968, n14957, n14964, n25630, 
            rx_data_ready, VCC_net, n18503, n14946, n14945) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output n14794;
    output n14921;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input RX_N_2;
    input n14995;
    output [7:0]rx_data;
    output \r_SM_Main_2__N_3262[2] ;
    output \r_Bit_Index[0] ;
    output n13657;
    input GND_net;
    output n4;
    output n4_adj_1;
    output n13652;
    output n4_adj_2;
    input n25972;
    input n14971;
    input n14970;
    input n14969;
    input n14968;
    input n14957;
    input n14964;
    input n25630;
    output rx_data_ready;
    input VCC_net;
    output n18503;
    input n14946;
    input n14945;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    
    wire n14758;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n14871;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n30559, r_Rx_Data_R, n13484, n26006, n10, n28381;
    wire [2:0]r_SM_Main_2__N_3268;
    
    wire n26790, n6, n18742, n29307, n19057, n22431, n22430, n22429, 
        n22428, n22427, n22426, n22425, n29310, n30556;
    
    SB_DFFESR r_Clock_Count_1130__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n14758), .D(n37[7]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n14758), .D(n37[6]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n14758), .D(n37[5]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n14758), .D(n37[4]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n14758), .D(n37[3]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n14758), .D(n37[2]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1130__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n14758), .D(n37[1]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n14794), 
            .D(n326[2]), .R(n14921));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n14794), 
            .D(n326[1]), .R(n14921));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n30559), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1130__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n14758), .D(n37[0]), .R(n14871));   // verilog/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n14995));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(\r_SM_Main_2__N_3262[2] ), .O(n13484));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(n13484), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n13657));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_95_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_95_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_832 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n26006));
    defparam i1_2_lut_adj_832.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut (.I0(r_Clock_Count[3]), .I1(n26006), .I2(n10), .I3(r_Clock_Count[4]), 
            .O(\r_SM_Main_2__N_3262[2] ));
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i23291_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[4]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[0]), .O(n28381));
    defparam i23291_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut_adj_833 (.I0(r_Clock_Count[2]), .I1(n26006), .I2(n28381), 
            .I3(r_Clock_Count[5]), .O(r_SM_Main_2__N_3268[0]));
    defparam i3_4_lut_adj_833.LUT_INIT = 16'hffdf;
    SB_LUT4 i21711_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3268[0]), 
            .I3(GND_net), .O(n26790));
    defparam i21711_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_834 (.I0(r_SM_Main[2]), .I1(n26790), .I2(\r_SM_Main_2__N_3262[2] ), 
            .I3(r_SM_Main[1]), .O(n14871));
    defparam i1_4_lut_adj_834.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3268[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i25055_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n14758));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i25055_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i1193_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1193_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n18742));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_91_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_91_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_835 (.I0(\r_Bit_Index[0] ), .I1(n13484), .I2(GND_net), 
            .I3(GND_net), .O(n13652));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_835.LUT_INIT = 16'heeee;
    SB_LUT4 equal_94_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_94_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i11090_3_lut (.I0(n14794), .I1(n18742), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n14921));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i11090_3_lut.LUT_INIT = 16'h8a8a;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3262[2] ), 
            .R(n25972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3262[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n14794));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i24498_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3268[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n29307));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i24498_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n29307), .I1(\r_SM_Main_2__N_3262[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n19057));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n19057), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1200_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1200_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n14971));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n14970));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n14969));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n14968));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n14957));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1130_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n22431), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1130_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n22430), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n14964));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n25630));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1130_add_4_8 (.CI(n22430), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n22431));
    SB_LUT4 r_Clock_Count_1130_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n22429), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_7 (.CI(n22429), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n22430));
    SB_LUT4 r_Clock_Count_1130_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n22428), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_6 (.CI(n22428), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n22429));
    SB_LUT4 r_Clock_Count_1130_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n22427), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_5 (.CI(n22427), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n22428));
    SB_LUT4 r_Clock_Count_1130_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n22426), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_4 (.CI(n22426), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n22427));
    SB_LUT4 r_Clock_Count_1130_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n22425), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_3 (.CI(n22425), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n22426));
    SB_LUT4 r_Clock_Count_1130_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1130_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1130_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n22425));
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(\r_SM_Main_2__N_3262[2] ), .I1(r_SM_Main[1]), 
            .I2(n29310), .I3(r_SM_Main[0]), .O(n30556));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 n30556_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(r_SM_Main_2__N_3268[0]), 
            .I3(n30556), .O(n30559));   // verilog/uart_rx.v(70[21:38])
    defparam n30556_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i24511_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(\r_SM_Main_2__N_3262[2] ), .O(n29310));
    defparam i24511_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i14681_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n18503));
    defparam i14681_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n14946));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n14945));   // verilog/uart_rx.v(49[10] 144[8])
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n30021, VCC_net, INHA_c, clk32MHz, n13483, pwm_counter, 
            GND_net, n13481) /* synthesis syn_module_defined=1 */ ;
    input n30021;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n13483;
    output [31:0]pwm_counter;
    input GND_net;
    input n13481;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n27607, n8, n7, n27418, n28070, n10, pwm_counter_31__N_531;
    wire [31:0]n133;
    
    wire n22394, n22393, n22392, n22391, n22390, n22389, n22388, 
        n22387, n22386, n22385, n22384, n22383, n22382, n22381, 
        n22380, n22379, n22378, n22377, n22376, n22375, n22374, 
        n22373, n22372, n22371, n22370, n22369, n22368, n22367, 
        n22366, n22365, n22364;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n30021), 
            .R(n13483));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n27607));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(n27607), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n8));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut (.I0(pwm_counter[21]), .I1(pwm_counter[12]), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[22]), .I2(pwm_counter[19]), 
            .I3(pwm_counter[18]), .O(n27418));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[11]), .I1(n7), .I2(pwm_counter[20]), 
            .I3(n8), .O(n28070));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n28070), .I1(n13481), .I2(n27418), .I3(pwm_counter[15]), 
            .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14663_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[31]), .I2(n10), 
            .I3(pwm_counter[14]), .O(pwm_counter_31__N_531));   // verilog/pwm.v(18[8:40])
    defparam i14663_4_lut.LUT_INIT = 16'h3332;
    SB_DFFSR pwm_counter_1127__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1127_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n22394), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1127_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n22393), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_32 (.CI(n22393), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n22394));
    SB_LUT4 pwm_counter_1127_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n22392), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_31 (.CI(n22392), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n22393));
    SB_LUT4 pwm_counter_1127_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n22391), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_counter_1127__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_1127_add_4_30 (.CI(n22391), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n22392));
    SB_LUT4 pwm_counter_1127_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n22390), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_counter_1127__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1127__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_531));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_1127_add_4_29 (.CI(n22390), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n22391));
    SB_LUT4 pwm_counter_1127_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n22389), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_28 (.CI(n22389), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n22390));
    SB_LUT4 pwm_counter_1127_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n22388), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_27 (.CI(n22388), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n22389));
    SB_LUT4 pwm_counter_1127_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n22387), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_26 (.CI(n22387), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n22388));
    SB_LUT4 pwm_counter_1127_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n22386), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_25 (.CI(n22386), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n22387));
    SB_LUT4 pwm_counter_1127_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n22385), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_24 (.CI(n22385), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n22386));
    SB_LUT4 pwm_counter_1127_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n22384), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_23 (.CI(n22384), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n22385));
    SB_LUT4 pwm_counter_1127_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n22383), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_22 (.CI(n22383), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n22384));
    SB_LUT4 pwm_counter_1127_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n22382), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_21 (.CI(n22382), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n22383));
    SB_LUT4 pwm_counter_1127_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n22381), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_20 (.CI(n22381), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n22382));
    SB_LUT4 pwm_counter_1127_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n22380), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_19 (.CI(n22380), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n22381));
    SB_LUT4 pwm_counter_1127_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n22379), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_18 (.CI(n22379), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n22380));
    SB_LUT4 pwm_counter_1127_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n22378), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_17 (.CI(n22378), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n22379));
    SB_LUT4 pwm_counter_1127_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n22377), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_16 (.CI(n22377), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n22378));
    SB_LUT4 pwm_counter_1127_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n22376), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_15 (.CI(n22376), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n22377));
    SB_LUT4 pwm_counter_1127_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n22375), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_14 (.CI(n22375), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n22376));
    SB_LUT4 pwm_counter_1127_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n22374), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_13 (.CI(n22374), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n22375));
    SB_LUT4 pwm_counter_1127_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n22373), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_12 (.CI(n22373), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n22374));
    SB_LUT4 pwm_counter_1127_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n22372), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_11 (.CI(n22372), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n22373));
    SB_LUT4 pwm_counter_1127_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n22371), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_10 (.CI(n22371), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n22372));
    SB_LUT4 pwm_counter_1127_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n22370), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_9 (.CI(n22370), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n22371));
    SB_LUT4 pwm_counter_1127_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n22369), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_8 (.CI(n22369), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n22370));
    SB_LUT4 pwm_counter_1127_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n22368), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_7 (.CI(n22368), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n22369));
    SB_LUT4 pwm_counter_1127_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n22367), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_6 (.CI(n22367), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n22368));
    SB_LUT4 pwm_counter_1127_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n22366), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_5 (.CI(n22366), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n22367));
    SB_LUT4 pwm_counter_1127_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n22365), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_4 (.CI(n22365), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n22366));
    SB_LUT4 pwm_counter_1127_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n22364), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_3 (.CI(n22364), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n22365));
    SB_LUT4 pwm_counter_1127_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1127_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1127_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n22364));
    
endmodule
