// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Oct 23 21:04:31 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    input PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_0, PIN_7_c_1, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(42[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(43[12:17])
    
    wire n7, n27859, n27858;
    wire [7:0]blue;   // verilog/TinyFPGA_B.v(44[11:15])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(110[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(111[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(148[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(149[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(150[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(151[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(152[22:24])
    
    wire n27771, n17748, n27770, n27769;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(155[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(156[22:30])
    
    wire n27768, n27857, n27767, n27570, n27856;
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(159[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(183[22:33])
    
    wire n1225, n16532, n40881, color_23__N_34, n27766, n27765, 
        n27569;
    wire [22:0]pwm_setpoint_22__N_58;
    
    wire PIN_13_N_106;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_107;
    wire [24:0]displacement_23__N_205;
    wire [23:0]displacement_23__N_81;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n39563, start;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n28, n15;
    wire [3:0]state_3__N_337;
    
    wire n18367, n18371, n18370, n27855, n40100, n40098, n39559, 
        n18369, n18368, n11518, n11517, n11516, n32680, n27568, 
        n18366, n40092, n2, n32684, n2755, n27854, n27764, n27763, 
        n10705, n1220, n1219, n18365, n2754, n2753, n2682, n2683, 
        n2752, n28574, n28573, n28572, n28571, n28570, n28569, 
        n28568, n28567, n28566, n2751, n2750, n28565, n28564, 
        n2685, n2684, n28563, n28562, n28561, n28560, n28559, 
        n2749, n27853, n2748, n2747, n2746, n2745, n2744, n2743, 
        n2742, n2741, n2740, n2739, n2738, n2737, n28558, n2736, 
        n2735, n2734, n2733, n2732, n2705, n2704, n2703, n2702, 
        n2701, n2700, n28557, n4, n2699, n2698, n2697, n28556, 
        n34680, n28555, n2696, n27852, n27762, n28554, n28553, 
        n28552, n28551, n28550, n32692, n27851, n393, n392, n391, 
        n390, n389, n388, n387, n386, n385, n384, n383, n382, 
        n381, n380, n379, n378, n377, n376, n375, n374, n373, 
        n372, n371, n370, n369, n1155, n1154, n1153, n1152, 
        n1151, n28549, n2695, n28548, n28547, n28546, n28545, 
        n28544, n28543;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n28542;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n27850, n28541, n28540, n28539, n28538, n28537, n28536, 
        n28535, n28534, n28533, n28532, n28531, n28530, n28529, 
        n28528, n28527, n28526, n28525, n28524, n2694, n2693, 
        n2692, n27761, n27849, n28523, n28522, n28521, n28520, 
        n28519, n28518, n28517, n28516, n28515, n28514, n28513, 
        n28512, n28511, n28510, n3, n4_adj_3930, n5, n6, n7_adj_3931, 
        n8, n9, n10, n11, n12, n13, n14, n15_adj_3932, n16, 
        n17, n18, n19, n20, n21, n22, n23, n24, n25, n28509, 
        n28508, n28507, n28506, n28505, n28504, n28503, n28502, 
        n28501, n28500, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n27848, n39549;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n16523, n16520, n16517, n16508, n16505, n16502, n16498;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n1125, n1124, n1123, n1122, n1121, n1120, n123, n40052, 
        n28499, n27847, n27846, n27845, n37, n27844, n27843, n27760, 
        n35, n9783, n27759, n34, n32, n31, n27758, n27842, n25_adj_3933, 
        n28498, n28497, n27757, n28496, n28495, n28494, n28493, 
        n40487, n28492, n28491, n28490, n28489, n40463, n40003, 
        n28488, n27841, n27840, n27839, n40001, n27838, n27837, 
        n28487, n28486, n28485, n28484, n28483, n6_adj_3934, n28482, 
        n25598, n28481, n28480, n28479, n28478, n34667, n6_adj_3935, 
        n28477, n28476, n4_adj_3936, n27836, n39993, n28475, n28474, 
        n39991, n40878, n39981, n39537, n34769, n39979, n39975, 
        n16495, n16544, n39973, n16491, n16541, n39969, n2_adj_3937, 
        n39967, n27835, n40488, n39527, n27834, n24632, n28473, 
        n28472, n28471, n28470, n16485, n16538, n39523, n39955, 
        n39953, n39951, n40515, n16475, n47, n46, n16535, n39948, 
        n43, n39946, n42, n40, n39, n28469, n38, n27833, n29221, 
        n16809, n16472, n28468, n28467, n28466, n28465, n28464, 
        n28463, n28462, n28461, n28460, n31_adj_3938, n28459, n28458, 
        n29220, n2691, n2690, n2346, n28457, n29219, n28456, n2689, 
        n28455, n28454, n28453, n28452, n28451, n28450, n2857, 
        n39519, n44, n43_adj_3939, n28449, n28448, n28447, n28446, 
        n29218, n34624, n34730, n42_adj_3940, n41, n40_adj_3941, 
        n38_adj_3942, n28445, n28444, n29217, n15_adj_3943, n27832, 
        n28443, n29216, n29215, n3761, n39904, n30, n29214, n29213, 
        n26, n16_adj_3944, n11_adj_3945, n10_adj_3946, n21_adj_3947, 
        n155, n131, n175, n29212, n39808, n40482, n29211, n29210, 
        n29209, n42_adj_3948, n41_adj_3949, n40_adj_3950, n39_adj_3951, 
        n37_adj_3952, n29208, n36, n29207, n40480, n29, n39507, 
        n27831, n39501, n27830, n27829, n27828, n27827, n27826, 
        n27825, n27824, n27823, n27822, n27821, n39499, n27820, 
        n27819, n16424, n27818, n27817, n39495, n39491, n40467, 
        n28442, n28441, n28440, n28439, n28438, n28437, n28436, 
        n28435, n28434, n28433, n28432, n29206, n2_adj_3953, n28431, 
        n28430, n28429, n28428, n28427, n28426, n28425, n28424, 
        n28423, n28422, n28421, n28420, n28419, n28418, n28417, 
        n28416, n28415, n28414, n28413, n28412, n28411, n28410, 
        n28409, n28408, n28407, n28406, n28405, n28404, n28403, 
        n29205, n28402, n28401, n29204, n29203, n28400, n28399, 
        n28398, n28397, n4684, n28396, n18245, n18244, n18243, 
        n18242, n18241, n18240, n18239, n29202, n18238, n18237, 
        n18236, n18235, n18234, n18233, n18232, n18231, n18230, 
        n18229, n18228, n18227, n18226, n18225, n18224, n18223, 
        n18222, n18221, n18220, n18219, n18218, n18217, n18216, 
        n18215, n18214, n18213, n18212, n18211, n18210, n18209, 
        n18208, n18207, n18206, n18205, n18204, n18203, n18202, 
        n18201, n18200, n18199, n18198, n18197, n18196, n18195, 
        n18194, n18193, n18192, n18191, n18190, n18189, n18188, 
        n18187, n18186, n18185, n18184, n18183, n18182, n18181, 
        n18180, n18179, n18178, n18177, n18176, n18175, n18174, 
        n18173, n18172, n18171, n18170, n18169, n18168, n18167, 
        n18166, n18165, n18164, n18163, n18162, n18161, n18160, 
        n18159, n18158, n18157, n18156, n18155, n18154, n18153, 
        n18152, n18151, n18150, n18149, n18148, n18147, n18146, 
        n18145, n18144, n18143, n18142, n18141, n18140, n18139, 
        n18138, n18137, n18136, n18135, n18134, n18133, n18132, 
        n18131, n18130, n18129, n18128, n18127, n18126, n18125, 
        n18124, n18123, n18122, n18121, n18120, n18119, n18118, 
        n18114, n18113, n18112, n18111, n18110, n18109, n18108, 
        n18107, n18106, n18105, n18104, n18103, n18102, n18101, 
        n18100, n18099, n18098, n18097, n18096, n18095, n18094, 
        n18093, n18092, n18091, n18090, n18089, n18088, n18087, 
        n18086, n18085, n18084, n18083, n18082, n18081, n18080, 
        n18079, n18078, n18077, n18075, n18074, n18073, n18072, 
        n18071, n18070, n18069, n18068, n18067, n18066, n18065, 
        n18064, n18063, n18062, n18061, n18060, n18059, n18058, 
        n18057, n18056, n18055, n18054, n18053, n18052, n18051, 
        n18050, n18049, n18048, n18047, n18046, n18045, n18044, 
        n18043, n18042, n18041, n18040, n18039, n18038, n18037, 
        n18036, n18035, n18034, n18033, n18032, n18031, n32742, 
        n39485, n29201, n249, n248, n39479, n224, n1085, n29200, 
        n39475, n1184, n29199, n39896, n29198, n1058, n1057, n1056, 
        n18030, n18029, n11515, n1055, n1054, n1053, n1052, n18028, 
        n99, n98, n97, n96, n95, n94, n93, n92, n91, n90, 
        n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, 
        n79, n18027, n18026, n18025, n18024, n18023, n78, n77, 
        n75, n74, n73, n72, n71, n70, n69, n68, n67, n66, 
        n65, n64, n63, n62, n61, n60, n59, n58, n57, n56, 
        n55, n54, n39467, n2688, n2687, n2686, n40471, n1035, 
        n53, n1250, n1251, n1252, n16514, n28395, n4706, n29197, 
        n28394, n16429, n39460, n33766, n40479, n33, n32_adj_3954, 
        n31_adj_3955, n30_adj_3956, n29_adj_3957, n28_adj_3958, n27, 
        n26_adj_3959, n25_adj_3960, n24_adj_3961, n23_adj_3962, n22_adj_3963, 
        n21_adj_3964, n20_adj_3965, n19_adj_3966, n18_adj_3967, n17_adj_3968, 
        n16_adj_3969, n15_adj_3970, n14_adj_3971, n13_adj_3972, n12_adj_3973, 
        n11_adj_3974, n10_adj_3975, n9_adj_3976, n8_adj_3977, n7_adj_3978, 
        n6_adj_3979, n5_adj_3980, n4_adj_3981, n3_adj_3982, n13950, 
        n28393, n2_adj_3983, n32694, n28392, n29196, n28391, n28390, 
        n28389, n28388, n28387, n29195, n27816, n29194, n27815, 
        n40850, n29193, n29192, n29191, n28386, n4446, n4445, 
        n4444, n4443, n4442, n4441, n4440, n4439, n4438, n4437, 
        n4436, n4435, n4434, n4433, n4432, n4431, n4430, n4429, 
        n4428, n4427, n4426, n4425, n4424, n4423, n29190, n27814, 
        n27813, n29189, n27589, n34749, n27812, n28385, n27811, 
        n28384, n27588, n28383, quadA_debounced, quadB_debounced, 
        count_enable, n28382, n3_adj_3984, n28381, n28380, n28379, 
        n28378, n27810, n15_adj_3985, n28377, n25_adj_3986, n24_adj_3987, 
        n23_adj_3988, n22_adj_3989, n21_adj_3990, n20_adj_3991, n19_adj_3992, 
        n18_adj_3993, n17_adj_3994, n16_adj_3995, n15_adj_3996, n14_adj_3997, 
        n13_adj_3998, n12_adj_3999, n11_adj_4000, n10_adj_4001, n9_adj_4002, 
        n8_adj_4003, n7_adj_4004, n6_adj_4005, n5_adj_4006, n4_adj_4007, 
        n28376, n6_adj_4008, n28375, n28374, n28373, n28372, n28371, 
        quadA_debounced_adj_4009, quadB_debounced_adj_4010, count_enable_adj_4011, 
        n39455, n28370, n28369, n28368, n28367, n28366, n28365, 
        n28364, n28363, n28362, n28361, n28360, n28359, n28358, 
        n28357, n28356, n3_adj_4012, n8_adj_4013, n28355, n28354, 
        n29188, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n29187, n29186, n27809, n220, n222, n224_adj_4014, n225, 
        n226, n16417, n32696;
    wire [2:0]r_SM_Main_adj_4662;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_4664;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3298;
    wire [2:0]r_SM_Main_2__N_3295;
    
    wire n39657, n18003, n18000;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    wire [1:0]reg_B_adj_4672;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n6666, n39653, n6665, n6664, n6663, n6662, n6661, n4_adj_4022, 
        n6673, n6672, n6671, n4_adj_4023, n28312, n28311, n6670, 
        n6669, n28310, n28309, n28308, n28307, n28306, n28305, 
        n28304, n28303, n27808, n28302, n28301, n28300, n40470, 
        n28299, n28298, n28297, n28296, n28295, n28294, n28293, 
        n39440, n28292, n28291, n28290, n28289, n28288, n28287, 
        n28286, n28285, n28284, n28283, n28282, n10710, n39436, 
        n28281, n39434, n10709, n10708, n10707, n28280, n10706, 
        n1258, n1257, n28279, n1256, n1255, n28278, n1254, n1253, 
        n28277, n28276, n28275, n8_adj_4024, n9_adj_4025, n10_adj_4026, 
        n11_adj_4027, n12_adj_4028, n13_adj_4029, n14_adj_4030, n15_adj_4031, 
        n16_adj_4032, n17_adj_4033, n18_adj_4034, n19_adj_4035, n20_adj_4036, 
        n21_adj_4037, n22_adj_4038, n23_adj_4039, n24_adj_4040, n25_adj_4041, 
        n16421, n28274, n1025, n1024, n1023, n1022, n1021, n41916, 
        n40469, n27807, n39432, n40492, n986, n28273, n510, n533, 
        n534, n558, n40304, n40973, n958, n957, n956, n955, 
        n954, n953, n13_adj_4042, n648, n649, n28272, n11_adj_4043, 
        n671, n672, n27806, n28271, n17721, n39418, n783, n784, 
        n785, n27805, n806, n807, n27804, n38_adj_4044, n37_adj_4045, 
        n36_adj_4046, n6708, n35_adj_4047, n914, n915, n916, n917, 
        n918, n938, n939, n33_adj_4048, n855, n852, n6674, n6675, 
        n6685, n6696, n26_adj_4049, n1043, n1044, n1045, n1046, 
        n1047, n1048, n40334, n1067, n1068, n3477, n22_adj_4050, 
        n28_adj_4051, n32708, n6678, n6679, n6680, n6681, n6682, 
        n6683, n6684, n1169, n1170, n1171, n1172, n1173, n1174, 
        n1175, n3459, n3458, n3457, n3456, n3455, n3454, n3453, 
        n3452, n26_adj_4052, n1193, n1194, n24_adj_4053, n6688, 
        n6689, n6690, n6691, n6692, n6693, n6694, n6695, n19_adj_4054, 
        n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n39374, n7_adj_4055, n16_adj_4056, n1316, n1317, n16404, 
        n6718, n6717, n6716, n6715, n6714, n6713, n6712, n6711, 
        n749, n748, n746, n6699, n6700, n6701, n6702, n6703, 
        n6704, n6705, n6706, n6707, n6726, n6727, n6728, n6729, 
        n6730, n6731, n6732, n6733, n6734, n6735, n6750, n11748, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n6725, n3362, n28270, n3358, n3357, n3356, n3355, 
        n3354, n3353, n3351, n1436, n1437, n3346, n3344, n3343, 
        n3340, n3337, n39372, n6719, n6720, n6721, n3321, n3322, 
        n3323, n3324, n3325, n3330, n39370, n39368, n1529, n1530, 
        n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
        n3320, n3319, n3318, n3317, n3316, n3315, n3314, n3313, 
        n3312, n3311, n3310, n3309, n3308, n3307, n1553, n1554, 
        n39366, n3305, n3304, n3303, n3302, n3301, n3300, n3299, 
        n3298, n6765, n6758, n6759, n6760, n6761, n6762, n6763, 
        n6764, n28269, n1643, n1644, n1645, n1646, n1647, n1648, 
        n1649, n1650, n1651, n1652, n1653, n6757, n6756, n6755, 
        n6754, n6753, n6780, n6779, n6778, n6777, n6776, n6775, 
        n6774, n6773, n1667, n1668, n6771, n6770, n3263, n28268, 
        n3258, n3257, n3256, n3255, n3254, n28267, n6738, n6739, 
        n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, 
        n6748, n6749, n28266, n3243, n3244, n3245, n3246, n3247, 
        n3248, n3249, n3250, n3251, n3252, n3253, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n3242, n3241, n3240, n3239, n3238, n3237, 
        n3236, n3235, n3234, n3233, n3232, n3231, n1778, n1779, 
        n34_adj_4057, n33_adj_4058, n32_adj_4059, n31_adj_4060, n3225, 
        n3224, n3223, n3222, n3221, n3220, n3219, n30_adj_4061, 
        n6766, n3209, n3210, n3211, n3212, n3213, n3214, n3215, 
        n3216, n3217, n3218, n1862, n1863, n1864, n1865, n1866, 
        n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
        n3208, n3207, n3206, n3205, n3204, n3203, n3202, n3201, 
        n3200, n3199, n1886, n1887, n6804, n6834, n6781, n6782, 
        n6783, n6801, n6825, n6826, n6827, n6828, n6829, n6830, 
        n6831, n6832, n6833, n1967, n1968, n1969, n1970, n1971, 
        n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n6824, n6823, n6852, n6851, n6850, n6849, n6848, 
        n6847, n6846, n6845, n1991, n1992, n6843, n3164, n28265, 
        n3158, n3157, n6786, n6787, n6788, n6789, n6790, n6791, 
        n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, 
        n6800, n3149, n3150, n3151, n3152, n3153, n3154, n3155, 
        n3156, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
        n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
        n3148, n3147, n3146, n3145, n3144, n3143, n3142, n3141, 
        n3140, n2093, n2094, n3138, n3137, n3136, n3135, n3134, 
        n3133, n3132, n3131, n6806, n6807, n6808, n6809, n6810, 
        n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, 
        n6819, n6820, n3124, n3125, n40491, n2168, n2169, n2170, 
        n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
        n2179, n2180, n2181, n2182, n2183, n3123, n3122, n3121, 
        n3120, n3119, n3118, n3117, n3116, n2192, n2193, n28264, 
        n3114, n3113, n3112, n3111, n3110, n3109, n3108, n6835, 
        n6836, n6837, n6838, n6839, n6840, n3102, n3103, n3104, 
        n3105, n3106, n3107, n2264, n2265, n2266, n2267, n2268, 
        n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
        n2277, n2278, n2279, n2280, n3101, n3100, n2288, n2289, 
        n28263, n28262, n28261, n6853, n6854, n6855, n6856, n6857, 
        n6858, n6859, n6860, n6861, n6883, n6906, n6930, n6955, 
        n39342, n27587, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
        n2371, n2372, n2373, n2374, n2381, n2382, n6864, n6865, 
        n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
        n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
        n6882, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
        n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, 
        n2462, n2463, n2464, n2465, n3065, n28260, n2471, n2472, 
        n3058, n3057, n3056, n6886, n6887, n6888, n6889, n6890, 
        n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, 
        n6899, n6900, n6901, n6902, n6903, n6904, n6905, n3053, 
        n3054, n3055, n2534, n2535, n2536, n2537, n2538, n2539, 
        n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
        n2548, n2549, n2550, n2551, n2552, n2553, n3052, n3051, 
        n3050, n3049, n2558, n2559, n8_adj_4062, n3047, n3046, 
        n3045, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
        n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
        n6924, n6925, n6926, n6927, n6928, n6929, n3043, n3044, 
        n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
        n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
        n2634, n2635, n2636, n2637, n2638, n3042, n3041, n3040, 
        n2642, n2643, n7_adj_4063, n26_adj_4064, n3038, n3037, n6933, 
        n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
        n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
        n6950, n6951, n6952, n6953, n6954, n3036, n2699_adj_4065, 
        n2700_adj_4066, n2701_adj_4067, n2702_adj_4068, n2703_adj_4069, 
        n2704_adj_4070, n2705_adj_4071, n2706, n2707, n2708, n2709, 
        n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
        n2718, n2719, n2720, n3035, n3034, n2723, n2724, n39306, 
        n24_adj_4072, n22_adj_4073, n3033, n3032, n2777, n2798, 
        n2799, n2801, n2802, n18_adj_4074, n28259, n32698, n17992, 
        n17989, n32700, n17980, n17974, n17973, n17972, n17971, 
        n17970, n3025, n3024, n3023, n3022, n3021, n3020, n3019, 
        n3018, n3017, n3016, n3015, n3014, n3013, n3012, n3011, 
        n3010, n3009, n3008, n3007, n3006, n3005, n17969, n28258, 
        n28257, n3004, n28256, n28255, n3003, n3002, n28254, n28253, 
        n28252, n3001, n28251, n28250, n16529, n28249, n28248, 
        n28247, n28246, n12_adj_4075, n28245, n28244, n2966, n28243, 
        n28242, n28241, n28240, n28239, n2958, n2957, n39291, 
        n63_adj_4076, n2956, n2955, n2954, n2953, n2952, n2951, 
        n2950, n2949, n2948, n40028, n2947, n2946, n2945, n2944, 
        n2943, n2942, n2941, n2940, n2939, n2938, n2937, n2936, 
        n2935, n2934, n2933, n17968, n2925, n2924, n5_adj_4077, 
        n2923, n2922, n2921, n1224, n2920, n1223, n2919, n2918, 
        n2917, n2916, n2915, n2914, n39630, n2913, n2912, n2911, 
        n2910, n2909, n2908, n2907, n2906, n2905, n2904, n2903, 
        n2902, n28238, n39287, n28237, n18539, n28236, n28235, 
        n28234, n1222, n1221, n1158, n1157, n28233, n28232, n28231, 
        n28230, n28229, n28228, n28227, n28226, n32686, n2867, 
        n18518, n28225, n18517, n33775, n18515, n18514, n18513, 
        n18512, n28224, n18510, n2858, n18509, n2857_adj_4078, n2856, 
        n2855, n2854, n2853, n34715, n2852, n32682, n2851, n32690, 
        n2850, n2849, n2848, n2847, n2846, n2845, n2844, n2843, 
        n2842, n2841, n2840, n2839, n2838, n2837, n2836, n2835, 
        n2834, n32688, n2825, n2824, n2823, n2822, n18498, n18497, 
        n18496, n18495, n18494, n18493, n18492, n18491, n18490, 
        n18489, n18488, n18487, n18486, n18485, n18484, n18483, 
        n18482, n18481, n18480, n18479, n18478, n18477, n18476, 
        n18475, n34622, n18473, n18472, n2821, n2820, n2819, n2818, 
        n2817, n2816, n2815, n2814, n2813, n2812, n2811, n2810, 
        n2809, n2808, n2807, n2806, n2805, n2804, n2803, n18471, 
        n18470, n18469, n18468, n18467, n18466, n18465, n18464, 
        n18463, n18462, n18461, n18460, n18459, n18458, n18457, 
        n18456, n18455, n18454, n18453, n18452, n18451, n18450, 
        n18449, n18448, n18447, n18446, n18445, n18444, n18443, 
        n18442, n18441, n18440, n28223, n28222, n40535, n17967, 
        n17966, n17965, n17964, n17963, n17962, n17961, n17960, 
        n17959, n17958, n17957, n17956, n17955, n17954, n17953, 
        n17952, n17951, n17950, n17949, n28221, n17948, n17947, 
        n17946, n17945, n28220, n17943, n17942, n40501, n17936, 
        n28219, n17932, n17931, n28218, n32702, n28217, n17922, 
        n32710, n17911, n28216, n32712, n39283, n32714, n17900, 
        n17899, n17897, n28215, n17896, n17895, n17893, n17892, 
        n32722, n30686, n32724, n32726, n32728, n28214, n32730, 
        n32732, n32734, n32736, n32738, n28213, n32744, n39281, 
        n18439, n18438, n18437, n18436, n18435, n18434, n18433, 
        n18432, n18431, n18430, n18429, n18428, n18427, n18426, 
        n18425, n18424, n18423, n18422, n18421, n39277, n2768, 
        n28212, n2758, n2757, n2756, n2755_adj_4079, n2754_adj_4080, 
        n2753_adj_4081, n2752_adj_4082, n2751_adj_4083, n2750_adj_4084, 
        n2749_adj_4085, n2748_adj_4086, n2747_adj_4087, n2746_adj_4088, 
        n2745_adj_4089, n2744_adj_4090, n2743_adj_4091, n2742_adj_4092, 
        n2741_adj_4093, n2740_adj_4094, n2739_adj_4095, n2738_adj_4096, 
        n2737_adj_4097, n2736_adj_4098, n2735_adj_4099, n2725, n2724_adj_4100, 
        n2723_adj_4101, n2722, n2721, n2720_adj_4102, n18372, n2719_adj_4103, 
        n2718_adj_4104, n2717_adj_4105, n2716_adj_4106, n2715_adj_4107, 
        n2714_adj_4108, n2713_adj_4109, n2712_adj_4110, n2711_adj_4111, 
        n2710_adj_4112, n2709_adj_4113, n2708_adj_4114, n2707_adj_4115, 
        n17625, n2706_adj_4116, n2705_adj_4117, n2704_adj_4118, n17619, 
        n28211, n28210, n28209, n28208, n28207, n2669, n28206, 
        n2658, n2657, n2656, n2655, n2654, n2653, n2652, n2651, 
        n2650, n2649, n2648, n2647, n2646, n28205, n1580, n28_adj_4119, 
        n2643_adj_4120, n1646_adj_4121, n1615, n1647_adj_4122, n1616, 
        n1648_adj_4123, n1617, n1649_adj_4124, n1618, n1650_adj_4125, 
        n1619, n1651_adj_4126, n1620, n1652_adj_4127, n1621, n1653_adj_4128, 
        n1622, n1654, n1623, n1655, n1624, n1656, n1625, n1657, 
        n1658, n39265, n2644, n2645, n134, n135, n136, n137, 
        n138, n139, n140, n141, n142, n143, n144, n145, n146, 
        n147, n148, n149, n150, n151, n152, n153, n154, n155_adj_4129, 
        n156, n157, n158, n159, n160, n161, n162, n163, n164, 
        n165, n1547, n1548, n1549, n1550, n1551, n1552, n1553_adj_4130, 
        n1554_adj_4131, n1555, n1556, n1557, n1558, n27_adj_4132, 
        n26_adj_4133, n2642_adj_4134, n1516, n1517, n1518, n1519, 
        n1520, n1521, n1522, n1523, n1524, n1525, n25_adj_4135, 
        n2641, n2639, n2638_adj_4136, n2637_adj_4137, n2636_adj_4138, 
        n28204, n17746, n2625_adj_4139, n2624_adj_4140, n2623_adj_4141, 
        n2622_adj_4142, n17561, n2621_adj_4143, n2620_adj_4144, n2619_adj_4145, 
        n2618_adj_4146, n2617, n2616, n28203, n34698, n2615, n2614, 
        n34777, n2613, n2612, n28202, n2611, n2610, n2609, n2608, 
        n2607, n2606, n2605, n28201, n28200, n17843, n28199, n17842, 
        n2640, n38_adj_4147, n39_adj_4148, n40_adj_4149, n41_adj_4150, 
        n42_adj_4151, n43_adj_4152, n44_adj_4153, n45, n17841, n28198, 
        n1481, n40523, n1448, n1417_adj_4154, n1449, n1418_adj_4155, 
        n1450, n1419_adj_4156, n1451, n1420_adj_4157, n1452, n1421, 
        n1453, n1422, n1454, n1423, n1455, n1424, n1456, n1425, 
        n1457, n1458, n17840, n17536, n28197, n1353, n1354, n1355, 
        n1356, n1357, n1358, n28196, n28195, n28194, n1382, n2570, 
        n1322, n1323, n1324, n1325, n17839, n17522, n1349, n1350, 
        n1351, n1352, n28193, n1318, n1319, n1320, n1321, n32716, 
        n32718, n32720, n17793, n17792, n17838, n17837, n17836, 
        n17833, n17830, n17827, n1283, n2556, n28192, n2557, n2558_adj_4158, 
        n32746, n1156, n2555, n2554, n2553_adj_4159, n2552_adj_4160, 
        n2551_adj_4161, n2550_adj_4162, n2549_adj_4163, n2548_adj_4164, 
        n2547_adj_4165, n2546_adj_4166, n2545_adj_4167, n2544_adj_4168, 
        n2543_adj_4169, n2542_adj_4170, n2541_adj_4171, n2540_adj_4172, 
        n2539_adj_4173, n2538_adj_4174, n2537_adj_4175, n2525, n2524, 
        n2523, n2522, n2521, n2520, n2519, n2518, n2517, n2516, 
        n2515, n2514, n2513, n2512, n2511, n2510, n2509, n2508, 
        n2507, n2506, n32748, n39232, n39230, n2_adj_4176, n3_adj_4177, 
        n4_adj_4178, n5_adj_4179, n6_adj_4180, n7_adj_4181, n8_adj_4182, 
        n9_adj_4183, n10_adj_4184, n11_adj_4185, n12_adj_4186, n13_adj_4187, 
        n14_adj_4188, n15_adj_4189, n16_adj_4190, n17_adj_4191, n18_adj_4192, 
        n19_adj_4193, n20_adj_4194, n21_adj_4195, n22_adj_4196, n23_adj_4197, 
        n24_adj_4198, n25_adj_4199, n2_adj_4200, n3_adj_4201, n4_adj_4202, 
        n5_adj_4203, n6_adj_4204, n7_adj_4205, n8_adj_4206, n9_adj_4207, 
        n10_adj_4208, n11_adj_4209, n12_adj_4210, n13_adj_4211, n14_adj_4212, 
        n15_adj_4213, n16_adj_4214, n17_adj_4215, n18_adj_4216, n19_adj_4217, 
        n20_adj_4218, n21_adj_4219, n22_adj_4220, n23_adj_4221, n24_adj_4222, 
        n25_adj_4223, n2471_adj_4224, n28191, n2458_adj_4225, n2457_adj_4226, 
        n2456_adj_4227, n2455_adj_4228, n2454_adj_4229, n2453_adj_4230, 
        n2452_adj_4231, n2451_adj_4232, n2450_adj_4233, n2449_adj_4234, 
        n2448_adj_4235, n2447_adj_4236, n2446, n2445, n2444, n2443, 
        n2442, n2441, n2440, n2439, n2438, n28190, n28189, n28188, 
        n2425, n2424, n28187, n2423, n2422, n2421, n2420, n2419, 
        n2418, n2417, n2416, n2415, n2414, n2413, n2412, n2411, 
        n2410, n2409, n2408, n2407, n28186, n28185, n2372_adj_4237, 
        n28184, n28183, n39226, n28182, n40874, n2358_adj_4238, 
        n2357_adj_4239, n2356, n2355, n2354, n2353, n2352, n2351, 
        n2350, n2349, n2348, n2347, n2346_adj_4240, n2345, n2344, 
        n2343, n2342, n2341, n2340, n2339, n2325, n2324, n2323, 
        n2322, n2321, n2320, n2319, n2318, n2317, n2316, n2315, 
        n2314, n2313, n2312, n2311, n2310, n2309, n2308, n46_adj_4241, 
        n39220, n28181, n28180, n28179, n28178, n2273_adj_4242, 
        n28177, n2258, n2257, n2256, n2255, n2254, n2253, n2252, 
        n2251, n2250, n2249, n2248, n2247, n28176, n44_adj_4243, 
        n40555, n2246, n28175, n2245, n2244, n2243, n2242, n2241, 
        n2240, n2225, n2224, n2223, n2222, n2221, n2220, n2219, 
        n2218, n2217, n2216, n2215, n2214, n2213, n2212, n2211, 
        n2210, n2209, n28174, n42_adj_4244, n2174_adj_4245, n28173, 
        n2158, n2157, n2156, n2155, n2154, n2153, n2152, n2151, 
        n2150, n2149, n2148, n2147, n2146, n2145, n2144, n2143, 
        n2142, n2141, n28172, n28171, n28170, n40_adj_4246, n42_adj_4247, 
        n44_adj_4248, n45_adj_4249, n28169, n28168, n28167, n2125, 
        n2124, n2123, n2122, n2121, n2120, n2119, n2118, n2117, 
        n2116, n2115, n2114, n2113, n2112, n2111, n2110, n39216, 
        n38_adj_4250, n40_adj_4251, n42_adj_4252, n43_adj_4253, n40561, 
        n40818, n2075_adj_4254, n28166, n27803, n40856, n2058, n2057, 
        n2056, n2055, n2054, n2053, n2052, n2051, n2050, n2049, 
        n2048, n2047, n2046, n2045, n2044, n2043, n2042, n28165, 
        n36_adj_4255, n38_adj_4256, n40_adj_4257, n41_adj_4258, n39212, 
        n2025, n2024, n2023, n2022, n2021, n2020, n2019, n2018, 
        n2017, n2016, n2015, n2014, n2013, n2012, n2011, n28164, 
        n34_adj_4259, n36_adj_4260, n38_adj_4261, n39_adj_4262, n41_adj_4263, 
        n43_adj_4264, n40517, n45_adj_4265, n40563, n1976_adj_4266, 
        n28163, n28162, n28161, n1958, n1957, n1956, n1955, n1954, 
        n1953, n1952, n1951, n1950, n1949, n1948, n1947, n28160, 
        n32_adj_4267, n34_adj_4268, n37_adj_4269, n39_adj_4270, n41_adj_4271, 
        n40826, n43_adj_4272, n1946, n1945, n1944, n1943, n40967, 
        n1925, n1924, n1923, n1922, n1921, n1920, n1919, n1918, 
        n1917, n1916, n1915, n1914, n1913, n1912, n28159, n30_adj_4273, 
        n31_adj_4274, n32_adj_4275, n33_adj_4276, n34_adj_4277, n35_adj_4278, 
        n37_adj_4279, n39_adj_4280, n41_adj_4281, n42_adj_4282, n43_adj_4283, 
        n45_adj_4284, n40858, n3306, n28158, n1877, n28157, n28156, 
        n28_adj_4285, n29_adj_4286, n30_adj_4287, n31_adj_4288, n32_adj_4289, 
        n33_adj_4290, n35_adj_4291, n37_adj_4292, n40507, n39_adj_4293, 
        n40_adj_4294, n41_adj_4295, n43_adj_4296, n40816, n6772, n1858, 
        n1857, n1856, n1855, n1854, n1853, n1852, n1851, n1850, 
        n1849, n1848, n1847, n1846, n1845, n1844, n28155, n26_adj_4297, 
        n27_adj_4298, n28_adj_4299, n29_adj_4300, n30_adj_4301, n31_adj_4302, 
        n33_adj_4303, n35_adj_4304, n37_adj_4305, n38_adj_4306, n39_adj_4307, 
        n41_adj_4308, n40935, n3230, n28154, n24_adj_4309, n25_adj_4310, 
        n26_adj_4311, n27_adj_4312, n28_adj_4313, n29_adj_4314, n30_adj_4315, 
        n31_adj_4316, n32_adj_4317, n33_adj_4318, n35_adj_4319, n36_adj_4320, 
        n37_adj_4321, n39_adj_4322, n41_adj_4323, n43_adj_4324, n44_adj_4325, 
        n45_adj_4326, n40336, n39669, n6805, n22_adj_4327, n23_adj_4328, 
        n24_adj_4329, n25_adj_4330, n26_adj_4331, n27_adj_4332, n28_adj_4333, 
        n29_adj_4334, n30_adj_4335, n31_adj_4336, n33_adj_4337, n34_adj_4338, 
        n35_adj_4339, n37_adj_4340, n39_adj_4341, n41_adj_4342, n42_adj_4343, 
        n43_adj_4344, n40340, n40882, n40682, n1778_adj_4345, n28153, 
        n28152, n34782, n28151, n6844, n34645, n28150, n1758_adj_4346, 
        n1757_adj_4347, n1756_adj_4348, n28149, n20_adj_4349, n21_adj_4350, 
        n22_adj_4351, n23_adj_4352, n24_adj_4353, n25_adj_4354, n26_adj_4355, 
        n27_adj_4356, n28_adj_4357, n29_adj_4358, n31_adj_4359, n32_adj_4360, 
        n33_adj_4361, n35_adj_4362, n37_adj_4363, n39_adj_4364, n41_adj_4365, 
        n40877, n1755_adj_4366, n1754_adj_4367, n1753, n39189, n1752, 
        n1751, n1750, n1749, n1748, n3139, n1747, n1746, n1745, 
        n28148, n18_adj_4368, n19_adj_4369, n20_adj_4370, n21_adj_4371, 
        n22_adj_4372, n23_adj_4373, n24_adj_4374, n25_adj_4375, n26_adj_4376, 
        n27_adj_4377, n29_adj_4378, n30_adj_4379, n31_adj_4380, n33_adj_4381, 
        n35_adj_4382, n37_adj_4383, n39_adj_4384, n41_adj_4385, n42_adj_4386, 
        n43_adj_4387, n45_adj_4388, n40342, n39187, n3115, n1725, 
        n1724, n1723, n1722, n1721, n1720, n1719, n1718, n1717, 
        n28147, n16_adj_4389, n17_adj_4390, n18_adj_4391, n19_adj_4392, 
        n20_adj_4393, n21_adj_4394, n22_adj_4395, n23_adj_4396, n25_adj_4397, 
        n27_adj_4398, n28_adj_4399, n29_adj_4400, n31_adj_4401, n33_adj_4402, 
        n35_adj_4403, n40883, n37_adj_4404, n39_adj_4405, n40589, 
        n41_adj_4406, n43_adj_4407, n1716, n1715, n1714, n14_adj_4408, 
        n16_adj_4409, n17_adj_4410, n18_adj_4411, n19_adj_4412, n20_adj_4413, 
        n21_adj_4414, n22_adj_4415, n23_adj_4416, n25_adj_4417, n26_adj_4418, 
        n27_adj_4419, n29_adj_4420, n31_adj_4421, n33_adj_4422, n35_adj_4423, 
        n37_adj_4424, n39_adj_4425, n40_adj_4426, n41_adj_4427, n43_adj_4428, 
        n45_adj_4429, n40860, n39185, n28146, n12_adj_4430, n14_adj_4431, 
        n15_adj_4432, n16_adj_4433, n17_adj_4434, n18_adj_4435, n19_adj_4436, 
        n20_adj_4437, n21_adj_4438, n23_adj_4439, n24_adj_4440, n25_adj_4441, 
        n27_adj_4442, n29_adj_4443, n40830, n31_adj_4444, n33_adj_4445, 
        n35_adj_4446, n37_adj_4447, n38_adj_4448, n39_adj_4449, n41_adj_4450, 
        n40668, n43_adj_4451, n40800, n40971, n39183, n39181, n28145, 
        n10_adj_4452, n12_adj_4453, n13_adj_4454, n14_adj_4455, n15_adj_4456, 
        n16_adj_4457, n17_adj_4458, n18_adj_4459, n19_adj_4460, n21_adj_4461, 
        n22_adj_4462, n23_adj_4463, n25_adj_4464, n27_adj_4465, n29_adj_4466, 
        n31_adj_4467, n33_adj_4468, n35_adj_4469, n36_adj_4470, n37_adj_4471, 
        n39_adj_4472, n41_adj_4473, n40972, n40483, n1679, n28144, 
        n3048, n28143, n8_adj_4474, n10_adj_4475, n11_adj_4476, n12_adj_4477, 
        n13_adj_4478, n14_adj_4479, n15_adj_4480, n16_adj_4481, n17_adj_4482, 
        n19_adj_4483, n20_adj_4484, n21_adj_4485, n23_adj_4486, n25_adj_4487, 
        n40481, n27_adj_4488, n29_adj_4489, n31_adj_4490, n33_adj_4491, 
        n34_adj_4492, n35_adj_4493, n37_adj_4494, n39_adj_4495, n40345, 
        n40666, n3039, n28142, n6_adj_4496, n8_adj_4497, n9_adj_4498, 
        n10_adj_4499, n11_adj_4500, n12_adj_4501, n13_adj_4502, n14_adj_4503, 
        n15_adj_4504, n17_adj_4505, n19_adj_4506, n21_adj_4507, n23_adj_4508, 
        n40472, n25_adj_4509, n40347, n27_adj_4510, n29_adj_4511, 
        n31_adj_4512, n32_adj_4513, n33_adj_4514, n35_adj_4515, n37_adj_4516, 
        n40885, n40848, n28141, n4_adj_4517, n6_adj_4518, n7_adj_4519, 
        n8_adj_4520, n9_adj_4521, n10_adj_4522, n11_adj_4523, n12_adj_4524, 
        n13_adj_4525, n15_adj_4526, n16_adj_4527, n17_adj_4528, n19_adj_4529, 
        n21_adj_4530, n40658, n23_adj_4531, n24_adj_4532, n25_adj_4533, 
        n27_adj_4534, n40656, n29_adj_4535, n30_adj_4536, n31_adj_4537, 
        n33_adj_4538, n35_adj_4539, n37_adj_4540, n40766, n39_adj_4541, 
        n40_adj_4542, n41_adj_4543, n43_adj_4544, n45_adj_4545, n40768, 
        n39691, n19_adj_4546, n39171, n39168, n35990, n28140, n28139, 
        n28138, n34616, n27586, n18308, n18307, n28137, n32678, 
        n40614, n28136, n37188, n40_adj_4547, n39_adj_4548, n39133, 
        n38_adj_4549, n37_adj_4550, n39131, n35_adj_4551, n34_adj_4552, 
        n28135, n40872, n39571, n5_adj_4553, n39127, n28134, n28_adj_4554, 
        n39125, n40671, n28133, n40363, n28132, n40514, n40369, 
        n28131, n28130, n40524, n28129, n28128, n28127, n40518, 
        n40513, n40675, n28126, n40974, n40393, n40667, n39095, 
        n39094, n39093, n28125, n28124, n39092, n39091, n39090, 
        n39089, n39088, n40516, n28123, n24_adj_4555, n40508, n21_adj_4556, 
        n20_adj_4557, n39087, n17_adj_4558, n28122, n39086, n39085, 
        n39084, n39083, n40506, n39082, n37153, n39081, n28121, 
        n39080, n40122, n39079, n28120, n40626, n39078, n28119, 
        n39077, n39076, n28118, n39075, n28117, n39074, n39073, 
        n28116, n39072, n28115, n39071, n28114, n40670, n40870, 
        n39070, n28113, n32_adj_4559, n31_adj_4560, n34612, n30_adj_4561, 
        n29_adj_4562, n28112, n28_adj_4563, n18306, n28111, n28110, 
        n28109, n39069, n39068, n39067, n39065, n28108, n21_adj_4564, 
        n39064, n17791, n39063, n39062, n40397, n28107, n28106, 
        n37047, n34618, n6_adj_4565, n27585, n28105, n34761, n40505, 
        n37033, n28104, n40968, n39047, n39045, n28103, n28102, 
        n28101, n39042, n39040, n39039, n39038, n28100, n40632, 
        n28099, n28098, n28097, n18305, n28096, n28095, n34725, 
        n18304, n18303, n28094, n18302, n28093, n28092, n18301, 
        n10_adj_4566, n34684, n40888, n39569, n36953, n40662, n6_adj_4567, 
        n40869, n28091, n28090, n28089, n28088, n40411, n6724, 
        n28087, n27584, n28086, n28085, n28084, n6769, n28083, 
        n28082, n28081, n16526, n40963, n28080, n40961, n39416, 
        n28079, n28078, n28077, n28076, n40958, n28075, n40947, 
        n28074, n28073, n28072, n28071, n27583, n40946, n28070, 
        n40415, n28069, n28068, n28067, n28066, n28065, n27582, 
        n27581, n40969, n40936, n40930, n40929, n28064, n28063, 
        n28062, n28061, n27802, n40924, n28060, n40962, n28059, 
        n28058, n28057, n28056, n28055, n28054, n40960, n40927, 
        n34344, n34342, n34642, n40902, n40937, n28053, n34678, 
        n40939, n2_adj_4568, n3_adj_4569, n4_adj_4570, n5_adj_4571, 
        n6_adj_4572, n7_adj_4573, n8_adj_4574, n9_adj_4575, n10_adj_4576, 
        n11_adj_4577, n12_adj_4578, n13_adj_4579, n14_adj_4580, n15_adj_4581, 
        n16_adj_4582, n17_adj_4583, n18_adj_4584, n19_adj_4585, n20_adj_4586, 
        n21_adj_4587, n22_adj_4588, n23_adj_4589, n24_adj_4590, n25_adj_4591, 
        n26_adj_4592, n27_adj_4593, n28_adj_4594, n29_adj_4595, n30_adj_4596, 
        n31_adj_4597, n33_adj_4598, n40849, n28052, n28051, n28050, 
        n27580, n40847, n40846, n28049, n27801, n28048, n28047, 
        n28046, n28045, n28044, n28043, n40836, n40833, n28042, 
        n28041, n28040, n28039, n40831, n40829, n28038, n28037, 
        n28036, n28035, n41713, n28034, n27713, n28033, n28032, 
        n27712, n28031, n28030, n28029, n40825, n28028, n27800, 
        n28027, n27711, n28026, n28025, n28024, n28023, n22_adj_4599, 
        n19_adj_4600, n18_adj_4601, n15_adj_4602, n28022, n27799, 
        n28021, n28020, n28019, n27798, n28018, n28017, n40819, 
        n28016, n28015, n28014, n36865, n28013, n28012, n28011, 
        n28010, n27710, n40815, n40813, n40642, n28009, n28008, 
        n28007, n40893, n40811, n40875, n38981, n28006, n28005, 
        n28004, n27797, n27579, n40975, n28003, n28002, n28001, 
        n40807, n28000, n27999, n27998, n40803, n27997, n27996, 
        n27995, n40894, n27994, n27993, n27796, n27992, n27991, 
        n27990, n27989, n27988, n27795, n27987, n27986, n40659, 
        n27985, n27984, n27983, n36316, n27982, n27981, n27794, 
        n27980, n40759, n27979, n27978, n40757, n27977, n32_adj_4603, 
        n39812, n40751, n29_adj_4604, n28_adj_4605, n40873, n40871, 
        n26_adj_4606, n40437, n20_adj_4607, n19_adj_4608, n36817, 
        n27976, n27975, n34659, n27793, n27974, n34672, n34555, 
        n27792, n27709, n27973, n27972, n27708, n40824, n27971, 
        n27970, n27969, n36797, n27791, n27968, n27967, n27966, 
        n27965, n27964, n27963, n27962, n27961, n27960, n27707, 
        n27959, n27958, n27957, n27956, n27955, n35420, n40439, 
        n27790, n27954, n27953, n27578, n27706, n27789, n27952, 
        n27705, n27951, n27950, n40657, n27949, n27948, n27947, 
        n37078, n33144, n40729, n27704, n27788, n27946, n27945, 
        n27577, n27944, n27943, n27942, n40727, n27941, n35752, 
        n27576, n27787, n27940, n27703, n27786, n27939, n27575, 
        n27574, n27938, n27937, n27936, n27935, n27934, n27785, 
        n27933, n40726, n27702, n27932, n40724, n27931, n27930, 
        n27929, n27573, n27572, n27928, n27927, n27926, n27784, 
        n27925, n27924, n27923, n27783, n27782, n27781, n27922, 
        n40828, n40719, n27921, n27920, n40717, n40832, n27919, 
        n27918, n40713, n27701, n36763, n36757, n27780, n40838, 
        n27917, n27916, n27915, n27914, n27913, n27912, n27911, 
        n27700, n27910, n27909, n33923, n27908, n27907, n34743, 
        n27906, n27905, n27904, n27903, n27902, n27901, n27900, 
        n27899, n27898, n27897, n39782, n36727, n27779, n34073, 
        n34651, n27896, n27895, n27699, n39709, n35922, n39780, 
        n23387, n27894, n27893, n27778, n39726, n27777, n27892, 
        n27776, n27698, n16405, n27891, n27890, n27889, n27775, 
        n27888, n27571, n34710, n36703, n36701, n39713, n36699, 
        n27887, n27886, n36697, n27697, n16420, n27696, n39722, 
        n36695, n27695, n27885, n36693, n27884, n34346, n8_adj_4609, 
        n27883, n27882, n27774, n27773, n4_adj_4610, n6_adj_4611, 
        n27694, n27881, n27880, n27879, n27878, n27877, n27693, 
        n27692, n27876, n27691, n27875, n27874, n37137, n27873, 
        n27872, n4_adj_4612, n27871, n27870, n27869, n27868, n27867, 
        n27866, n27865, n27864, n27863, n40609, n27862, n27861, 
        n36653, n36651, n40607, n27860, n16547, n27772, n36645, 
        n36643, n36641, n40594, n36629, n36625, n40588, n36621, 
        n20_adj_4613, n18_adj_4614, n16_adj_4615, n36615, n40674, 
        n36613, n36607, n34961, n41708, n19_adj_4616, n40565, n34307, 
        n39736, n34976, n40648, n40553, n18_adj_4617, n39673, n16_adj_4618, 
        n13_adj_4619, n5_adj_4620, n40343, n40254, n36485, n36483, 
        n36481, n36479, n36477, n33787, n42588, n33396, n36236, 
        n40212, n40455, n40498, n41718, n47_adj_4621, n46_adj_4622, 
        n40457, n40164, n40497, n36216;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 div_46_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4443));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_DFF h2_62 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_LUT4 i13447_3_lut (.I0(setpoint[21]), .I1(n4444), .I2(n36216), 
            .I3(GND_net), .O(n17954));   // verilog/coms.v(126[12] 289[6])
    defparam i13447_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_81[0]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_63 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF dir_67 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_LUT4 div_46_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i17_3_lut (.I0(n2949), .I1(n34_adj_4552), .I2(n2950), .I3(GND_net), 
            .O(n39_adj_4548));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    neopixel nx (.timer({timer}), .clk32MHz(clk32MHz), .n32678(n32678), 
            .VCC_net(VCC_net), .bit_ctr({bit_ctr}), .GND_net(GND_net), 
            .n32688(n32688), .n32680(n32680), .n32744(n32744), .n32746(n32746), 
            .n32748(n32748), .n32682(n32682), .n32734(n32734), .n32736(n32736), 
            .n32738(n32738), .n32742(n32742), .n32730(n32730), .n32732(n32732), 
            .n32726(n32726), .n32728(n32728), .n32722(n32722), .n32724(n32724), 
            .n32718(n32718), .n32720(n32720), .n32684(n32684), .start(start), 
            .n32716(n32716), .n32714(n32714), .n32686(n32686), .n39074(n39074), 
            .n19(n19_adj_4546), .n39095(n39095), .\state[0] (state[0]), 
            .n155(n155), .n39081(n39081), .n39092(n39092), .n39091(n39091), 
            .n39090(n39090), .\state[1] (state[1]), .n37153(n37153), .n39089(n39089), 
            .n39088(n39088), .n32712(n32712), .n18052(n18052), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n18051(n18051), .n18050(n18050), .n18049(n18049), .n18048(n18048), 
            .n18047(n18047), .n18046(n18046), .n18045(n18045), .n18044(n18044), 
            .n18043(n18043), .n18042(n18042), .n18041(n18041), .n18040(n18040), 
            .n18039(n18039), .n18038(n18038), .n18037(n18037), .n18036(n18036), 
            .n18035(n18035), .n18034(n18034), .n18033(n18033), .n18032(n18032), 
            .n18031(n18031), .n18030(n18030), .n18029(n18029), .n18028(n18028), 
            .n18027(n18027), .n18026(n18026), .n18025(n18025), .n18024(n18024), 
            .n18023(n18023), .n32710(n32710), .n32708(n32708), .n39080(n39080), 
            .n39087(n39087), .n39094(n39094), .n32702(n32702), .n32700(n32700), 
            .n32694(n32694), .n32698(n32698), .n32696(n32696), .n18000(n18000), 
            .n32692(n32692), .n39079(n39079), .n39086(n39086), .n39093(n39093), 
            .n39085(n39085), .n39070(n39070), .n32690(n32690), .n17922(n17922), 
            .n39084(n39084), .n39083(n39083), .n39069(n39069), .\state_3__N_337[1] (state_3__N_337[1]), 
            .n131(n131), .n17536(n17536), .n39082(n39082), .n21(n21_adj_3947), 
            .n17792(n17792), .n17561(n17561), .n17721(n17721), .n39078(n39078), 
            .n39077(n39077), .n39072(n39072), .n39071(n39071), .\color[16] (color[16]), 
            .\color[17] (color[17]), .\color[18] (color[18]), .\color[19] (color[19]), 
            .\color[22] (color[22]), .\color[23] (color[23]), .\color[20] (color[20]), 
            .\color[21] (color[21]), .n39067(n39067), .n39065(n39065), 
            .n39068(n39068), .n39073(n39073), .n39064(n39064), .PIN_8_c(PIN_8_c), 
            .n39063(n39063), .n39076(n39076), .n39075(n39075), .n175(n175), 
            .n39062(n39062)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(57[10] 63[2])
    SB_LUT4 i13448_3_lut (.I0(setpoint[20]), .I1(n4443), .I2(n36216), 
            .I3(GND_net), .O(n17955));   // verilog/coms.v(126[12] 289[6])
    defparam i13448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15_4_lut (.I0(n2943), .I1(n2944), .I2(n2952), .I3(n2947), 
            .O(n37_adj_4550));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13449_3_lut (.I0(setpoint[19]), .I1(n4442), .I2(n36216), 
            .I3(GND_net), .O(n17956));   // verilog/coms.v(126[12] 289[6])
    defparam i13449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3182_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n28061), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13450_3_lut (.I0(setpoint[18]), .I1(n4441), .I2(n36216), 
            .I3(GND_net), .O(n17957));   // verilog/coms.v(126[12] 289[6])
    defparam i13450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1854_21_lut (.I0(GND_net), .I1(n2739_adj_4095), 
            .I2(VCC_net), .I3(n28184), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13451_3_lut (.I0(setpoint[17]), .I1(n4440), .I2(n36216), 
            .I3(GND_net), .O(n17958));   // verilog/coms.v(126[12] 289[6])
    defparam i13451_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3182_9 (.CI(n28061), .I0(n2547), .I1(n93), .CO(n28062));
    SB_LUT4 i13452_3_lut (.I0(setpoint[16]), .I1(n4439), .I2(n36216), 
            .I3(GND_net), .O(n17959));   // verilog/coms.v(126[12] 289[6])
    defparam i13452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4218), .I3(n28400), .O(n20_adj_3991)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut (.I0(n37_adj_4550), .I1(n39_adj_4548), .I2(n38_adj_4549), 
            .I3(n40_adj_4547), .O(n2966));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13453_3_lut (.I0(setpoint[15]), .I1(n4438), .I2(n36216), 
            .I3(GND_net), .O(n17960));   // verilog/coms.v(126[12] 289[6])
    defparam i13453_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_1854_21 (.CI(n28184), .I0(n2739_adj_4095), 
            .I1(VCC_net), .CO(n28185));
    SB_LUT4 i13454_3_lut (.I0(setpoint[14]), .I1(n4437), .I2(n36216), 
            .I3(GND_net), .O(n17961));   // verilog/coms.v(126[12] 289[6])
    defparam i13454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3182_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n28060), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13943_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[5] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18450));   // verilog/coms.v(126[12] 289[6])
    defparam i13943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13455_3_lut (.I0(setpoint[13]), .I1(n4436), .I2(n36216), 
            .I3(GND_net), .O(n17962));   // verilog/coms.v(126[12] 289[6])
    defparam i13455_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_2_add_3_7 (.CI(n28400), .I0(GND_net), .I1(n20_adj_4218), 
            .CO(n28401));
    SB_LUT4 div_46_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4219), .I3(n28399), .O(n21_adj_3990)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_6 (.CI(n28399), .I0(GND_net), .I1(n21_adj_4219), 
            .CO(n28400));
    SB_LUT4 communication_counter_31__I_0_add_1854_20_lut (.I0(GND_net), .I1(n2740_adj_4094), 
            .I2(VCC_net), .I3(n28183), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4220), .I3(n28398), .O(n22_adj_3989)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_5 (.CI(n28398), .I0(GND_net), .I1(n22_adj_4220), 
            .CO(n28399));
    SB_LUT4 div_46_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4221), .I3(n28397), .O(n23_adj_3988)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_20 (.CI(n28183), .I0(n2740_adj_4094), 
            .I1(VCC_net), .CO(n28184));
    SB_CARRY div_46_unary_minus_2_add_3_4 (.CI(n28397), .I0(GND_net), .I1(n23_adj_4221), 
            .CO(n28398));
    SB_LUT4 div_46_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4222), .I3(n28396), .O(n24_adj_3987)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_3 (.CI(n28396), .I0(GND_net), .I1(n24_adj_4222), 
            .CO(n28397));
    SB_LUT4 communication_counter_31__I_0_add_1854_19_lut (.I0(GND_net), .I1(n2741_adj_4093), 
            .I2(VCC_net), .I3(n28182), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4223), .I3(VCC_net), .O(n25_adj_3986)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_19 (.CI(n28182), .I0(n2741_adj_4093), 
            .I1(VCC_net), .CO(n28183));
    SB_CARRY div_46_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4223), 
            .CO(n28396));
    SB_LUT4 communication_counter_31__I_0_add_1854_18_lut (.I0(GND_net), .I1(n2742_adj_4092), 
            .I2(VCC_net), .I3(n28181), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4176), .I3(n28395), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4177), .I3(n28394), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_18 (.CI(n28181), .I0(n2742_adj_4092), 
            .I1(VCC_net), .CO(n28182));
    SB_CARRY div_46_unary_minus_4_add_3_24 (.CI(n28394), .I0(GND_net), .I1(n3_adj_4177), 
            .CO(n28395));
    SB_LUT4 communication_counter_31__I_0_add_1854_17_lut (.I0(GND_net), .I1(n2743_adj_4091), 
            .I2(VCC_net), .I3(n28180), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_17 (.CI(n28180), .I0(n2743_adj_4091), 
            .I1(VCC_net), .CO(n28181));
    SB_LUT4 div_46_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4178), .I3(n28393), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_23 (.CI(n28393), .I0(GND_net), .I1(n4_adj_4178), 
            .CO(n28394));
    SB_LUT4 communication_counter_31__I_0_add_1854_16_lut (.I0(GND_net), .I1(n2744_adj_4090), 
            .I2(VCC_net), .I3(n28179), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4179), .I3(n28392), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_22 (.CI(n28392), .I0(GND_net), .I1(n5_adj_4179), 
            .CO(n28393));
    SB_CARRY communication_counter_31__I_0_add_1854_16 (.CI(n28179), .I0(n2744_adj_4090), 
            .I1(VCC_net), .CO(n28180));
    SB_LUT4 div_46_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4180), .I3(n28391), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_21 (.CI(n28391), .I0(GND_net), .I1(n6_adj_4180), 
            .CO(n28392));
    SB_LUT4 div_46_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4181), .I3(n28390), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_15_lut (.I0(GND_net), .I1(n2745_adj_4089), 
            .I2(VCC_net), .I3(n28178), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_20 (.CI(n28390), .I0(GND_net), .I1(n7_adj_4181), 
            .CO(n28391));
    SB_LUT4 div_46_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4182), .I3(n28389), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_15 (.CI(n28178), .I0(n2745_adj_4089), 
            .I1(VCC_net), .CO(n28179));
    SB_LUT4 add_3182_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n28066), 
            .O(n6894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_14 (.CI(n28066), .I0(n2542), .I1(n88), .CO(n28067));
    SB_LUT4 i13456_3_lut (.I0(setpoint[12]), .I1(n4435), .I2(n36216), 
            .I3(GND_net), .O(n17963));   // verilog/coms.v(126[12] 289[6])
    defparam i13456_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_4_add_3_19 (.CI(n28389), .I0(GND_net), .I1(n8_adj_4182), 
            .CO(n28390));
    SB_LUT4 div_46_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4183), .I3(n28388), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_14_lut (.I0(GND_net), .I1(n2746_adj_4088), 
            .I2(VCC_net), .I3(n28177), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_14 (.CI(n28177), .I0(n2746_adj_4088), 
            .I1(VCC_net), .CO(n28178));
    SB_LUT4 add_3182_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n28065), 
            .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1806_3_lut (.I0(n2653), .I1(n2720_adj_4102), 
            .I2(n2669), .I3(GND_net), .O(n2752_adj_4082));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1854_13_lut (.I0(GND_net), .I1(n2747_adj_4087), 
            .I2(VCC_net), .I3(n28176), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13942_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[5] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18449));   // verilog/coms.v(126[12] 289[6])
    defparam i13942_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_4_add_3_18 (.CI(n28388), .I0(GND_net), .I1(n9_adj_4183), 
            .CO(n28389));
    SB_LUT4 div_46_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4184), .I3(n28387), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13457_3_lut (.I0(setpoint[11]), .I1(n4434), .I2(n36216), 
            .I3(GND_net), .O(n17964));   // verilog/coms.v(126[12] 289[6])
    defparam i13457_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_46_unary_minus_4_add_3_17 (.CI(n28387), .I0(GND_net), .I1(n10_adj_4184), 
            .CO(n28388));
    SB_CARRY communication_counter_31__I_0_add_1854_13 (.CI(n28176), .I0(n2747_adj_4087), 
            .I1(VCC_net), .CO(n28177));
    SB_LUT4 i13458_3_lut (.I0(setpoint[10]), .I1(n4433), .I2(n36216), 
            .I3(GND_net), .O(n17965));   // verilog/coms.v(126[12] 289[6])
    defparam i13458_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3182_13 (.CI(n28065), .I0(n2543), .I1(n89), .CO(n28066));
    SB_LUT4 div_46_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4185), .I3(n28386), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3182_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n28064), 
            .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4568));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13676_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13950), .I3(GND_net), .O(n18183));   // verilog/coms.v(126[12] 289[6])
    defparam i13676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13459_3_lut (.I0(setpoint[9]), .I1(n4432), .I2(n36216), .I3(GND_net), 
            .O(n17966));   // verilog/coms.v(126[12] 289[6])
    defparam i13459_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13460_3_lut (.I0(setpoint[8]), .I1(n4431), .I2(n36216), .I3(GND_net), 
            .O(n17967));   // verilog/coms.v(126[12] 289[6])
    defparam i13460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13461_3_lut (.I0(setpoint[7]), .I1(n4430), .I2(n36216), .I3(GND_net), 
            .O(n17968));   // verilog/coms.v(126[12] 289[6])
    defparam i13461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13462_3_lut (.I0(setpoint[6]), .I1(n4429), .I2(n36216), .I3(GND_net), 
            .O(n17969));   // verilog/coms.v(126[12] 289[6])
    defparam i13462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13859_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n33775), .I3(GND_net), .O(n18366));   // verilog/coms.v(126[12] 289[6])
    defparam i13859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13463_3_lut (.I0(setpoint[5]), .I1(n4428), .I2(n36216), .I3(GND_net), 
            .O(n17970));   // verilog/coms.v(126[12] 289[6])
    defparam i13463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13941_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[5] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18448));   // verilog/coms.v(126[12] 289[6])
    defparam i13941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13677_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13950), .I3(GND_net), .O(n18184));   // verilog/coms.v(126[12] 289[6])
    defparam i13677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4191));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13464_3_lut (.I0(setpoint[4]), .I1(n4427), .I2(n36216), .I3(GND_net), 
            .O(n17971));   // verilog/coms.v(126[12] 289[6])
    defparam i13464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1653_3_lut (.I0(n2458), .I1(n6875), .I2(n2471), .I3(GND_net), 
            .O(n2545));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13940_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[5] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18447));   // verilog/coms.v(126[12] 289[6])
    defparam i13940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13465_3_lut (.I0(setpoint[3]), .I1(n4426), .I2(n36216), .I3(GND_net), 
            .O(n17972));   // verilog/coms.v(126[12] 289[6])
    defparam i13465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i963_3_lut (.I0(n1413), .I1(n6700), .I2(n1436), .I3(GND_net), 
            .O(n1530));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13466_3_lut (.I0(setpoint[2]), .I1(n4425), .I2(n36216), .I3(GND_net), 
            .O(n17973));   // verilog/coms.v(126[12] 289[6])
    defparam i13466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4190));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13678_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13950), .I3(GND_net), .O(n18185));   // verilog/coms.v(126[12] 289[6])
    defparam i13678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13954_3_lut (.I0(encoder0_position[11]), .I1(n2744), .I2(count_enable), 
            .I3(GND_net), .O(n18461));   // quad.v(35[10] 41[6])
    defparam i13954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[6]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_107[6]), 
            .I2(n15), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13953_3_lut (.I0(encoder0_position[10]), .I1(n2745), .I2(count_enable), 
            .I3(GND_net), .O(n18460));   // quad.v(35[10] 41[6])
    defparam i13953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3932));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13679_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13950), .I3(GND_net), .O(n18186));   // verilog/coms.v(126[12] 289[6])
    defparam i13679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13952_3_lut (.I0(encoder0_position[9]), .I1(n2746), .I2(count_enable), 
            .I3(GND_net), .O(n18459));   // quad.v(35[10] 41[6])
    defparam i13952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13951_3_lut (.I0(encoder0_position[8]), .I1(n2747), .I2(count_enable), 
            .I3(GND_net), .O(n18458));   // quad.v(35[10] 41[6])
    defparam i13951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13680_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13950), .I3(GND_net), .O(n18187));   // verilog/coms.v(126[12] 289[6])
    defparam i13680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i41_4_lut (.I0(n2702_adj_4068), .I1(n80), 
            .I2(n6936), .I3(n2724), .O(n41_adj_4543));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i39_4_lut (.I0(n2703_adj_4069), .I1(n81), 
            .I2(n6937), .I3(n2724), .O(n39_adj_4541));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_3986), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13950_3_lut (.I0(encoder0_position[7]), .I1(n2748), .I2(count_enable), 
            .I3(GND_net), .O(n18457));   // quad.v(35[10] 41[6])
    defparam i13950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13949_3_lut (.I0(encoder0_position[6]), .I1(n2749), .I2(count_enable), 
            .I3(GND_net), .O(n18456));   // quad.v(35[10] 41[6])
    defparam i13949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i45_4_lut (.I0(n2700_adj_4066), .I1(n78), 
            .I2(n6934), .I3(n2724), .O(n45_adj_4545));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13948_3_lut (.I0(encoder0_position[5]), .I1(n2750), .I2(count_enable), 
            .I3(GND_net), .O(n18455));   // quad.v(35[10] 41[6])
    defparam i13948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13681_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13950), .I3(GND_net), .O(n18188));   // verilog/coms.v(126[12] 289[6])
    defparam i13681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i43_4_lut (.I0(n2701_adj_4067), .I1(n79), 
            .I2(n6935), .I3(n2724), .O(n43_adj_4544));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i37_4_lut (.I0(n2704_adj_4070), .I1(n82), 
            .I2(n6938), .I3(n2724), .O(n37_adj_4540));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13947_3_lut (.I0(encoder0_position[4]), .I1(n2751), .I2(count_enable), 
            .I3(GND_net), .O(n18454));   // quad.v(35[10] 41[6])
    defparam i13947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13946_3_lut (.I0(encoder0_position[3]), .I1(n2752), .I2(count_enable), 
            .I3(GND_net), .O(n18453));   // quad.v(35[10] 41[6])
    defparam i13946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6942), 
            .I3(n2724), .O(n29_adj_4535));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6941), 
            .I3(n2724), .O(n31_adj_4537));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6946), 
            .I3(n2724), .O(n21_adj_4530));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6945), 
            .I3(n2724), .O(n23_adj_4531));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY div_46_unary_minus_4_add_3_16 (.CI(n28386), .I0(GND_net), .I1(n11_adj_4185), 
            .CO(n28387));
    SB_LUT4 div_46_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6944), 
            .I3(n2724), .O(n25_adj_4533));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13958_3_lut (.I0(encoder0_position[15]), .I1(n2740), .I2(count_enable), 
            .I3(GND_net), .O(n18465));   // quad.v(35[10] 41[6])
    defparam i13958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6948), 
            .I3(n2724), .O(n17_adj_4528));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13957_3_lut (.I0(encoder0_position[14]), .I1(n2741), .I2(count_enable), 
            .I3(GND_net), .O(n18464));   // quad.v(35[10] 41[6])
    defparam i13957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13956_3_lut (.I0(encoder0_position[13]), .I1(n2742), .I2(count_enable), 
            .I3(GND_net), .O(n18463));   // quad.v(35[10] 41[6])
    defparam i13956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6947), 
            .I3(n2724), .O(n19_adj_4529));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY add_3182_8 (.CI(n28060), .I0(n2548), .I1(n94), .CO(n28061));
    SB_LUT4 i13955_3_lut (.I0(encoder0_position[12]), .I1(n2743), .I2(count_enable), 
            .I3(GND_net), .O(n18462));   // quad.v(35[10] 41[6])
    defparam i13955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6952), 
            .I3(n2724), .O(n9_adj_4521));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i18892_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[22] [0]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n23387));   // verilog/coms.v(100[12:33])
    defparam i18892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6953), 
            .I3(n2724), .O(n7_adj_4519));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13966_3_lut (.I0(encoder0_position[23]), .I1(n2732), .I2(count_enable), 
            .I3(GND_net), .O(n18473));   // quad.v(35[10] 41[6])
    defparam i13966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18895_4_lut (.I0(n23387), .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(byte_transmit_counter[1]), .O(n21_adj_4564));   // verilog/coms.v(100[12:33])
    defparam i18895_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13965_3_lut (.I0(encoder0_position[22]), .I1(n2733), .I2(count_enable), 
            .I3(GND_net), .O(n18472));   // quad.v(35[10] 41[6])
    defparam i13965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13860_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n33775), .I3(GND_net), .O(n18367));   // verilog/coms.v(126[12] 289[6])
    defparam i13860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1830_i35_4_lut (.I0(n2705_adj_4071), .I1(n83), 
            .I2(n6939), .I3(n2724), .O(n35_adj_4539));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i13976_3_lut (.I0(encoder1_position[9]), .I1(n2696), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18483));   // quad.v(35[10] 41[6])
    defparam i13976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13975_3_lut (.I0(encoder1_position[8]), .I1(n2697), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18482));   // quad.v(35[10] 41[6])
    defparam i13975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13974_3_lut (.I0(encoder1_position[7]), .I1(n2698), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18481));   // quad.v(35[10] 41[6])
    defparam i13974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6951), 
            .I3(n2724), .O(n11_adj_4523));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6950), 
            .I3(n2724), .O(n13_adj_4525));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6943), 
            .I3(n2724), .O(n27_adj_4534));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6949), 
            .I3(n2724), .O(n15_adj_4526));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6940), 
            .I3(n2724), .O(n33_adj_4538));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1595_3_lut (.I0(n2369), .I1(n6855), .I2(n2381), .I3(GND_net), 
            .O(n2459));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1595_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13978_3_lut (.I0(encoder1_position[11]), .I1(n2694), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18485));   // quad.v(35[10] 41[6])
    defparam i13978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1854_12_lut (.I0(GND_net), .I1(n2748_adj_4086), 
            .I2(VCC_net), .I3(n28175), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32945_4_lut (.I0(n27_adj_4534), .I1(n15_adj_4526), .I2(n13_adj_4525), 
            .I3(n11_adj_4523), .O(n39265));
    defparam i32945_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4538), 
            .I3(GND_net), .O(n12_adj_4524));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_3182_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n28059), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13977_3_lut (.I0(encoder1_position[10]), .I1(n2695), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18484));   // quad.v(35[10] 41[6])
    defparam i13977_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1854_12 (.CI(n28175), .I0(n2748_adj_4086), 
            .I1(VCC_net), .CO(n28176));
    SB_LUT4 i32892_2_lut (.I0(n33_adj_4538), .I1(n15_adj_4526), .I2(GND_net), 
            .I3(GND_net), .O(n39212));
    defparam i32892_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13980_3_lut (.I0(encoder1_position[13]), .I1(n2692), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18487));   // quad.v(35[10] 41[6])
    defparam i13980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13979_3_lut (.I0(encoder1_position[12]), .I1(n2693), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18486));   // quad.v(35[10] 41[6])
    defparam i13979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4525), 
            .I3(GND_net), .O(n10_adj_4522));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13982_3_lut (.I0(encoder1_position[15]), .I1(n2690), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18489));   // quad.v(35[10] 41[6])
    defparam i13982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13981_3_lut (.I0(encoder1_position[14]), .I1(n2691), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18488));   // quad.v(35[10] 41[6])
    defparam i13981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13984_3_lut (.I0(encoder1_position[17]), .I1(n2688), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18491));   // quad.v(35[10] 41[6])
    defparam i13984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13983_3_lut (.I0(encoder1_position[16]), .I1(n2689), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18490));   // quad.v(35[10] 41[6])
    defparam i13983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13986_3_lut (.I0(encoder1_position[19]), .I1(n2686), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18493));   // quad.v(35[10] 41[6])
    defparam i13986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i30_3_lut (.I0(n12_adj_4524), .I1(n83), 
            .I2(n35_adj_4539), .I3(GND_net), .O(n30_adj_4536));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1828_3_lut (.I0(n2720), .I1(n6954), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13985_3_lut (.I0(encoder1_position[18]), .I1(n2687), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18492));   // quad.v(35[10] 41[6])
    defparam i13985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32986_3_lut (.I0(n7_adj_4519), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n39306));
    defparam i32986_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i33582_4_lut (.I0(n13_adj_4525), .I1(n11_adj_4523), .I2(n9_adj_4521), 
            .I3(n39306), .O(n39904));
    defparam i33582_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i13917_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18424));   // verilog/coms.v(126[12] 289[6])
    defparam i13917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13916_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18423));   // verilog/coms.v(126[12] 289[6])
    defparam i13916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33574_4_lut (.I0(n19_adj_4529), .I1(n17_adj_4528), .I2(n15_adj_4526), 
            .I3(n39904), .O(n39896));
    defparam i33574_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34402_4_lut (.I0(n25_adj_4533), .I1(n23_adj_4531), .I2(n21_adj_4530), 
            .I3(n39896), .O(n40724));
    defparam i34402_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33982_4_lut (.I0(n31_adj_4537), .I1(n29_adj_4535), .I2(n27_adj_4534), 
            .I3(n40724), .O(n40304));
    defparam i33982_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i13682_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13950), .I3(GND_net), .O(n18189));   // verilog/coms.v(126[12] 289[6])
    defparam i13682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13683_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13950), .I3(GND_net), .O(n18190));   // verilog/coms.v(126[12] 289[6])
    defparam i13683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34528_4_lut (.I0(n37_adj_4540), .I1(n35_adj_4539), .I2(n33_adj_4538), 
            .I3(n40304), .O(n40850));
    defparam i34528_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4544), 
            .I3(GND_net), .O(n16_adj_4527));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4519), 
            .I3(GND_net), .O(n6_adj_4518));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13915_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18422));   // verilog/coms.v(126[12] 289[6])
    defparam i13915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34336_3_lut (.I0(n6_adj_4518), .I1(n90), .I2(n21_adj_4530), 
            .I3(GND_net), .O(n40658));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34336_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34337_3_lut (.I0(n40658), .I1(n89), .I2(n23_adj_4531), .I3(GND_net), 
            .O(n40659));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34337_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32957_4_lut (.I0(n21_adj_4530), .I1(n19_adj_4529), .I2(n17_adj_4528), 
            .I3(n9_adj_4521), .O(n39277));
    defparam i32957_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32865_2_lut (.I0(n43_adj_4544), .I1(n19_adj_4529), .I2(GND_net), 
            .I3(GND_net), .O(n39185));
    defparam i32865_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4528), 
            .I3(GND_net), .O(n8_adj_4520));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i24_3_lut (.I0(n16_adj_4527), .I1(n78), 
            .I2(n45_adj_4545), .I3(GND_net), .O(n24_adj_4532));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32867_4_lut (.I0(n43_adj_4544), .I1(n25_adj_4533), .I2(n23_adj_4531), 
            .I3(n39277), .O(n39187));
    defparam i32867_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34025_4_lut (.I0(n24_adj_4532), .I1(n8_adj_4520), .I2(n45_adj_4545), 
            .I3(n39185), .O(n40347));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34025_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34285_3_lut (.I0(n40659), .I1(n88), .I2(n25_adj_4533), .I3(GND_net), 
            .O(n40607));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34285_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1829_3_lut (.I0(n390), .I1(n6955), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13684_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13950), .I3(GND_net), .O(n18191));   // verilog/coms.v(126[12] 289[6])
    defparam i13684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4189));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13914_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18421));   // verilog/coms.v(126[12] 289[6])
    defparam i13914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4517));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34334_3_lut (.I0(n4_adj_4517), .I1(n87), .I2(n27_adj_4534), 
            .I3(GND_net), .O(n40656));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34334_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34335_3_lut (.I0(n40656), .I1(n86), .I2(n29_adj_4535), .I3(GND_net), 
            .O(n40657));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34335_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32906_4_lut (.I0(n33_adj_4538), .I1(n31_adj_4537), .I2(n29_adj_4535), 
            .I3(n39265), .O(n39226));
    defparam i32906_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34563_4_lut (.I0(n30_adj_4536), .I1(n10_adj_4522), .I2(n35_adj_4539), 
            .I3(n39212), .O(n40885));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34563_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34287_3_lut (.I0(n40657), .I1(n85), .I2(n31_adj_4537), .I3(GND_net), 
            .O(n40609));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34287_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34638_4_lut (.I0(n40609), .I1(n40885), .I2(n35_adj_4539), 
            .I3(n39226), .O(n40960));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34638_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34639_3_lut (.I0(n40960), .I1(n82), .I2(n37_adj_4540), .I3(GND_net), 
            .O(n40961));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34639_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34602_3_lut (.I0(n40961), .I1(n81), .I2(n39_adj_4541), .I3(GND_net), 
            .O(n40924));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34602_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32869_4_lut (.I0(n43_adj_4544), .I1(n41_adj_4543), .I2(n39_adj_4541), 
            .I3(n40850), .O(n39189));
    defparam i32869_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34444_4_lut (.I0(n40607), .I1(n40347), .I2(n45_adj_4545), 
            .I3(n39187), .O(n40766));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34444_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34593_3_lut (.I0(n40924), .I1(n80), .I2(n41_adj_4543), .I3(GND_net), 
            .O(n40_adj_4542));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34593_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13926_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[7] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18433));   // verilog/coms.v(126[12] 289[6])
    defparam i13926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1807_3_lut (.I0(n2699_adj_4065), .I1(n6933), .I2(n2724), 
            .I3(GND_net), .O(n2777));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_3989), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_106));   // verilog/TinyFPGA_B.v(166[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34446_4_lut (.I0(n40_adj_4542), .I1(n40766), .I2(n45_adj_4545), 
            .I3(n39189), .O(n40768));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34446_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34447_3_lut (.I0(n40768), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34447_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30901_1_lut (.I0(n36607), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36629));
    defparam i30901_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13925_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[7] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18432));   // verilog/coms.v(126[12] 289[6])
    defparam i13925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1805_3_lut (.I0(n2652), .I1(n2719_adj_4103), 
            .I2(n2669), .I3(GND_net), .O(n2751_adj_4083));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13924_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[7] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18431));   // verilog/coms.v(126[12] 289[6])
    defparam i13924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1661_3_lut (.I0(n387), .I1(n6883), .I2(n2471), .I3(GND_net), 
            .O(n2553));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13923_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[7] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18430));   // verilog/coms.v(126[12] 289[6])
    defparam i13923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4514));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4512));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4188));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1777_i37_2_lut (.I0(n2704_adj_4070), .I1(n83), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4516));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1040_3_lut (.I0(n1530), .I1(n6712), .I2(n1553), .I3(GND_net), 
            .O(n1644));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13922_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[7] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18429));   // verilog/coms.v(126[12] 289[6])
    defparam i13922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1777_i35_2_lut (.I0(n2705_adj_4071), .I1(n84), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4515));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13921_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[7] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18428));   // verilog/coms.v(126[12] 289[6])
    defparam i13921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_3987), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13685_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13950), .I3(GND_net), .O(n18192));   // verilog/coms.v(126[12] 289[6])
    defparam i13685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4509));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1660_3_lut (.I0(n2465), .I1(n6882), .I2(n2471), .I3(GND_net), 
            .O(n2552));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13920_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18427));   // verilog/coms.v(126[12] 289[6])
    defparam i13920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13686_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13950), .I3(GND_net), .O(n18193));   // verilog/coms.v(126[12] 289[6])
    defparam i13686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_3_lut (.I0(bit_ctr[16]), .I1(n39067), .I2(n17536), .I3(GND_net), 
            .O(n32686));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4510));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4507));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4508));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1854_11_lut (.I0(GND_net), .I1(n2749_adj_4085), 
            .I2(VCC_net), .I3(n28174), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1115_3_lut (.I0(n1644), .I1(n6725), .I2(n1667), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4498));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4500));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4506));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4186), .I3(n28385), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_15 (.CI(n28385), .I0(GND_net), .I1(n12_adj_4186), 
            .CO(n28386));
    SB_LUT4 div_46_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4187), .I3(n28384), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_7 (.CI(n28059), .I0(n2549), .I1(n95), .CO(n28060));
    SB_LUT4 div_46_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4502));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1854_11 (.CI(n28174), .I0(n2749_adj_4085), 
            .I1(VCC_net), .CO(n28175));
    SB_LUT4 div_46_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4504));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4505));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4511));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3182_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n28058), 
            .O(n6902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_10_lut (.I0(GND_net), .I1(n2750_adj_4084), 
            .I2(VCC_net), .I3(n28173), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33094_4_lut (.I0(n29_adj_4511), .I1(n17_adj_4505), .I2(n15_adj_4504), 
            .I3(n13_adj_4502), .O(n39416));
    defparam i33094_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY div_46_unary_minus_4_add_3_14 (.CI(n28384), .I0(GND_net), .I1(n13_adj_4187), 
            .CO(n28385));
    SB_CARRY add_3182_6 (.CI(n28058), .I0(n2550), .I1(n96), .CO(n28059));
    SB_LUT4 add_3182_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n28057), 
            .O(n6903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33730_4_lut (.I0(n11_adj_4500), .I1(n9_adj_4498), .I2(n2719), 
            .I3(n98), .O(n40052));
    defparam i33730_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY add_3182_5 (.CI(n28057), .I0(n2551), .I1(n97), .CO(n28058));
    SB_LUT4 i13991_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n34976), 
            .I3(GND_net), .O(n18498));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3182_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n28056), 
            .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34047_4_lut (.I0(n17_adj_4505), .I1(n15_adj_4504), .I2(n13_adj_4502), 
            .I3(n40052), .O(n40369));
    defparam i34047_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34041_4_lut (.I0(n23_adj_4508), .I1(n21_adj_4507), .I2(n19_adj_4506), 
            .I3(n40369), .O(n40363));
    defparam i34041_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33096_4_lut (.I0(n29_adj_4511), .I1(n27_adj_4510), .I2(n25_adj_4509), 
            .I3(n40363), .O(n39418));
    defparam i33096_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4496));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34147_3_lut (.I0(n6_adj_4496), .I1(n87), .I2(n29_adj_4511), 
            .I3(GND_net), .O(n40469));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34147_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13990_3_lut (.I0(encoder1_position[23]), .I1(n2682), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18497));   // quad.v(35[10] 41[6])
    defparam i13990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13989_3_lut (.I0(encoder1_position[22]), .I1(n2683), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18496));   // quad.v(35[10] 41[6])
    defparam i13989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i32_3_lut (.I0(n14_adj_4503), .I1(n83), 
            .I2(n37_adj_4516), .I3(GND_net), .O(n32_adj_4513));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4188), .I3(n28383), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_12 (.CI(n28064), .I0(n2544), .I1(n90), .CO(n28065));
    SB_CARRY add_3182_4 (.CI(n28056), .I0(n2552), .I1(n98), .CO(n28057));
    SB_CARRY div_46_unary_minus_4_add_3_13 (.CI(n28383), .I0(GND_net), .I1(n14_adj_4188), 
            .CO(n28384));
    SB_CARRY communication_counter_31__I_0_add_1854_10 (.CI(n28173), .I0(n2750_adj_4084), 
            .I1(VCC_net), .CO(n28174));
    SB_LUT4 add_3182_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n28055), 
            .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_3 (.CI(n28055), .I0(n2553), .I1(n99), .CO(n28056));
    SB_LUT4 communication_counter_31__I_0_add_1854_9_lut (.I0(GND_net), .I1(n2751_adj_4083), 
            .I2(VCC_net), .I3(n28172), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3182_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34148_3_lut (.I0(n40469), .I1(n86), .I2(n31_adj_4512), .I3(GND_net), 
            .O(n40470));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34148_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4189), .I3(n28382), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_12 (.CI(n28382), .I0(GND_net), .I1(n15_adj_4189), 
            .CO(n28383));
    SB_LUT4 i33049_4_lut (.I0(n35_adj_4515), .I1(n33_adj_4514), .I2(n31_adj_4512), 
            .I3(n39416), .O(n39370));
    defparam i33049_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34561_4_lut (.I0(n32_adj_4513), .I1(n12_adj_4501), .I2(n37_adj_4516), 
            .I3(n39368), .O(n40883));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34561_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33681_3_lut (.I0(n40470), .I1(n85), .I2(n33_adj_4514), .I3(GND_net), 
            .O(n40003));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33681_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34149_3_lut (.I0(n8_adj_4497), .I1(n90), .I2(n23_adj_4508), 
            .I3(GND_net), .O(n40471));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34149_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14005_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1035), .I3(GND_net), .O(n18512));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34150_3_lut (.I0(n40471), .I1(n89), .I2(n25_adj_4509), .I3(GND_net), 
            .O(n40472));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34150_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i22_3_lut (.I0(bit_ctr[8]), .I1(n39079), .I2(n17536), .I3(GND_net), 
            .O(n32714));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33706_4_lut (.I0(n25_adj_4509), .I1(n23_adj_4508), .I2(n21_adj_4507), 
            .I3(n39436), .O(n40028));
    defparam i33706_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34023_3_lut (.I0(n10_adj_4499), .I1(n91), .I2(n21_adj_4507), 
            .I3(GND_net), .O(n40345));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34023_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33679_3_lut (.I0(n40472), .I1(n88), .I2(n27_adj_4510), .I3(GND_net), 
            .O(n40001));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33679_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34292_4_lut (.I0(n35_adj_4515), .I1(n33_adj_4514), .I2(n31_adj_4512), 
            .I3(n39418), .O(n40614));
    defparam i34292_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34636_4_lut (.I0(n40003), .I1(n40883), .I2(n37_adj_4516), 
            .I3(n39370), .O(n40958));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34636_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34340_4_lut (.I0(n40001), .I1(n40345), .I2(n27_adj_4510), 
            .I3(n40028), .O(n40662));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34340_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34650_4_lut (.I0(n40662), .I1(n40958), .I2(n37_adj_4516), 
            .I3(n40614), .O(n40972));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34650_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34651_3_lut (.I0(n40972), .I1(n82), .I2(n2703_adj_4069), 
            .I3(GND_net), .O(n40973));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34651_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34645_3_lut (.I0(n40973), .I1(n81), .I2(n2702_adj_4068), 
            .I3(GND_net), .O(n40967));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34645_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34524_3_lut (.I0(n40967), .I1(n80), .I2(n2701_adj_4067), 
            .I3(GND_net), .O(n40846));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34524_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i13945_3_lut (.I0(encoder0_position[2]), .I1(n2753), .I2(count_enable), 
            .I3(GND_net), .O(n18452));   // quad.v(35[10] 41[6])
    defparam i13945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13944_3_lut (.I0(encoder0_position[1]), .I1(n2754), .I2(count_enable), 
            .I3(GND_net), .O(n18451));   // quad.v(35[10] 41[6])
    defparam i13944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34525_3_lut (.I0(n40846), .I1(n79), .I2(n2700_adj_4066), 
            .I3(GND_net), .O(n40847));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34525_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1983_4_lut (.I0(n40847), .I1(n77), .I2(n78), .I3(n2699_adj_4065), 
            .O(n2723));
    defparam i1983_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i13467_3_lut (.I0(setpoint[1]), .I1(n4424), .I2(n36216), .I3(GND_net), 
            .O(n17974));   // verilog/coms.v(126[12] 289[6])
    defparam i13467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1512 (.I0(bit_ctr[9]), .I1(n39080), .I2(n17536), 
            .I3(GND_net), .O(n32716));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1512.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4190), .I3(n28381), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_11 (.CI(n28381), .I0(GND_net), .I1(n16_adj_4190), 
            .CO(n28382));
    SB_LUT4 add_3182_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n28063), 
            .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4191), .I3(n28380), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_10 (.CI(n28380), .I0(GND_net), .I1(n17_adj_4191), 
            .CO(n28381));
    SB_LUT4 div_46_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4493));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1854_9 (.CI(n28172), .I0(n2751_adj_4083), 
            .I1(VCC_net), .CO(n28173));
    SB_LUT4 div_46_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4495));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4491));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_3988), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4494));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1854_8_lut (.I0(GND_net), .I1(n2752_adj_4082), 
            .I2(VCC_net), .I3(n28171), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_8 (.CI(n28171), .I0(n2752_adj_4082), 
            .I1(VCC_net), .CO(n28172));
    SB_CARRY add_3182_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n28055));
    SB_LUT4 div_46_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4488));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1988_27_lut (.I0(n2966), .I1(n2933), 
            .I2(VCC_net), .I3(n28054), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3182_11 (.CI(n28063), .I0(n2545), .I1(n91), .CO(n28064));
    SB_LUT4 div_46_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4489));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1988_26_lut (.I0(GND_net), .I1(n2934), 
            .I2(VCC_net), .I3(n28053), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_26 (.CI(n28053), .I0(n2934), 
            .I1(VCC_net), .CO(n28054));
    SB_LUT4 communication_counter_31__I_0_add_1988_25_lut (.I0(GND_net), .I1(n2935), 
            .I2(VCC_net), .I3(n28052), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4192), .I3(n28379), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_25 (.CI(n28052), .I0(n2935), 
            .I1(VCC_net), .CO(n28053));
    SB_LUT4 communication_counter_31__I_0_add_1988_24_lut (.I0(GND_net), .I1(n2936), 
            .I2(VCC_net), .I3(n28051), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_24 (.CI(n28051), .I0(n2936), 
            .I1(VCC_net), .CO(n28052));
    SB_LUT4 add_3182_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n28062), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_7_lut (.I0(GND_net), .I1(n2753_adj_4081), 
            .I2(VCC_net), .I3(n28170), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_9 (.CI(n28379), .I0(GND_net), .I1(n18_adj_4192), 
            .CO(n28380));
    SB_LUT4 add_555_24_lut (.I0(duty[22]), .I1(n41708), .I2(n3), .I3(n27589), 
            .O(pwm_setpoint_22__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_555_23_lut (.I0(duty[21]), .I1(n41708), .I2(n4_adj_3930), 
            .I3(n27588), .O(pwm_setpoint_22__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4486));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i18_4_lut (.I0(n175), .I1(n155), .I2(state[1]), .I3(start), 
            .O(n32684));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 div_46_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4487));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4193), .I3(n28378), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1513 (.I0(bit_ctr[21]), .I1(n39082), .I2(n17536), 
            .I3(GND_net), .O(n32720));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1513.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_8 (.CI(n28378), .I0(GND_net), .I1(n19_adj_4193), 
            .CO(n28379));
    SB_LUT4 communication_counter_31__I_0_add_1988_23_lut (.I0(GND_net), .I1(n2937), 
            .I2(VCC_net), .I3(n28050), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_23 (.CI(n27588), .I0(n41708), .I1(n4_adj_3930), .CO(n27589));
    SB_LUT4 div_46_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4194), .I3(n28377), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4476));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1188_3_lut (.I0(n1755), .I1(n6739), .I2(n1778), .I3(GND_net), 
            .O(n1863));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4478));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4485));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1514 (.I0(bit_ctr[10]), .I1(n39081), .I2(n17536), 
            .I3(GND_net), .O(n32718));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1514.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1515 (.I0(bit_ctr[23]), .I1(n39084), .I2(n17536), 
            .I3(GND_net), .O(n32724));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1515.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1516 (.I0(bit_ctr[22]), .I1(n39083), .I2(n17536), 
            .I3(GND_net), .O(n32722));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1516.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4480));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1517 (.I0(bit_ctr[25]), .I1(n39086), .I2(n17536), 
            .I3(GND_net), .O(n32728));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1517.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4482));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4483));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1518 (.I0(bit_ctr[24]), .I1(n39085), .I2(n17536), 
            .I3(GND_net), .O(n32726));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1518.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4490));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22_3_lut_adj_1519 (.I0(bit_ctr[27]), .I1(n39088), .I2(n17536), 
            .I3(GND_net), .O(n32732));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1519.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33177_4_lut (.I0(n31_adj_4490), .I1(n19_adj_4483), .I2(n17_adj_4482), 
            .I3(n15_adj_4480), .O(n39499));
    defparam i33177_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i22_3_lut_adj_1520 (.I0(bit_ctr[26]), .I1(n39087), .I2(n17536), 
            .I3(GND_net), .O(n32730));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1520.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_7 (.CI(n28377), .I0(GND_net), .I1(n20_adj_4194), 
            .CO(n28378));
    SB_LUT4 i13964_3_lut (.I0(encoder0_position[21]), .I1(n2734), .I2(count_enable), 
            .I3(GND_net), .O(n18471));   // quad.v(35[10] 41[6])
    defparam i13964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13963_3_lut (.I0(encoder0_position[20]), .I1(n2735), .I2(count_enable), 
            .I3(GND_net), .O(n18470));   // quad.v(35[10] 41[6])
    defparam i13963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33800_4_lut (.I0(n13_adj_4478), .I1(n11_adj_4476), .I2(n2637), 
            .I3(n98), .O(n40122));
    defparam i33800_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34075_4_lut (.I0(n19_adj_4483), .I1(n17_adj_4482), .I2(n15_adj_4480), 
            .I3(n40122), .O(n40397));
    defparam i34075_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_555_22_lut (.I0(duty[20]), .I1(n41708), .I2(n5), .I3(n27587), 
            .O(pwm_setpoint_22__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_1854_7 (.CI(n28170), .I0(n2753_adj_4081), 
            .I1(VCC_net), .CO(n28171));
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13962_3_lut (.I0(encoder0_position[19]), .I1(n2736), .I2(count_enable), 
            .I3(GND_net), .O(n18469));   // quad.v(35[10] 41[6])
    defparam i13962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4195), .I3(n28376), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_6_lut (.I0(GND_net), .I1(n2754_adj_4080), 
            .I2(GND_net), .I3(n28169), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_6 (.CI(n28376), .I0(GND_net), .I1(n21_adj_4195), 
            .CO(n28377));
    SB_LUT4 i13961_3_lut (.I0(encoder0_position[18]), .I1(n2737), .I2(count_enable), 
            .I3(GND_net), .O(n18468));   // quad.v(35[10] 41[6])
    defparam i13961_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1988_23 (.CI(n28050), .I0(n2937), 
            .I1(VCC_net), .CO(n28051));
    SB_CARRY add_555_22 (.CI(n27587), .I0(n41708), .I1(n5), .CO(n27588));
    SB_LUT4 i13960_3_lut (.I0(encoder0_position[17]), .I1(n2738), .I2(count_enable), 
            .I3(GND_net), .O(n18467));   // quad.v(35[10] 41[6])
    defparam i13960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1988_22_lut (.I0(GND_net), .I1(n2938), 
            .I2(VCC_net), .I3(n28049), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34071_4_lut (.I0(n25_adj_4487), .I1(n23_adj_4486), .I2(n21_adj_4485), 
            .I3(n40397), .O(n40393));
    defparam i34071_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33179_4_lut (.I0(n31_adj_4490), .I1(n29_adj_4489), .I2(n27_adj_4488), 
            .I3(n40393), .O(n39501));
    defparam i33179_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY communication_counter_31__I_0_add_1854_6 (.CI(n28169), .I0(n2754_adj_4080), 
            .I1(GND_net), .CO(n28170));
    SB_CARRY communication_counter_31__I_0_add_1988_22 (.CI(n28049), .I0(n2938), 
            .I1(VCC_net), .CO(n28050));
    SB_LUT4 communication_counter_31__I_0_add_1988_21_lut (.I0(GND_net), .I1(n2939), 
            .I2(VCC_net), .I3(n28048), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_21_lut (.I0(duty[19]), .I1(n41708), .I2(n6), .I3(n27586), 
            .O(pwm_setpoint_22__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4196), .I3(n28375), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_5_lut (.I0(GND_net), .I1(n2755_adj_4079), 
            .I2(GND_net), .I3(n28168), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13959_3_lut (.I0(encoder0_position[16]), .I1(n2739), .I2(count_enable), 
            .I3(GND_net), .O(n18466));   // quad.v(35[10] 41[6])
    defparam i13959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4474));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY div_46_unary_minus_4_add_3_5 (.CI(n28375), .I0(GND_net), .I1(n22_adj_4196), 
            .CO(n28376));
    SB_LUT4 i22_3_lut_adj_1521 (.I0(bit_ctr[31]), .I1(n39092), .I2(n17536), 
            .I3(GND_net), .O(n32742));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1521.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4197), .I3(n28374), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_5 (.CI(n28168), .I0(n2755_adj_4079), 
            .I1(GND_net), .CO(n28169));
    SB_CARRY div_46_unary_minus_4_add_3_4 (.CI(n28374), .I0(GND_net), .I1(n23_adj_4197), 
            .CO(n28375));
    SB_LUT4 div_46_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_3999), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1049_3_lut (.I0(n378), .I1(n6721), .I2(n1553), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4198), .I3(n28373), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_21 (.CI(n27586), .I0(n41708), .I1(n6), .CO(n27587));
    SB_LUT4 communication_counter_31__I_0_add_1854_4_lut (.I0(GND_net), .I1(n2756), 
            .I2(VCC_net), .I3(n28167), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34157_3_lut (.I0(n8_adj_4474), .I1(n87), .I2(n31_adj_4490), 
            .I3(GND_net), .O(n40479));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34157_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4439));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1854_4 (.CI(n28167), .I0(n2756), 
            .I1(VCC_net), .CO(n28168));
    SB_LUT4 i34158_3_lut (.I0(n40479), .I1(n86), .I2(n33_adj_4491), .I3(GND_net), 
            .O(n40480));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34158_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i22_3_lut_adj_1522 (.I0(bit_ctr[30]), .I1(n39091), .I2(n17536), 
            .I3(GND_net), .O(n32738));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1522.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1523 (.I0(bit_ctr[29]), .I1(n39090), .I2(n17536), 
            .I3(GND_net), .O(n32736));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1523.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1524 (.I0(bit_ctr[28]), .I1(n39089), .I2(n17536), 
            .I3(GND_net), .O(n32734));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1524.LUT_INIT = 16'hcaca;
    SB_LUT4 i13973_3_lut (.I0(encoder1_position[6]), .I1(n2699), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18480));   // quad.v(35[10] 41[6])
    defparam i13973_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1988_21 (.CI(n28048), .I0(n2939), 
            .I1(VCC_net), .CO(n28049));
    SB_LUT4 communication_counter_31__I_0_add_1988_20_lut (.I0(GND_net), .I1(n2940), 
            .I2(VCC_net), .I3(n28047), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_20 (.CI(n28047), .I0(n2940), 
            .I1(VCC_net), .CO(n28048));
    SB_CARRY div_46_unary_minus_4_add_3_3 (.CI(n28373), .I0(GND_net), .I1(n24_adj_4198), 
            .CO(n28374));
    SB_LUT4 div_46_LessThan_1722_i34_3_lut (.I0(n16_adj_4481), .I1(n83), 
            .I2(n39_adj_4495), .I3(GND_net), .O(n34_adj_4492));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33173_4_lut (.I0(n37_adj_4494), .I1(n35_adj_4493), .I2(n33_adj_4491), 
            .I3(n39499), .O(n39495));
    defparam i33173_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13972_3_lut (.I0(encoder1_position[5]), .I1(n2700), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18479));   // quad.v(35[10] 41[6])
    defparam i13972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13971_3_lut (.I0(encoder1_position[4]), .I1(n2701), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18478));   // quad.v(35[10] 41[6])
    defparam i13971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34516_4_lut (.I0(n34_adj_4492), .I1(n14_adj_4479), .I2(n39_adj_4495), 
            .I3(n39491), .O(n40838));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34516_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4199), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33671_3_lut (.I0(n40480), .I1(n85), .I2(n35_adj_4493), .I3(GND_net), 
            .O(n39993));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33671_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13970_3_lut (.I0(encoder1_position[3]), .I1(n2702), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18477));   // quad.v(35[10] 41[6])
    defparam i13970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1988_19_lut (.I0(GND_net), .I1(n2941), 
            .I2(VCC_net), .I3(n28046), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_20_lut (.I0(duty[18]), .I1(n41708), .I2(n7_adj_3931), 
            .I3(n27585), .O(pwm_setpoint_22__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13969_3_lut (.I0(encoder1_position[2]), .I1(n2703), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18476));   // quad.v(35[10] 41[6])
    defparam i13969_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1988_19 (.CI(n28046), .I0(n2941), 
            .I1(VCC_net), .CO(n28047));
    SB_LUT4 communication_counter_31__I_0_add_1988_18_lut (.I0(GND_net), .I1(n2942), 
            .I2(VCC_net), .I3(n28045), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_18 (.CI(n28045), .I0(n2942), 
            .I1(VCC_net), .CO(n28046));
    SB_LUT4 communication_counter_31__I_0_add_1988_17_lut (.I0(GND_net), .I1(n2943), 
            .I2(VCC_net), .I3(n28044), .O(n3010)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_17 (.CI(n28044), .I0(n2943), 
            .I1(VCC_net), .CO(n28045));
    SB_LUT4 communication_counter_31__I_0_add_1988_16_lut (.I0(GND_net), .I1(n2944), 
            .I2(VCC_net), .I3(n28043), .O(n3011)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34159_3_lut (.I0(n10_adj_4475), .I1(n90), .I2(n25_adj_4487), 
            .I3(GND_net), .O(n40481));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34159_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_add_1854_3_lut (.I0(GND_net), .I1(n2757), 
            .I2(VCC_net), .I3(n28166), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_3 (.CI(n28166), .I0(n2757), 
            .I1(VCC_net), .CO(n28167));
    SB_LUT4 i13968_3_lut (.I0(encoder1_position[1]), .I1(n2704), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18475));   // quad.v(35[10] 41[6])
    defparam i13968_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1988_16 (.CI(n28043), .I0(n2944), 
            .I1(VCC_net), .CO(n28044));
    SB_LUT4 communication_counter_31__I_0_add_1988_15_lut (.I0(GND_net), .I1(n2945), 
            .I2(VCC_net), .I3(n28042), .O(n3012)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4199), 
            .CO(n28373));
    SB_LUT4 i34160_3_lut (.I0(n40481), .I1(n89), .I2(n27_adj_4488), .I3(GND_net), 
            .O(n40482));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34160_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_add_1854_2_lut (.I0(GND_net), .I1(n2758), 
            .I2(GND_net), .I3(VCC_net), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_15 (.CI(n28042), .I0(n2945), 
            .I1(VCC_net), .CO(n28043));
    SB_LUT4 communication_counter_31__I_0_add_1988_14_lut (.I0(GND_net), .I1(n2946), 
            .I2(VCC_net), .I3(n28041), .O(n3013)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_14 (.CI(n28041), .I0(n2946), 
            .I1(VCC_net), .CO(n28042));
    SB_LUT4 communication_counter_31__I_0_add_1519_21_lut (.I0(n2273_adj_4242), 
            .I1(n2240), .I2(VCC_net), .I3(n28372), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33776_4_lut (.I0(n27_adj_4488), .I1(n25_adj_4487), .I2(n23_adj_4486), 
            .I3(n39523), .O(n40098));
    defparam i33776_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 communication_counter_31__I_0_add_1519_20_lut (.I0(GND_net), .I1(n2241), 
            .I2(VCC_net), .I3(n28371), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i20_3_lut (.I0(n12_adj_4477), .I1(n91), 
            .I2(n23_adj_4486), .I3(GND_net), .O(n20_adj_4484));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_add_1988_13_lut (.I0(GND_net), .I1(n2947), 
            .I2(VCC_net), .I3(n28040), .O(n3014)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_2 (.CI(VCC_net), .I0(n2758), 
            .I1(GND_net), .CO(n28166));
    SB_CARRY communication_counter_31__I_0_add_1988_13 (.CI(n28040), .I0(n2947), 
            .I1(VCC_net), .CO(n28041));
    SB_LUT4 i33669_3_lut (.I0(n40482), .I1(n88), .I2(n29_adj_4489), .I3(GND_net), 
            .O(n39991));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33669_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY communication_counter_31__I_0_add_1519_20 (.CI(n28371), .I0(n2241), 
            .I1(VCC_net), .CO(n28372));
    SB_LUT4 communication_counter_31__I_0_add_1988_12_lut (.I0(GND_net), .I1(n2948), 
            .I2(VCC_net), .I3(n28039), .O(n3015)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34304_4_lut (.I0(n37_adj_4494), .I1(n35_adj_4493), .I2(n33_adj_4491), 
            .I3(n39501), .O(n40626));
    defparam i34304_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_add_1519_19_lut (.I0(GND_net), .I1(n2242), 
            .I2(VCC_net), .I3(n28370), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_12 (.CI(n28039), .I0(n2948), 
            .I1(VCC_net), .CO(n28040));
    SB_LUT4 communication_counter_31__I_0_add_1921_26_lut (.I0(n2867), .I1(n2834), 
            .I2(VCC_net), .I3(n28165), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_1988_11_lut (.I0(GND_net), .I1(n2949), 
            .I2(VCC_net), .I3(n28038), .O(n3016)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34617_4_lut (.I0(n39993), .I1(n40838), .I2(n39_adj_4495), 
            .I3(n39495), .O(n40939));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34617_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 communication_counter_31__I_0_add_1921_25_lut (.I0(GND_net), .I1(n2835), 
            .I2(VCC_net), .I3(n28164), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_19 (.CI(n28370), .I0(n2242), 
            .I1(VCC_net), .CO(n28371));
    SB_LUT4 communication_counter_31__I_0_add_1519_18_lut (.I0(GND_net), .I1(n2243), 
            .I2(VCC_net), .I3(n28369), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_18 (.CI(n28369), .I0(n2243), 
            .I1(VCC_net), .CO(n28370));
    SB_CARRY communication_counter_31__I_0_add_1921_25 (.CI(n28164), .I0(n2835), 
            .I1(VCC_net), .CO(n28165));
    SB_LUT4 i34021_4_lut (.I0(n39991), .I1(n20_adj_4484), .I2(n29_adj_4489), 
            .I3(n40098), .O(n40343));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34021_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 communication_counter_31__I_0_add_1921_24_lut (.I0(GND_net), .I1(n2836), 
            .I2(VCC_net), .I3(n28163), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_11 (.CI(n28038), .I0(n2949), 
            .I1(VCC_net), .CO(n28039));
    SB_LUT4 i34640_4_lut (.I0(n40343), .I1(n40939), .I2(n39_adj_4495), 
            .I3(n40626), .O(n40962));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34640_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY communication_counter_31__I_0_add_1921_24 (.CI(n28163), .I0(n2836), 
            .I1(VCC_net), .CO(n28164));
    SB_LUT4 i34641_3_lut (.I0(n40962), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n40963));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34641_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 communication_counter_31__I_0_add_1988_10_lut (.I0(GND_net), .I1(n2950), 
            .I2(VCC_net), .I3(n28037), .O(n3017)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1519_17_lut (.I0(GND_net), .I1(n2244), 
            .I2(VCC_net), .I3(n28368), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_10 (.CI(n28037), .I0(n2950), 
            .I1(VCC_net), .CO(n28038));
    SB_LUT4 communication_counter_31__I_0_add_1988_9_lut (.I0(GND_net), .I1(n2951), 
            .I2(VCC_net), .I3(n28036), .O(n3018)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_9 (.CI(n28036), .I0(n2951), 
            .I1(VCC_net), .CO(n28037));
    SB_LUT4 communication_counter_31__I_0_add_1921_23_lut (.I0(GND_net), .I1(n2837), 
            .I2(VCC_net), .I3(n28162), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34344_3_lut (.I0(n40963), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n40666));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34344_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 communication_counter_31__I_0_add_1988_8_lut (.I0(GND_net), .I1(n2952), 
            .I2(VCC_net), .I3(n28035), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34345_3_lut (.I0(n40666), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n40667));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34345_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY communication_counter_31__I_0_add_1921_23 (.CI(n28162), .I0(n2837), 
            .I1(VCC_net), .CO(n28163));
    SB_LUT4 i1_4_lut (.I0(n40667), .I1(n16508), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_CARRY communication_counter_31__I_0_add_1988_8 (.CI(n28035), .I0(n2952), 
            .I1(VCC_net), .CO(n28036));
    SB_LUT4 i22_3_lut_adj_1525 (.I0(bit_ctr[7]), .I1(n39070), .I2(n17536), 
            .I3(GND_net), .O(n32692));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1525.LUT_INIT = 16'hcaca;
    SB_LUT4 i13493_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n37153), .I3(GND_net), .O(n18000));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1988_7_lut (.I0(GND_net), .I1(n2953), 
            .I2(VCC_net), .I3(n28034), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_17 (.CI(n28368), .I0(n2244), 
            .I1(VCC_net), .CO(n28369));
    SB_CARRY communication_counter_31__I_0_add_1988_7 (.CI(n28034), .I0(n2953), 
            .I1(VCC_net), .CO(n28035));
    SB_LUT4 communication_counter_31__I_0_add_1519_16_lut (.I0(GND_net), .I1(n2245), 
            .I2(VCC_net), .I3(n28367), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1921_22_lut (.I0(GND_net), .I1(n2838), 
            .I2(VCC_net), .I3(n28161), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY communication_counter_31__I_0_add_1519_16 (.CI(n28367), .I0(n2245), 
            .I1(VCC_net), .CO(n28368));
    SB_LUT4 communication_counter_31__I_0_add_1519_15_lut (.I0(GND_net), .I1(n2246), 
            .I2(VCC_net), .I3(n28366), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1988_6_lut (.I0(GND_net), .I1(n2954), 
            .I2(GND_net), .I3(n28033), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4471));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1921_22 (.CI(n28161), .I0(n2838), 
            .I1(VCC_net), .CO(n28162));
    SB_LUT4 communication_counter_31__I_0_add_1921_21_lut (.I0(GND_net), .I1(n2839), 
            .I2(VCC_net), .I3(n28160), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_15 (.CI(n28366), .I0(n2246), 
            .I1(VCC_net), .CO(n28367));
    SB_LUT4 div_46_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4473));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1519_14_lut (.I0(GND_net), .I1(n2247), 
            .I2(VCC_net), .I3(n28365), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_21 (.CI(n28160), .I0(n2839), 
            .I1(VCC_net), .CO(n28161));
    SB_CARRY communication_counter_31__I_0_add_1988_6 (.CI(n28033), .I0(n2954), 
            .I1(GND_net), .CO(n28034));
    SB_LUT4 div_46_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4469));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1519_14 (.CI(n28365), .I0(n2247), 
            .I1(VCC_net), .CO(n28366));
    SB_LUT4 div_46_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4472));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1988_5_lut (.I0(GND_net), .I1(n2955), 
            .I2(GND_net), .I3(n28032), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_5 (.CI(n28032), .I0(n2955), 
            .I1(GND_net), .CO(n28033));
    SB_LUT4 communication_counter_31__I_0_add_1988_4_lut (.I0(GND_net), .I1(n2956), 
            .I2(VCC_net), .I3(n28031), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_4 (.CI(n28031), .I0(n2956), 
            .I1(VCC_net), .CO(n28032));
    SB_LUT4 communication_counter_31__I_0_add_1988_3_lut (.I0(GND_net), .I1(n2957), 
            .I2(VCC_net), .I3(n28030), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4466));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1921_20_lut (.I0(GND_net), .I1(n2840), 
            .I2(VCC_net), .I3(n28159), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_3 (.CI(n28030), .I0(n2957), 
            .I1(VCC_net), .CO(n28031));
    SB_LUT4 communication_counter_31__I_0_add_1988_2_lut (.I0(GND_net), .I1(n2958), 
            .I2(GND_net), .I3(VCC_net), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1988_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1988_2 (.CI(VCC_net), .I0(n2958), 
            .I1(GND_net), .CO(n28030));
    SB_LUT4 communication_counter_31__I_0_add_1519_13_lut (.I0(GND_net), .I1(n2248), 
            .I2(VCC_net), .I3(n28364), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4467));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4463));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3181_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n28029), 
            .O(n6864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_13 (.CI(n28364), .I0(n2248), 
            .I1(VCC_net), .CO(n28365));
    SB_LUT4 add_3181_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n28028), 
            .O(n6865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_61 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_CARRY add_3181_20 (.CI(n28028), .I0(n2448), .I1(n82), .CO(n28029));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_81[23]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_LUT4 add_3181_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n28027), 
            .O(n6866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4464));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1519_12_lut (.I0(GND_net), .I1(n2249), 
            .I2(VCC_net), .I3(n28363), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_12 (.CI(n28363), .I0(n2249), 
            .I1(VCC_net), .CO(n28364));
    SB_CARRY communication_counter_31__I_0_add_1921_20 (.CI(n28159), .I0(n2840), 
            .I1(VCC_net), .CO(n28160));
    SB_LUT4 div_46_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4465));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1519_11_lut (.I0(GND_net), .I1(n2250), 
            .I2(VCC_net), .I3(n28362), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_11 (.CI(n28362), .I0(n2250), 
            .I1(VCC_net), .CO(n28363));
    SB_CARRY add_3181_19 (.CI(n28027), .I0(n2449), .I1(n83), .CO(n28028));
    SB_LUT4 communication_counter_31__I_0_add_1519_10_lut (.I0(GND_net), .I1(n2251), 
            .I2(VCC_net), .I3(n28361), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1921_19_lut (.I0(GND_net), .I1(n2841), 
            .I2(VCC_net), .I3(n28158), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_10 (.CI(n28361), .I0(n2251), 
            .I1(VCC_net), .CO(n28362));
    SB_LUT4 communication_counter_31__I_0_add_1519_9_lut (.I0(GND_net), .I1(n2252), 
            .I2(VCC_net), .I3(n28360), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4454));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4456));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1519_9 (.CI(n28360), .I0(n2252), 
            .I1(VCC_net), .CO(n28361));
    SB_LUT4 div_46_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4458));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4460));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1519_8_lut (.I0(GND_net), .I1(n2253), 
            .I2(VCC_net), .I3(n28359), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_19 (.CI(n28158), .I0(n2841), 
            .I1(VCC_net), .CO(n28159));
    SB_CARRY communication_counter_31__I_0_add_1519_8 (.CI(n28359), .I0(n2253), 
            .I1(VCC_net), .CO(n28360));
    SB_LUT4 communication_counter_31__I_0_add_1519_7_lut (.I0(GND_net), .I1(n2254), 
            .I2(GND_net), .I3(n28358), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_7 (.CI(n28358), .I0(n2254), 
            .I1(GND_net), .CO(n28359));
    SB_LUT4 communication_counter_31__I_0_add_1519_6_lut (.I0(GND_net), .I1(n2255), 
            .I2(GND_net), .I3(n28357), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1921_18_lut (.I0(GND_net), .I1(n2842), 
            .I2(VCC_net), .I3(n28157), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4461));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4468));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3181_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n28026), 
            .O(n6867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_6 (.CI(n28357), .I0(n2255), 
            .I1(GND_net), .CO(n28358));
    SB_CARRY add_555_20 (.CI(n27585), .I0(n41708), .I1(n7_adj_3931), .CO(n27586));
    SB_LUT4 communication_counter_31__I_0_add_1519_5_lut (.I0(GND_net), .I1(n2256), 
            .I2(VCC_net), .I3(n28356), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_1921_18 (.CI(n28157), .I0(n2842), 
            .I1(VCC_net), .CO(n28158));
    SB_LUT4 i33247_4_lut (.I0(n33_adj_4468), .I1(n21_adj_4461), .I2(n19_adj_4460), 
            .I3(n17_adj_4458), .O(n39569));
    defparam i33247_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33842_4_lut (.I0(n15_adj_4456), .I1(n13_adj_4454), .I2(n2552), 
            .I3(n98), .O(n40164));
    defparam i33842_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY add_3181_18 (.CI(n28026), .I0(n2450), .I1(n84), .CO(n28027));
    SB_LUT4 i34093_4_lut (.I0(n21_adj_4461), .I1(n19_adj_4460), .I2(n17_adj_4458), 
            .I3(n40164), .O(n40415));
    defparam i34093_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34089_4_lut (.I0(n27_adj_4465), .I1(n25_adj_4464), .I2(n23_adj_4463), 
            .I3(n40415), .O(n40411));
    defparam i34089_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY communication_counter_31__I_0_add_1519_5 (.CI(n28356), .I0(n2256), 
            .I1(VCC_net), .CO(n28357));
    SB_LUT4 communication_counter_31__I_0_add_1921_17_lut (.I0(GND_net), .I1(n2843), 
            .I2(VCC_net), .I3(n28156), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1519_4_lut (.I0(GND_net), .I1(n2257), 
            .I2(VCC_net), .I3(n28355), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1519_4 (.CI(n28355), .I0(n2257), 
            .I1(VCC_net), .CO(n28356));
    SB_CARRY communication_counter_31__I_0_add_1921_17 (.CI(n28156), .I0(n2843), 
            .I1(VCC_net), .CO(n28157));
    SB_LUT4 communication_counter_31__I_0_add_1921_16_lut (.I0(GND_net), .I1(n2844), 
            .I2(VCC_net), .I3(n28155), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33249_4_lut (.I0(n33_adj_4468), .I1(n31_adj_4467), .I2(n29_adj_4466), 
            .I3(n40411), .O(n39571));
    defparam i33249_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4452));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34165_3_lut (.I0(n10_adj_4452), .I1(n87), .I2(n33_adj_4468), 
            .I3(GND_net), .O(n40487));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34165_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_add_1519_3_lut (.I0(GND_net), .I1(n2258), 
            .I2(GND_net), .I3(n28354), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34166_3_lut (.I0(n40487), .I1(n86), .I2(n35_adj_4469), .I3(GND_net), 
            .O(n40488));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34166_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i36_3_lut (.I0(n18_adj_4459), .I1(n83), 
            .I2(n41_adj_4473), .I3(GND_net), .O(n36_adj_4470));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33241_4_lut (.I0(n39_adj_4472), .I1(n37_adj_4471), .I2(n35_adj_4469), 
            .I3(n39569), .O(n39563));
    defparam i33241_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34514_4_lut (.I0(n36_adj_4470), .I1(n16_adj_4457), .I2(n41_adj_4473), 
            .I3(n39559), .O(n40836));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34514_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33659_3_lut (.I0(n40488), .I1(n85), .I2(n37_adj_4471), .I3(GND_net), 
            .O(n39981));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33659_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY communication_counter_31__I_0_add_1519_3 (.CI(n28354), .I0(n2258), 
            .I1(GND_net), .CO(n28355));
    SB_CARRY communication_counter_31__I_0_add_1921_16 (.CI(n28155), .I0(n2844), 
            .I1(VCC_net), .CO(n28156));
    SB_LUT4 div_46_i1648_3_lut_3_lut (.I0(n2471), .I1(n6870), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_31__I_0_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4238), 
            .I1(VCC_net), .CO(n28354));
    SB_LUT4 div_46_LessThan_1665_i22_3_lut (.I0(n14_adj_4455), .I1(n91), 
            .I2(n25_adj_4464), .I3(GND_net), .O(n22_adj_4462));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34510_4_lut (.I0(n22_adj_4462), .I1(n12_adj_4453), .I2(n25_adj_4464), 
            .I3(n39630), .O(n40832));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34510_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34511_3_lut (.I0(n40832), .I1(n90), .I2(n27_adj_4465), .I3(GND_net), 
            .O(n40833));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34511_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34391_3_lut (.I0(n40833), .I1(n89), .I2(n29_adj_4466), .I3(GND_net), 
            .O(n40713));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34391_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34310_4_lut (.I0(n39_adj_4472), .I1(n37_adj_4471), .I2(n35_adj_4469), 
            .I3(n39571), .O(n40632));
    defparam i34310_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34615_4_lut (.I0(n39981), .I1(n40836), .I2(n41_adj_4473), 
            .I3(n39563), .O(n40937));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34615_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33657_3_lut (.I0(n40713), .I1(n88), .I2(n31_adj_4467), .I3(GND_net), 
            .O(n39979));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33657_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34652_4_lut (.I0(n39979), .I1(n40937), .I2(n41_adj_4473), 
            .I3(n40632), .O(n40974));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34652_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34653_3_lut (.I0(n40974), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n40975));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34653_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34649_3_lut (.I0(n40975), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n40971));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34649_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1526 (.I0(n40971), .I1(n16505), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1526.LUT_INIT = 16'hceef;
    SB_LUT4 i22_3_lut_adj_1527 (.I0(bit_ctr[18]), .I1(n39072), .I2(n17536), 
            .I3(GND_net), .O(n32696));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1527.LUT_INIT = 16'hcaca;
    SB_LUT4 i13496_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4023), 
            .I3(n16429), .O(n18003));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13496_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13485_3_lut (.I0(n17746), .I1(r_Bit_Index[0]), .I2(n17619), 
            .I3(GND_net), .O(n17992));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13485_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 communication_counter_31__I_0_i786_3_lut (.I0(n1153), .I1(n1220), 
            .I2(n1184), .I3(GND_net), .O(n1252));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i787_3_lut (.I0(n1154), .I1(n1221), 
            .I2(n1184), .I3(GND_net), .O(n1253));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i785_3_lut (.I0(n1152), .I1(n1219), 
            .I2(n1184), .I3(GND_net), .O(n1251));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i789_3_lut (.I0(n1156), .I1(n1223), 
            .I2(n1184), .I3(GND_net), .O(n1255));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i788_3_lut (.I0(n1155), .I1(n1222), 
            .I2(n1184), .I3(GND_net), .O(n1254));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i791_3_lut (.I0(n1158), .I1(n1225), 
            .I2(n1184), .I3(GND_net), .O(n1257));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i790_rep_62_3_lut (.I0(n1157), .I1(n1224), 
            .I2(n1184), .I3(GND_net), .O(n1256));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i790_rep_62_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n34616));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1528 (.I0(n1254), .I1(n1250), .I2(n34616), .I3(n1255), 
            .O(n6_adj_4565));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i1_4_lut_adj_1528.LUT_INIT = 16'heccc;
    SB_LUT4 communication_counter_31__I_0_add_1921_15_lut (.I0(GND_net), .I1(n2845), 
            .I2(VCC_net), .I3(n28154), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1645_3_lut_3_lut (.I0(n2471), .I1(n6867), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_555_19_lut (.I0(duty[17]), .I1(n41708), .I2(n8), .I3(n27584), 
            .O(pwm_setpoint_22__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4565), 
            .O(n1283));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14032_4_lut (.I0(n35922), .I1(r_Clock_Count[0]), .I2(n226), 
            .I3(n2346), .O(n18539));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14032_4_lut.LUT_INIT = 16'h4450;
    SB_CARRY communication_counter_31__I_0_add_1921_15 (.CI(n28154), .I0(n2845), 
            .I1(VCC_net), .CO(n28155));
    SB_LUT4 communication_counter_31__I_0_add_1921_14_lut (.I0(GND_net), .I1(n2846), 
            .I2(VCC_net), .I3(n28153), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13482_3_lut (.I0(n17748), .I1(r_Bit_Index_adj_4664[0]), .I2(n17625), 
            .I3(GND_net), .O(n17989));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13482_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i22_3_lut_adj_1529 (.I0(bit_ctr[0]), .I1(n39073), .I2(n17536), 
            .I3(GND_net), .O(n32698));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1529.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1647_3_lut_3_lut (.I0(n2471), .I1(n6869), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13473_4_lut (.I0(n35922), .I1(r_Clock_Count[6]), .I2(n220), 
            .I3(n2346), .O(n17980));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13473_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 div_46_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_3991), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i24_3_lut (.I0(communication_counter[23]), 
            .I1(n10_adj_3975), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1258));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1530 (.I0(bit_ctr[3]), .I1(n39095), .I2(n17536), 
            .I3(GND_net), .O(n32748));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1530.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_81[22]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_LUT4 i22_3_lut_adj_1531 (.I0(bit_ctr[2]), .I1(n39094), .I2(n17536), 
            .I3(GND_net), .O(n32746));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1531.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1532 (.I0(bit_ctr[1]), .I1(n39093), .I2(n17536), 
            .I3(GND_net), .O(n32744));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1532.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1921_14 (.CI(n28153), .I0(n2846), 
            .I1(VCC_net), .CO(n28154));
    SB_LUT4 div_46_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_1921_13_lut (.I0(GND_net), .I1(n2847), 
            .I2(VCC_net), .I3(n28152), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1533 (.I0(bit_ctr[17]), .I1(n39071), .I2(n17536), 
            .I3(GND_net), .O(n32694));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1533.LUT_INIT = 16'hcaca;
    SB_LUT4 i13435_4_lut (.I0(n35922), .I1(r_Clock_Count[4]), .I2(n222), 
            .I3(n2346), .O(n17942));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13435_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 div_46_i1644_3_lut_3_lut (.I0(n2471), .I1(n6866), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_31__I_0_add_1921_13 (.CI(n28152), .I0(n2847), 
            .I1(VCC_net), .CO(n28153));
    SB_LUT4 i13320_4_lut (.I0(n17748), .I1(r_Bit_Index_adj_4664[2]), .I2(n4706), 
            .I3(n17625), .O(n17827));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13320_4_lut.LUT_INIT = 16'h1444;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_81[21]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_81[20]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_81[19]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_81[18]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_81[17]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_LUT4 i13429_4_lut (.I0(n35922), .I1(r_Clock_Count[2]), .I2(n224_adj_4014), 
            .I3(n2346), .O(n17936));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13429_4_lut.LUT_INIT = 16'h4450;
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_81[16]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_81[15]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_81[14]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_81[13]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_81[12]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_81[11]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_81[10]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_81[9]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_81[8]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_81[7]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_81[6]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_81[5]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_81[4]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_81[3]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_81[2]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_81[1]));   // verilog/TinyFPGA_B.v(207[10] 209[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[22]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[21]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[20]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_LUT4 communication_counter_31__I_0_add_1921_12_lut (.I0(GND_net), .I1(n2848), 
            .I2(VCC_net), .I3(n28151), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_12 (.CI(n28151), .I0(n2848), 
            .I1(VCC_net), .CO(n28152));
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[19]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[18]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[17]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[16]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[15]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[14]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[13]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[12]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[11]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[10]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[9]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[8]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[7]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[6]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[5]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[4]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[3]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_LUT4 i13862_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n33775), .I3(GND_net), .O(n18369));   // verilog/coms.v(126[12] 289[6])
    defparam i13862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13988_3_lut (.I0(encoder1_position[21]), .I1(n2684), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18495));   // quad.v(35[10] 41[6])
    defparam i13988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13987_3_lut (.I0(encoder1_position[20]), .I1(n2685), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n18494));   // quad.v(35[10] 41[6])
    defparam i13987_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[2]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[1]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_DFF communication_counter_1136__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_LUT4 div_46_i1124_3_lut (.I0(n1653), .I1(n6734), .I2(n1667), .I3(GND_net), 
            .O(n1764));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1197_3_lut (.I0(n1764), .I1(n6748), .I2(n1778), .I3(GND_net), 
            .O(n1872));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1268_3_lut (.I0(n1872), .I1(n6763), .I2(n1886), .I3(GND_net), 
            .O(n1977));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1337_3_lut (.I0(n1977), .I1(n6779), .I2(n1991), .I3(GND_net), 
            .O(n2079));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1337_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1404_3_lut (.I0(n2079), .I1(n6796), .I2(n2093), .I3(GND_net), 
            .O(n2178));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1469_3_lut (.I0(n2178), .I1(n6814), .I2(n2192), .I3(GND_net), 
            .O(n2274));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1469_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1532_3_lut (.I0(n2274), .I1(n6833), .I2(n2288), .I3(GND_net), 
            .O(n2367));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1532_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13424_4_lut (.I0(n35922), .I1(r_Clock_Count[1]), .I2(n225), 
            .I3(n2346), .O(n17931));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13424_4_lut.LUT_INIT = 16'h4450;
    SB_LUT4 div_46_i1593_3_lut (.I0(n2367), .I1(n6853), .I2(n2381), .I3(GND_net), 
            .O(n2457));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4442));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_3993), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1475_3_lut (.I0(n384), .I1(n6820), .I2(n2192), .I3(GND_net), 
            .O(n2280));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1538_3_lut (.I0(n2280), .I1(n6839), .I2(n2288), .I3(GND_net), 
            .O(n2373));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13863_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n33775), .I3(GND_net), .O(n18370));   // verilog/coms.v(126[12] 289[6])
    defparam i13863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1534 (.I0(bit_ctr[11]), .I1(n39074), .I2(n17536), 
            .I3(GND_net), .O(n32700));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1534.LUT_INIT = 16'hcaca;
    SB_LUT4 i13864_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n33775), .I3(GND_net), .O(n18371));   // verilog/coms.v(126[12] 289[6])
    defparam i13864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1535 (.I0(bit_ctr[12]), .I1(n39075), .I2(n17536), 
            .I3(GND_net), .O(n32702));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1535.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1643_3_lut_3_lut (.I0(n2471), .I1(n6865), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1649_3_lut_3_lut (.I0(n2471), .I1(n6871), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13865_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n33775), .I3(GND_net), .O(n18372));   // verilog/coms.v(126[12] 289[6])
    defparam i13865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1646_3_lut_3_lut (.I0(n2471), .I1(n6868), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14003_3_lut (.I0(quadA_debounced_adj_4009), .I1(reg_B_adj_4672[1]), 
            .I2(n34961), .I3(GND_net), .O(n18510));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1259_3_lut (.I0(n1863), .I1(n6754), .I2(n1886), .I3(GND_net), 
            .O(n1968));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1328_3_lut (.I0(n1968), .I1(n6770), .I2(n1991), .I3(GND_net), 
            .O(n2070));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1395_3_lut (.I0(n2070), .I1(n6787), .I2(n2093), .I3(GND_net), 
            .O(n2169));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1460_3_lut (.I0(n2169), .I1(n6805), .I2(n2192), .I3(GND_net), 
            .O(n2265));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1921_11_lut (.I0(GND_net), .I1(n2849), 
            .I2(VCC_net), .I3(n28150), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_19 (.CI(n27584), .I0(n41708), .I1(n8), .CO(n27585));
    SB_LUT4 div_46_i1642_3_lut_3_lut (.I0(n2471), .I1(n6864), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_31__I_0_add_1921_11 (.CI(n28150), .I0(n2849), 
            .I1(VCC_net), .CO(n28151));
    SB_LUT4 communication_counter_31__I_0_add_1921_10_lut (.I0(GND_net), .I1(n2850), 
            .I2(VCC_net), .I3(n28149), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1536 (.I0(bit_ctr[13]), .I1(n39076), .I2(n17536), 
            .I3(GND_net), .O(n32708));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1536.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1537 (.I0(bit_ctr[19]), .I1(n39077), .I2(n17536), 
            .I3(GND_net), .O(n32710));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1537.LUT_INIT = 16'hcaca;
    SB_LUT4 i13516_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n37153), .I3(GND_net), .O(n18023));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13516_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_1921_10 (.CI(n28149), .I0(n2850), 
            .I1(VCC_net), .CO(n28150));
    SB_LUT4 i21_3_lut_adj_1538 (.I0(bit_ctr[14]), .I1(n39064), .I2(n17536), 
            .I3(GND_net), .O(n32680));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21_3_lut_adj_1538.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_3_lut_adj_1539 (.I0(bit_ctr[15]), .I1(n39068), .I2(n17536), 
            .I3(GND_net), .O(n32688));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21_3_lut_adj_1539.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1921_9_lut (.I0(GND_net), .I1(n2851), 
            .I2(VCC_net), .I3(n28148), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_18_lut (.I0(duty[16]), .I1(n41708), .I2(n9), .I3(n27583), 
            .O(pwm_setpoint_22__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14011_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1035), .I3(GND_net), .O(n18518));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14010_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1035), .I3(GND_net), .O(n18517));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14010_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1921_9 (.CI(n28148), .I0(n2851), 
            .I1(VCC_net), .CO(n28149));
    SB_LUT4 i14008_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1035), .I3(GND_net), .O(n18515));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1921_8_lut (.I0(GND_net), .I1(n2852), 
            .I2(VCC_net), .I3(n28147), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14007_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1035), .I3(GND_net), .O(n18514));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13517_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n37153), .I3(GND_net), .O(n18024));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13518_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n37153), .I3(GND_net), .O(n18025));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13518_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_1921_8 (.CI(n28147), .I0(n2852), 
            .I1(VCC_net), .CO(n28148));
    SB_LUT4 i13519_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n37153), .I3(GND_net), .O(n18026));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13520_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n37153), .I3(GND_net), .O(n18027));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13521_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n37153), .I3(GND_net), .O(n18028));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1921_7_lut (.I0(GND_net), .I1(n2853), 
            .I2(VCC_net), .I3(n28146), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14006_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1035), .I3(GND_net), .O(n18513));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13522_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n37153), .I3(GND_net), .O(n18029));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_555_18 (.CI(n27583), .I0(n41708), .I1(n9), .CO(n27584));
    SB_LUT4 mux_78_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[7]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_107[7]), 
            .I2(n15), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_555_17_lut (.I0(duty[15]), .I1(n41708), .I2(n10), .I3(n27582), 
            .O(pwm_setpoint_22__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13523_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n37153), .I3(GND_net), .O(n18030));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13524_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n37153), .I3(GND_net), .O(n18031));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13524_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_1921_7 (.CI(n28146), .I0(n2853), 
            .I1(VCC_net), .CO(n28147));
    SB_LUT4 i13525_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n37153), .I3(GND_net), .O(n18032));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13526_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n37153), .I3(GND_net), .O(n18033));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13527_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n37153), .I3(GND_net), .O(n18034));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1921_6_lut (.I0(GND_net), .I1(n2854), 
            .I2(GND_net), .I3(n28145), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3181_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n28025), 
            .O(n6868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_6 (.CI(n28145), .I0(n2854), 
            .I1(GND_net), .CO(n28146));
    SB_LUT4 i13528_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n37153), .I3(GND_net), .O(n18035));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13528_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3181_17 (.CI(n28025), .I0(n2451), .I1(n85), .CO(n28026));
    SB_LUT4 div_46_i1523_3_lut (.I0(n2265), .I1(n6824), .I2(n2288), .I3(GND_net), 
            .O(n2358));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1584_3_lut (.I0(n2358), .I1(n6844), .I2(n2381), .I3(GND_net), 
            .O(n2448));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4003), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i725_3_lut (.I0(n374), .I1(n6675), .I2(n1067), .I3(GND_net), 
            .O(n1175));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i808_3_lut (.I0(n1175), .I1(n6684), .I2(n1193), .I3(GND_net), 
            .O(n1298));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i889_3_lut (.I0(n1298), .I1(n6694), .I2(n1316), .I3(GND_net), 
            .O(n1418));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i968_3_lut (.I0(n1418), .I1(n6705), .I2(n1436), .I3(GND_net), 
            .O(n1535));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1045_3_lut (.I0(n1535), .I1(n6717), .I2(n1553), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1120_3_lut (.I0(n1649), .I1(n6730), .I2(n1667), .I3(GND_net), 
            .O(n1760));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1193_3_lut (.I0(n1760), .I1(n6744), .I2(n1778), .I3(GND_net), 
            .O(n1868));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1264_3_lut (.I0(n1868), .I1(n6759), .I2(n1886), .I3(GND_net), 
            .O(n1973));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1921_5_lut (.I0(GND_net), .I1(n2855), 
            .I2(GND_net), .I3(n28144), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_5 (.CI(n28144), .I0(n2855), 
            .I1(GND_net), .CO(n28145));
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13529_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n37153), .I3(GND_net), .O(n18036));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3181_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n28024), 
            .O(n6869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_16_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1599_3_lut (.I0(n2373), .I1(n6859), .I2(n2381), .I3(GND_net), 
            .O(n2463));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1599_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4432));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_3994), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1409_3_lut (.I0(n383), .I1(n6801), .I2(n2093), .I3(GND_net), 
            .O(n2183));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1474_3_lut (.I0(n2183), .I1(n6819), .I2(n2192), .I3(GND_net), 
            .O(n2279));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1537_3_lut (.I0(n2279), .I1(n6838), .I2(n2288), .I3(GND_net), 
            .O(n2372));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1598_3_lut (.I0(n2372), .I1(n6858), .I2(n2381), .I3(GND_net), 
            .O(n2462));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1598_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4434));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_3998), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1125_3_lut (.I0(n379), .I1(n6735), .I2(n1667), .I3(GND_net), 
            .O(n1765));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1198_3_lut (.I0(n1765), .I1(n6749), .I2(n1778), .I3(GND_net), 
            .O(n1873));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1269_3_lut (.I0(n1873), .I1(n6764), .I2(n1886), .I3(GND_net), 
            .O(n1978));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1338_3_lut (.I0(n1978), .I1(n6780), .I2(n1991), .I3(GND_net), 
            .O(n2080));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1405_3_lut (.I0(n2080), .I1(n6797), .I2(n2093), .I3(GND_net), 
            .O(n2179));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1405_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3181_16 (.CI(n28024), .I0(n2452), .I1(n86), .CO(n28025));
    SB_LUT4 i13530_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n37153), .I3(GND_net), .O(n18037));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13530_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3181_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n28023), 
            .O(n6870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_15 (.CI(n28023), .I0(n2453), .I1(n87), .CO(n28024));
    SB_LUT4 add_3181_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n28022), 
            .O(n6871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_14 (.CI(n28022), .I0(n2454), .I1(n88), .CO(n28023));
    SB_LUT4 add_3181_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n28021), 
            .O(n6872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13531_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n37153), .I3(GND_net), .O(n18038));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13531_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3181_13 (.CI(n28021), .I0(n2455), .I1(n89), .CO(n28022));
    SB_LUT4 add_3181_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n28020), 
            .O(n6873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_12 (.CI(n28020), .I0(n2456), .I1(n90), .CO(n28021));
    SB_LUT4 div_46_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1652_3_lut (.I0(n2457), .I1(n6874), .I2(n2471), .I3(GND_net), 
            .O(n2544));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1921_4_lut (.I0(GND_net), .I1(n2856), 
            .I2(VCC_net), .I3(n28143), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13532_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n37153), .I3(GND_net), .O(n18039));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13532_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_1921_4 (.CI(n28143), .I0(n2856), 
            .I1(VCC_net), .CO(n28144));
    SB_LUT4 i1_4_lut_adj_1540 (.I0(n5_adj_4077), .I1(n123), .I2(n33787), 
            .I3(n63_adj_4076), .O(n6_adj_4008));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1540.LUT_INIT = 16'haeaa;
    SB_LUT4 add_3181_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n28019), 
            .O(n6874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_11 (.CI(n28019), .I0(n2457), .I1(n91), .CO(n28020));
    SB_CARRY add_555_17 (.CI(n27582), .I0(n41708), .I1(n10), .CO(n27583));
    SB_LUT4 communication_counter_31__I_0_add_1921_3_lut (.I0(GND_net), .I1(n2857_adj_4078), 
            .I2(VCC_net), .I3(n28142), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3181_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n28018), 
            .O(n6875)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_648_8_lut (.I0(n986), .I1(n953), 
            .I2(VCC_net), .I3(n28574), .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_648_7_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(n28573), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1921_3 (.CI(n28142), .I0(n2857_adj_4078), 
            .I1(VCC_net), .CO(n28143));
    SB_CARRY add_3181_10 (.CI(n28018), .I0(n2458), .I1(n92), .CO(n28019));
    SB_LUT4 add_3181_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n28017), 
            .O(n6876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_9 (.CI(n28017), .I0(n2459), .I1(n93), .CO(n28018));
    SB_LUT4 add_3181_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n28016), 
            .O(n6877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_8 (.CI(n28016), .I0(n2460), .I1(n94), .CO(n28017));
    SB_LUT4 add_3181_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n28015), 
            .O(n6878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4185));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_1921_2_lut (.I0(GND_net), .I1(n2858), 
            .I2(GND_net), .I3(VCC_net), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1921_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_16_lut (.I0(duty[14]), .I1(n41708), .I2(n11), .I3(n27581), 
            .O(pwm_setpoint_22__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3181_7 (.CI(n28015), .I0(n2461), .I1(n95), .CO(n28016));
    SB_CARRY communication_counter_31__I_0_add_1921_2 (.CI(VCC_net), .I0(n2858), 
            .I1(GND_net), .CO(n28142));
    SB_CARRY communication_counter_31__I_0_add_648_7 (.CI(n28573), .I0(n954), 
            .I1(GND_net), .CO(n28574));
    SB_LUT4 communication_counter_31__I_0_add_648_6_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(n28572), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_648_6 (.CI(n28572), .I0(n955), 
            .I1(GND_net), .CO(n28573));
    SB_LUT4 add_3181_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n28014), 
            .O(n6879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_6 (.CI(n28014), .I0(n2462), .I1(n96), .CO(n28015));
    SB_LUT4 add_3185_25_lut (.I0(n249), .I1(n41713), .I2(n248), .I3(n28141), 
            .O(displacement_23__N_205[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3185_24_lut (.I0(n393), .I1(n41713), .I2(n392), .I3(n28140), 
            .O(displacement_23__N_205[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 communication_counter_31__I_0_add_648_5_lut (.I0(GND_net), .I1(n956), 
            .I2(VCC_net), .I3(n28571), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_24 (.CI(n28140), .I0(n41713), .I1(n392), .CO(n28141));
    SB_LUT4 add_3185_23_lut (.I0(n534), .I1(n41713), .I2(n533), .I3(n28139), 
            .O(displacement_23__N_205[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1333_3_lut (.I0(n1973), .I1(n6775), .I2(n1991), .I3(GND_net), 
            .O(n2075));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1333_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3181_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n28013), 
            .O(n6880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_648_5 (.CI(n28571), .I0(n956), 
            .I1(VCC_net), .CO(n28572));
    SB_LUT4 i13533_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n37153), .I3(GND_net), .O(n18040));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13534_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n37153), .I3(GND_net), .O(n18041));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13534_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3181_5 (.CI(n28013), .I0(n2463), .I1(n97), .CO(n28014));
    SB_CARRY add_3185_23 (.CI(n28139), .I0(n41713), .I1(n533), .CO(n28140));
    SB_LUT4 communication_counter_31__I_0_add_648_4_lut (.I0(GND_net), .I1(n957), 
            .I2(VCC_net), .I3(n28570), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13535_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n37153), .I3(GND_net), .O(n18042));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3185_22_lut (.I0(n672), .I1(n41713), .I2(n671), .I3(n28138), 
            .O(displacement_23__N_205[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13536_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n37153), .I3(GND_net), .O(n18043));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3181_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n28012), 
            .O(n6881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_648_4 (.CI(n28570), .I0(n957), 
            .I1(VCC_net), .CO(n28571));
    SB_CARRY add_3181_4 (.CI(n28012), .I0(n2464), .I1(n98), .CO(n28013));
    SB_LUT4 i13537_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n37153), .I3(GND_net), .O(n18044));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13537_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13538_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n37153), .I3(GND_net), .O(n18045));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13538_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13539_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n37153), .I3(GND_net), .O(n18046));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13539_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1541 (.I0(n16405), .I1(n63_adj_4076), .I2(n9783), 
            .I3(n19_adj_4616), .O(n5_adj_4620));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1541.LUT_INIT = 16'hdc50;
    SB_LUT4 add_3181_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n28011), 
            .O(n6882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_22 (.CI(n28138), .I0(n41713), .I1(n671), .CO(n28139));
    SB_CARRY add_3181_3 (.CI(n28011), .I0(n2465), .I1(n99), .CO(n28012));
    SB_LUT4 add_3181_2_lut (.I0(GND_net), .I1(n387), .I2(n558), .I3(VCC_net), 
            .O(n6883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3181_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3181_2 (.CI(VCC_net), .I0(n387), .I1(n558), .CO(n28011));
    SB_LUT4 i13540_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n37153), .I3(GND_net), .O(n18047));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13540_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3180_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n28010), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3185_21_lut (.I0(n807), .I1(n41713), .I2(n806), .I3(n28137), 
            .O(displacement_23__N_205[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3180_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n28009), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_19 (.CI(n28009), .I0(n2358), .I1(n83), .CO(n28010));
    SB_LUT4 add_3180_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n28008), 
            .O(n6845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_21 (.CI(n28137), .I0(n41713), .I1(n806), .CO(n28138));
    SB_CARRY add_3180_18 (.CI(n28008), .I0(n2359), .I1(n84), .CO(n28009));
    SB_CARRY add_555_16 (.CI(n27581), .I0(n41708), .I1(n11), .CO(n27582));
    SB_LUT4 add_3180_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n28007), 
            .O(n6846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_17 (.CI(n28007), .I0(n2360), .I1(n85), .CO(n28008));
    SB_LUT4 i3_4_lut (.I0(n42588), .I1(n6_adj_4008), .I2(n16420), .I3(n3761), 
            .O(n8_adj_4013));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut.LUT_INIT = 16'hcfce;
    SB_LUT4 add_3185_20_lut (.I0(n939), .I1(n41713), .I2(n938), .I3(n28136), 
            .O(displacement_23__N_205[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 communication_counter_31__I_0_add_648_3_lut (.I0(GND_net), .I1(n958), 
            .I2(GND_net), .I3(n28569), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3180_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n28006), 
            .O(n6847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_16 (.CI(n28006), .I0(n2361), .I1(n86), .CO(n28007));
    SB_LUT4 i13541_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n37153), .I3(GND_net), .O(n18048));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13541_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_648_3 (.CI(n28569), .I0(n958), 
            .I1(GND_net), .CO(n28570));
    SB_CARRY add_3185_20 (.CI(n28136), .I0(n41713), .I1(n938), .CO(n28137));
    SB_LUT4 i13542_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n37153), .I3(GND_net), .O(n18049));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13542_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3180_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n28005), 
            .O(n6848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_15 (.CI(n28005), .I0(n2362), .I1(n87), .CO(n28006));
    SB_LUT4 div_46_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4184));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_648_2 (.CI(VCC_net), .I0(n1058), 
            .I1(VCC_net), .CO(n28569));
    SB_LUT4 communication_counter_31__I_0_add_715_9_lut (.I0(n1085), .I1(n1052), 
            .I2(VCC_net), .I3(n28568), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3185_19_lut (.I0(n1068), .I1(n41713), .I2(n1067), .I3(n28135), 
            .O(displacement_23__N_205[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3180_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n28004), 
            .O(n6849)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_14 (.CI(n28004), .I0(n2363), .I1(n88), .CO(n28005));
    SB_LUT4 communication_counter_31__I_0_add_715_8_lut (.I0(GND_net), .I1(n1053), 
            .I2(VCC_net), .I3(n28567), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_19 (.CI(n28135), .I0(n41713), .I1(n1067), .CO(n28136));
    SB_LUT4 i13543_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n37153), .I3(GND_net), .O(n18050));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13543_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3180_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n28003), 
            .O(n6850)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1542 (.I0(n123), .I1(n8_adj_4013), .I2(n35990), 
            .I3(n5_adj_4620), .O(n41916));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1542.LUT_INIT = 16'hefcf;
    SB_LUT4 div_46_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4450));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_555_15_lut (.I0(duty[13]), .I1(n41708), .I2(n12), .I3(n27580), 
            .O(pwm_setpoint_22__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3180_13 (.CI(n28003), .I0(n2364), .I1(n89), .CO(n28004));
    SB_LUT4 i13544_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n37153), .I3(GND_net), .O(n18051));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13544_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13545_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n37153), .I3(GND_net), .O(n18052));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13545_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13546_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[19] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18053));   // verilog/coms.v(126[12] 289[6])
    defparam i13546_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13547_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[19] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18054));   // verilog/coms.v(126[12] 289[6])
    defparam i13547_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13548_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[19] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18055));   // verilog/coms.v(126[12] 289[6])
    defparam i13548_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1601_3_lut (.I0(n386), .I1(n6861), .I2(n2381), .I3(GND_net), 
            .O(n2465));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13549_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[19] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18056));   // verilog/coms.v(126[12] 289[6])
    defparam i13549_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13550_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[19] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18057));   // verilog/coms.v(126[12] 289[6])
    defparam i13550_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13551_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[19] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18058));   // verilog/coms.v(126[12] 289[6])
    defparam i13551_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13552_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[19] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18059));   // verilog/coms.v(126[12] 289[6])
    defparam i13552_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3180_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n28002), 
            .O(n6851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_12 (.CI(n28002), .I0(n2365), .I1(n90), .CO(n28003));
    SB_LUT4 i13553_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[18] [0]), 
            .I2(n35752), .I3(GND_net), .O(n18060));   // verilog/coms.v(126[12] 289[6])
    defparam i13553_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13554_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[18] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18061));   // verilog/coms.v(126[12] 289[6])
    defparam i13554_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_715_8 (.CI(n28567), .I0(n1053), 
            .I1(VCC_net), .CO(n28568));
    SB_LUT4 communication_counter_31__I_0_add_715_7_lut (.I0(GND_net), .I1(n1054), 
            .I2(GND_net), .I3(n28566), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3185_18_lut (.I0(n1194), .I1(n41713), .I2(n1193), .I3(n28134), 
            .O(displacement_23__N_205[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3180_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n28001), 
            .O(n6852)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_715_7 (.CI(n28566), .I0(n1054), 
            .I1(GND_net), .CO(n28567));
    SB_CARRY add_3185_18 (.CI(n28134), .I0(n41713), .I1(n1193), .CO(n28135));
    SB_LUT4 add_3185_17_lut (.I0(n1317), .I1(n41713), .I2(n1316), .I3(n28133), 
            .O(displacement_23__N_205[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13555_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[18] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18062));   // verilog/coms.v(126[12] 289[6])
    defparam i13555_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3185_17 (.CI(n28133), .I0(n41713), .I1(n1316), .CO(n28134));
    SB_LUT4 i13556_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[18] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18063));   // verilog/coms.v(126[12] 289[6])
    defparam i13556_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13557_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[18] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18064));   // verilog/coms.v(126[12] 289[6])
    defparam i13557_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13558_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[18] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18065));   // verilog/coms.v(126[12] 289[6])
    defparam i13558_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13559_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[18] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18066));   // verilog/coms.v(126[12] 289[6])
    defparam i13559_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1713_3_lut_3_lut (.I0(n2558), .I1(n6900), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_555_15 (.CI(n27580), .I0(n41708), .I1(n12), .CO(n27581));
    SB_LUT4 i13560_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[18] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18067));   // verilog/coms.v(126[12] 289[6])
    defparam i13560_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_715_6_lut (.I0(GND_net), .I1(n1055), 
            .I2(GND_net), .I3(n28565), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_715_6 (.CI(n28565), .I0(n1055), 
            .I1(GND_net), .CO(n28566));
    SB_LUT4 add_3185_16_lut (.I0(n1437), .I1(n41713), .I2(n1436), .I3(n28132), 
            .O(displacement_23__N_205[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 communication_counter_31__I_0_add_715_5_lut (.I0(GND_net), .I1(n1056), 
            .I2(VCC_net), .I3(n28564), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13561_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[17] [0]), 
            .I2(n35752), .I3(GND_net), .O(n18068));   // verilog/coms.v(126[12] 289[6])
    defparam i13561_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13562_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[17] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18069));   // verilog/coms.v(126[12] 289[6])
    defparam i13562_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_715_5 (.CI(n28564), .I0(n1056), 
            .I1(VCC_net), .CO(n28565));
    SB_CARRY add_3185_16 (.CI(n28132), .I0(n41713), .I1(n1436), .CO(n28133));
    SB_LUT4 communication_counter_31__I_0_add_715_4_lut (.I0(GND_net), .I1(n1057), 
            .I2(VCC_net), .I3(n28563), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1400_3_lut (.I0(n2075), .I1(n6792), .I2(n2093), .I3(GND_net), 
            .O(n2174));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3185_15_lut (.I0(n1554), .I1(n41713), .I2(n1553), .I3(n28131), 
            .O(displacement_23__N_205[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13563_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[17] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18070));   // verilog/coms.v(126[12] 289[6])
    defparam i13563_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13564_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[17] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18071));   // verilog/coms.v(126[12] 289[6])
    defparam i13564_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13565_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[17] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18072));   // verilog/coms.v(126[12] 289[6])
    defparam i13565_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13566_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[17] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18073));   // verilog/coms.v(126[12] 289[6])
    defparam i13566_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3185_15 (.CI(n28131), .I0(n41713), .I1(n1553), .CO(n28132));
    SB_CARRY communication_counter_31__I_0_add_715_4 (.CI(n28563), .I0(n1057), 
            .I1(VCC_net), .CO(n28564));
    SB_LUT4 div_46_i1699_3_lut_3_lut (.I0(n2558), .I1(n6886), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_add_715_3_lut (.I0(GND_net), .I1(n1058), 
            .I2(GND_net), .I3(n28562), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_11 (.CI(n28001), .I0(n2366), .I1(n91), .CO(n28002));
    SB_LUT4 add_3185_14_lut (.I0(n1668), .I1(n41713), .I2(n1667), .I3(n28130), 
            .O(displacement_23__N_205[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3180_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n28000), 
            .O(n6853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_14 (.CI(n28130), .I0(n41713), .I1(n1667), .CO(n28131));
    SB_LUT4 communication_counter_31__I_0_i723_3_lut (.I0(n1058), .I1(n1125), 
            .I2(n1085), .I3(GND_net), .O(n1157));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i721_3_lut (.I0(n1056), .I1(n1123), 
            .I2(n1085), .I3(GND_net), .O(n1155));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i720_3_lut (.I0(n1055), .I1(n1122), 
            .I2(n1085), .I3(GND_net), .O(n1154));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i719_3_lut (.I0(n1054), .I1(n1121), 
            .I2(n1085), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1801_3_lut (.I0(n2648), .I1(n2715_adj_4107), 
            .I2(n2669), .I3(GND_net), .O(n2747_adj_4087));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1651_3_lut (.I0(n2456), .I1(n6873), .I2(n2471), .I3(GND_net), 
            .O(n2543));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3180_10 (.CI(n28000), .I0(n2367), .I1(n92), .CO(n28001));
    SB_LUT4 communication_counter_31__I_0_i718_3_lut (.I0(n1053), .I1(n1120), 
            .I2(n1085), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3180_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n27999), 
            .O(n6854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i722_rep_63_3_lut (.I0(n1057), .I1(n1124), 
            .I2(n1085), .I3(GND_net), .O(n1156));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i722_rep_63_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n36625));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1543 (.I0(n1154), .I1(n36625), .I2(n1155), .I3(n1157), 
            .O(n34618));
    defparam i1_4_lut_adj_1543.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_1544 (.I0(n34618), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i3_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_CARRY communication_counter_31__I_0_add_715_3 (.CI(n28562), .I0(n1058), 
            .I1(GND_net), .CO(n28563));
    SB_LUT4 communication_counter_31__I_0_mux_3_i25_3_lut (.I0(communication_counter[24]), 
            .I1(n9_adj_3976), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1158));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3185_13_lut (.I0(n1779), .I1(n41713), .I2(n1778), .I3(n28129), 
            .O(displacement_23__N_205[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13567_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[17] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18074));   // verilog/coms.v(126[12] 289[6])
    defparam i13567_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_715_2 (.CI(VCC_net), .I0(n1158), 
            .I1(VCC_net), .CO(n28562));
    SB_LUT4 communication_counter_31__I_0_add_782_10_lut (.I0(n1184), .I1(n1151), 
            .I2(VCC_net), .I3(n28561), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3185_13 (.CI(n28129), .I0(n41713), .I1(n1778), .CO(n28130));
    SB_LUT4 i13568_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[17] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18075));   // verilog/coms.v(126[12] 289[6])
    defparam i13568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1700_3_lut_3_lut (.I0(n2558), .I1(n6887), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_add_782_9_lut (.I0(GND_net), .I1(n1152), 
            .I2(VCC_net), .I3(n28560), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1545 (.I0(bit_ctr[20]), .I1(n39078), .I2(n17536), 
            .I3(GND_net), .O(n32712));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1545.LUT_INIT = 16'hcaca;
    SB_LUT4 i13570_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18077));   // verilog/coms.v(126[12] 289[6])
    defparam i13570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1800_3_lut (.I0(n2647), .I1(n2714_adj_4108), 
            .I2(n2669), .I3(GND_net), .O(n2746_adj_4088));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1800_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF blue_1137__i0 (.Q(blue[0]), .C(LED_c), .D(n45));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_LUT4 add_3185_12_lut (.I0(n1887), .I1(n41713), .I2(n1886), .I3(n28128), 
            .O(displacement_23__N_205[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13571_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18078));   // verilog/coms.v(126[12] 289[6])
    defparam i13571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13572_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18079));   // verilog/coms.v(126[12] 289[6])
    defparam i13572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13573_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18080));   // verilog/coms.v(126[12] 289[6])
    defparam i13573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13574_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18081));   // verilog/coms.v(126[12] 289[6])
    defparam i13574_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3185_12 (.CI(n28128), .I0(n41713), .I1(n1886), .CO(n28129));
    SB_LUT4 div_46_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3180_9 (.CI(n27999), .I0(n2368), .I1(n93), .CO(n28000));
    SB_LUT4 add_3180_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n27998), 
            .O(n6855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_8 (.CI(n27998), .I0(n2369), .I1(n94), .CO(n27999));
    SB_LUT4 add_3180_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n27997), 
            .O(n6856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_3_lut_adj_1546 (.I0(bit_ctr[5]), .I1(n39065), .I2(n17536), 
            .I3(GND_net), .O(n32682));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21_3_lut_adj_1546.LUT_INIT = 16'hcaca;
    SB_LUT4 i13323_4_lut (.I0(n17748), .I1(r_Bit_Index_adj_4664[1]), .I2(r_Bit_Index_adj_4664[0]), 
            .I3(n17625), .O(n17830));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13323_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 add_3185_11_lut (.I0(n1992), .I1(n41713), .I2(n1991), .I3(n28127), 
            .O(displacement_23__N_205[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1470_3_lut (.I0(n2179), .I1(n6815), .I2(n2192), .I3(GND_net), 
            .O(n2275));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_555_14_lut (.I0(duty[12]), .I1(n41708), .I2(n13), .I3(n27579), 
            .O(pwm_setpoint_22__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_782_9 (.CI(n28560), .I0(n1152), 
            .I1(VCC_net), .CO(n28561));
    SB_CARRY add_3185_11 (.CI(n28127), .I0(n41713), .I1(n1991), .CO(n28128));
    SB_LUT4 div_46_i1465_3_lut (.I0(n2174), .I1(n6810), .I2(n2192), .I3(GND_net), 
            .O(n2270));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3185_10_lut (.I0(n2094), .I1(n41713), .I2(n2093), .I3(n28126), 
            .O(displacement_23__N_205[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_555_14 (.CI(n27579), .I0(n41708), .I1(n13), .CO(n27580));
    SB_LUT4 i13326_4_lut (.I0(n17746), .I1(r_Bit_Index[2]), .I2(n4684), 
            .I3(n17619), .O(n17833));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13326_4_lut.LUT_INIT = 16'h1444;
    SB_CARRY add_3180_7 (.CI(n27997), .I0(n2370), .I1(n95), .CO(n27998));
    SB_LUT4 add_3180_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n27996), 
            .O(n6857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4183));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1701_3_lut_3_lut (.I0(n2558), .I1(n6888), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13575_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18082));   // verilog/coms.v(126[12] 289[6])
    defparam i13575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_782_8_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n28559), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13576_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18083));   // verilog/coms.v(126[12] 289[6])
    defparam i13576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13577_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18084));   // verilog/coms.v(126[12] 289[6])
    defparam i13577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13578_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18085));   // verilog/coms.v(126[12] 289[6])
    defparam i13578_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3185_10 (.CI(n28126), .I0(n41713), .I1(n2093), .CO(n28127));
    SB_CARRY add_3180_6 (.CI(n27996), .I0(n2371), .I1(n96), .CO(n27997));
    SB_LUT4 div_46_i1702_3_lut_3_lut (.I0(n2558), .I1(n6889), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13579_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18086));   // verilog/coms.v(126[12] 289[6])
    defparam i13579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13580_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18087));   // verilog/coms.v(126[12] 289[6])
    defparam i13580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13581_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18088));   // verilog/coms.v(126[12] 289[6])
    defparam i13581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13582_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18089));   // verilog/coms.v(126[12] 289[6])
    defparam i13582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13583_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18090));   // verilog/coms.v(126[12] 289[6])
    defparam i13583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13329_4_lut (.I0(n17746), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n17619), .O(n17836));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13329_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i13584_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18091));   // verilog/coms.v(126[12] 289[6])
    defparam i13584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13585_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18092));   // verilog/coms.v(126[12] 289[6])
    defparam i13585_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_782_8 (.CI(n28559), .I0(n1153), 
            .I1(VCC_net), .CO(n28560));
    SB_LUT4 add_3180_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n27995), 
            .O(n6858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13586_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18093));   // verilog/coms.v(126[12] 289[6])
    defparam i13586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13587_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18094));   // verilog/coms.v(126[12] 289[6])
    defparam i13587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13588_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18095));   // verilog/coms.v(126[12] 289[6])
    defparam i13588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_782_7_lut (.I0(GND_net), .I1(n1154), 
            .I2(GND_net), .I3(n28558), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_782_7 (.CI(n28558), .I0(n1154), 
            .I1(GND_net), .CO(n28559));
    SB_LUT4 add_3185_9_lut (.I0(n2193), .I1(n41713), .I2(n2192), .I3(n28125), 
            .O(displacement_23__N_205[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3185_9 (.CI(n28125), .I0(n41713), .I1(n2192), .CO(n28126));
    SB_CARRY add_3180_5 (.CI(n27995), .I0(n2372), .I1(n97), .CO(n27996));
    SB_LUT4 add_3185_8_lut (.I0(n2289), .I1(n41713), .I2(n2288), .I3(n28124), 
            .O(displacement_23__N_205[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 communication_counter_31__I_0_add_782_6_lut (.I0(GND_net), .I1(n1155), 
            .I2(GND_net), .I3(n28557), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_782_6 (.CI(n28557), .I0(n1155), 
            .I1(GND_net), .CO(n28558));
    SB_LUT4 mux_78_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[8]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_107[8]), 
            .I2(n15), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3180_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n27994), 
            .O(n6859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13589_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18096));   // verilog/coms.v(126[12] 289[6])
    defparam i13589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_782_5_lut (.I0(GND_net), .I1(n1156), 
            .I2(VCC_net), .I3(n28556), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_8 (.CI(n28124), .I0(n41713), .I1(n2288), .CO(n28125));
    SB_LUT4 i13590_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18097));   // verilog/coms.v(126[12] 289[6])
    defparam i13590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3185_7_lut (.I0(n2382), .I1(n41713), .I2(n2381), .I3(n28123), 
            .O(displacement_23__N_205[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_782_5 (.CI(n28556), .I0(n1156), 
            .I1(VCC_net), .CO(n28557));
    SB_LUT4 communication_counter_31__I_0_add_782_4_lut (.I0(GND_net), .I1(n1157), 
            .I2(VCC_net), .I3(n28555), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13591_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18098));   // verilog/coms.v(126[12] 289[6])
    defparam i13591_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3180_4 (.CI(n27994), .I0(n2373), .I1(n98), .CO(n27995));
    SB_LUT4 i13592_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18099));   // verilog/coms.v(126[12] 289[6])
    defparam i13592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i744_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_782_4 (.CI(n28555), .I0(n1157), 
            .I1(VCC_net), .CO(n28556));
    SB_LUT4 communication_counter_31__I_0_add_782_3_lut (.I0(GND_net), .I1(n1158), 
            .I2(GND_net), .I3(n28554), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3185_7 (.CI(n28123), .I0(n41713), .I1(n2381), .CO(n28124));
    SB_LUT4 i13593_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18100));   // verilog/coms.v(126[12] 289[6])
    defparam i13593_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_782_3 (.CI(n28554), .I0(n1158), 
            .I1(GND_net), .CO(n28555));
    SB_LUT4 add_3185_6_lut (.I0(n2472), .I1(n41713), .I2(n2471), .I3(n28122), 
            .O(displacement_23__N_205[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3185_6 (.CI(n28122), .I0(n41713), .I1(n2471), .CO(n28123));
    SB_LUT4 div_46_i1533_3_lut (.I0(n2275), .I1(n6834), .I2(n2288), .I3(GND_net), 
            .O(n2368));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1594_3_lut (.I0(n2368), .I1(n6854), .I2(n2381), .I3(GND_net), 
            .O(n2458));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1594_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4441));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4005), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33363_3_lut (.I0(n372), .I1(n558), .I2(n806), .I3(GND_net), 
            .O(n918));
    defparam i33363_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_46_i638_3_lut (.I0(n918), .I1(n6665), .I2(n938), .I3(GND_net), 
            .O(n1047));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i723_3_lut (.I0(n1047), .I1(n6673), .I2(n1067), .I3(GND_net), 
            .O(n1173));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i806_3_lut (.I0(n1173), .I1(n6682), .I2(n1193), .I3(GND_net), 
            .O(n1296));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13594_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18101));   // verilog/coms.v(126[12] 289[6])
    defparam i13594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3180_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n27993), 
            .O(n6860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_3 (.CI(n27993), .I0(n2374), .I1(n99), .CO(n27994));
    SB_LUT4 i13595_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18102));   // verilog/coms.v(126[12] 289[6])
    defparam i13595_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_782_2 (.CI(VCC_net), .I0(n1258), 
            .I1(VCC_net), .CO(n28554));
    SB_LUT4 i13596_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18103));   // verilog/coms.v(126[12] 289[6])
    defparam i13596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3180_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6861)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3180_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3180_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n27993));
    SB_LUT4 add_3179_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n27992), 
            .O(n6823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3179_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n27991), 
            .O(n6824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13597_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18104));   // verilog/coms.v(126[12] 289[6])
    defparam i13597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_849_11_lut (.I0(n1283), .I1(n1250), 
            .I2(VCC_net), .I3(n28553), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3179_18 (.CI(n27991), .I0(n2265), .I1(n84), .CO(n27992));
    SB_LUT4 communication_counter_31__I_0_i651_3_lut (.I0(n954), .I1(n1021), 
            .I2(n986), .I3(GND_net), .O(n1053));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_849_10_lut (.I0(GND_net), .I1(n1251), 
            .I2(VCC_net), .I3(n28552), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3179_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n27990), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i653_3_lut (.I0(n956), .I1(n1023), 
            .I2(n986), .I3(GND_net), .O(n1055));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i652_3_lut (.I0(n955), .I1(n1022), 
            .I2(n986), .I3(GND_net), .O(n1054));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3179_17 (.CI(n27990), .I0(n2266), .I1(n85), .CO(n27991));
    SB_LUT4 communication_counter_31__I_0_i655_3_lut (.I0(n958), .I1(n1025), 
            .I2(n986), .I3(GND_net), .O(n1057));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i654_rep_64_3_lut (.I0(n957), .I1(n1024), 
            .I2(n986), .I3(GND_net), .O(n1056));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i654_rep_64_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1547 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n34622));
    defparam i1_3_lut_adj_1547.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1548 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n36621));
    defparam i1_2_lut_adj_1548.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1549 (.I0(n1052), .I1(n36621), .I2(n1053), .I3(n34622), 
            .O(n1085));
    defparam i1_4_lut_adj_1549.LUT_INIT = 16'hfefa;
    SB_LUT4 communication_counter_31__I_0_mux_3_i26_3_lut (.I0(communication_counter[25]), 
            .I1(n8_adj_3977), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1058));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_849_10 (.CI(n28552), .I0(n1251), 
            .I1(VCC_net), .CO(n28553));
    SB_LUT4 add_3185_5_lut (.I0(n2559), .I1(n41713), .I2(n2558), .I3(n28121), 
            .O(displacement_23__N_205[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_555_13_lut (.I0(duty[11]), .I1(n41708), .I2(n14), .I3(n27578), 
            .O(pwm_setpoint_22__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3185_5 (.CI(n28121), .I0(n41713), .I1(n2558), .CO(n28122));
    SB_LUT4 div_46_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1705_3_lut_3_lut (.I0(n2558), .I1(n6892), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3179_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n27989), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_16 (.CI(n27989), .I0(n2267), .I1(n86), .CO(n27990));
    SB_LUT4 add_3179_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n27988), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_15 (.CI(n27988), .I0(n2268), .I1(n87), .CO(n27989));
    SB_LUT4 div_46_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3179_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n27987), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13598_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18105));   // verilog/coms.v(126[12] 289[6])
    defparam i13598_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3179_14 (.CI(n27987), .I0(n2269), .I1(n88), .CO(n27988));
    SB_LUT4 i13599_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18106));   // verilog/coms.v(126[12] 289[6])
    defparam i13599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13600_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18107));   // verilog/coms.v(126[12] 289[6])
    defparam i13600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3179_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n27986), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_849_9_lut (.I0(GND_net), .I1(n1252), 
            .I2(VCC_net), .I3(n28551), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i887_3_lut (.I0(n1296), .I1(n6692), .I2(n1316), .I3(GND_net), 
            .O(n1416));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13601_3_lut (.I0(Kp[1]), .I1(\data_in_frame[2] [1]), .I2(n35752), 
            .I3(GND_net), .O(n18108));   // verilog/coms.v(126[12] 289[6])
    defparam i13601_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i966_3_lut (.I0(n1416), .I1(n6703), .I2(n1436), .I3(GND_net), 
            .O(n1533));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3185_4_lut (.I0(n2643), .I1(n41713), .I2(n2642), .I3(n28120), 
            .O(displacement_23__N_205[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3185_4 (.CI(n28120), .I0(n41713), .I1(n2642), .CO(n28121));
    SB_CARRY communication_counter_31__I_0_add_849_9 (.CI(n28551), .I0(n1252), 
            .I1(VCC_net), .CO(n28552));
    SB_LUT4 i13602_3_lut (.I0(Kp[2]), .I1(\data_in_frame[2] [2]), .I2(n35752), 
            .I3(GND_net), .O(n18109));   // verilog/coms.v(126[12] 289[6])
    defparam i13602_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13603_3_lut (.I0(Kp[3]), .I1(\data_in_frame[2] [3]), .I2(n35752), 
            .I3(GND_net), .O(n18110));   // verilog/coms.v(126[12] 289[6])
    defparam i13603_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3179_13 (.CI(n27986), .I0(n2270), .I1(n89), .CO(n27987));
    SB_LUT4 add_3179_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n27985), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4001), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i891_3_lut (.I0(n376), .I1(n6696), .I2(n1316), .I3(GND_net), 
            .O(n1420));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i891_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3179_12 (.CI(n27985), .I0(n2271), .I1(n90), .CO(n27986));
    SB_LUT4 div_46_i1528_3_lut (.I0(n2270), .I1(n6829), .I2(n2288), .I3(GND_net), 
            .O(n2363));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1528_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13604_3_lut (.I0(Kp[4]), .I1(\data_in_frame[2] [4]), .I2(n35752), 
            .I3(GND_net), .O(n18111));   // verilog/coms.v(126[12] 289[6])
    defparam i13604_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3179_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n27984), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i970_3_lut (.I0(n1420), .I1(n6707), .I2(n1436), .I3(GND_net), 
            .O(n1537));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1047_3_lut (.I0(n1537), .I1(n6719), .I2(n1553), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3185_3_lut (.I0(n2724), .I1(n41713), .I2(n2723), .I3(n28119), 
            .O(displacement_23__N_205[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n16472), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_CARRY add_555_13 (.CI(n27578), .I0(n41708), .I1(n14), .CO(n27579));
    SB_LUT4 add_7128_7_lut (.I0(n36629), .I1(n746), .I2(GND_net), .I3(n29221), 
            .O(n36236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7128_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3185_3 (.CI(n28119), .I0(n41713), .I1(n2723), .CO(n28120));
    SB_LUT4 add_7128_6_lut (.I0(GND_net), .I1(n852), .I2(GND_net), .I3(n29220), 
            .O(n11515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7128_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_11 (.CI(n27984), .I0(n2272), .I1(n91), .CO(n27985));
    SB_LUT4 add_3179_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n27983), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_10 (.CI(n27983), .I0(n2273), .I1(n92), .CO(n27984));
    SB_LUT4 div_46_i1122_3_lut (.I0(n1651), .I1(n6732), .I2(n1667), .I3(GND_net), 
            .O(n1762));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1195_3_lut (.I0(n1762), .I1(n6746), .I2(n1778), .I3(GND_net), 
            .O(n1870));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1703_3_lut_3_lut (.I0(n2558), .I1(n6890), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35393_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n41713));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i35393_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3185_2_lut (.I0(n2802), .I1(n41713), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_205[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3185_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3179_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n27982), 
            .O(n6833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1266_3_lut (.I0(n1870), .I1(n6761), .I2(n1886), .I3(GND_net), 
            .O(n1975));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1335_3_lut (.I0(n1975), .I1(n6777), .I2(n1991), .I3(GND_net), 
            .O(n2077));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13605_3_lut (.I0(Kp[5]), .I1(\data_in_frame[2] [5]), .I2(n35752), 
            .I3(GND_net), .O(n18112));   // verilog/coms.v(126[12] 289[6])
    defparam i13605_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_7128_6 (.CI(n29220), .I0(n852), .I1(GND_net), .CO(n29221));
    SB_LUT4 add_7128_5_lut (.I0(GND_net), .I1(n748), .I2(VCC_net), .I3(n29219), 
            .O(n11516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7128_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_849_8_lut (.I0(GND_net), .I1(n1253), 
            .I2(VCC_net), .I3(n28550), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_9 (.CI(n27982), .I0(n2274), .I1(n93), .CO(n27983));
    SB_LUT4 div_46_i1402_3_lut (.I0(n2077), .I1(n6794), .I2(n2093), .I3(GND_net), 
            .O(n2176));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1467_3_lut (.I0(n2176), .I1(n6812), .I2(n2192), .I3(GND_net), 
            .O(n2272));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1530_3_lut (.I0(n2272), .I1(n6831), .I2(n2288), .I3(GND_net), 
            .O(n2365));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1530_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_849_8 (.CI(n28550), .I0(n1253), 
            .I1(VCC_net), .CO(n28551));
    SB_LUT4 add_3179_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n27981), 
            .O(n6834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1591_3_lut (.I0(n2365), .I1(n6851), .I2(n2381), .I3(GND_net), 
            .O(n2455));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1650_3_lut (.I0(n2455), .I1(n6872), .I2(n2471), .I3(GND_net), 
            .O(n2542));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_78_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[9]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_107[9]), 
            .I2(n15), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3179_8 (.CI(n27981), .I0(n2275), .I1(n94), .CO(n27982));
    SB_LUT4 mux_78_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[22]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_107[22]), 
            .I2(n15), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3185_2 (.CI(VCC_net), .I0(n41713), .I1(n2801), .CO(n28119));
    SB_LUT4 add_3179_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n27980), 
            .O(n6835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4182));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1799_3_lut (.I0(n2646), .I1(n2713_adj_4109), 
            .I2(n2669), .I3(GND_net), .O(n2745_adj_4089));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4181));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1706_3_lut_3_lut (.I0(n2558), .I1(n6893), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_7128_5 (.CI(n29219), .I0(n748), .I1(VCC_net), .CO(n29220));
    SB_CARRY add_3179_7 (.CI(n27980), .I0(n2276), .I1(n95), .CO(n27981));
    SB_LUT4 add_3179_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n27979), 
            .O(n6836)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4180));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4179));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1798_3_lut (.I0(n2645), .I1(n2712_adj_4110), 
            .I2(n2669), .I3(GND_net), .O(n2744_adj_4090));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4178));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1797_3_lut (.I0(n2644), .I1(n2711_adj_4111), 
            .I2(n2669), .I3(GND_net), .O(n2743_adj_4091));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_849_7_lut (.I0(GND_net), .I1(n1254), 
            .I2(GND_net), .I3(n28549), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_6 (.CI(n27979), .I0(n2277), .I1(n96), .CO(n27980));
    SB_LUT4 div_46_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4177));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4176));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_mux_3_i30_3_lut (.I0(communication_counter[29]), 
            .I1(n4_adj_3981), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n748));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1719_3_lut_3_lut (.I0(n2558), .I1(n6906), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3179_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n27978), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n16421), 
            .I3(GND_net), .O(n15_adj_3943));   // verilog/TinyFPGA_B.v(187[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4_4_lut_adj_1550 (.I0(control_mode[3]), .I1(control_mode[7]), 
            .I2(control_mode[4]), .I3(control_mode[5]), .O(n10_adj_4566));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i4_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[2]), .I1(n10_adj_4566), .I2(control_mode[6]), 
            .I3(GND_net), .O(n16421));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i29_3_lut (.I0(communication_counter[28]), 
            .I1(n5_adj_3980), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n749));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3179_5 (.CI(n27978), .I0(n2278), .I1(n97), .CO(n27979));
    SB_LUT4 mux_78_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[23]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_107[23]), 
            .I2(n15), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1796_3_lut (.I0(n2643_adj_4120), 
            .I1(n2710_adj_4112), .I2(n2669), .I3(GND_net), .O(n2742_adj_4092));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4223));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1795_3_lut (.I0(n2642_adj_4134), 
            .I1(n2709_adj_4113), .I2(n2669), .I3(GND_net), .O(n2741_adj_4093));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3179_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n27977), 
            .O(n6838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4222));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4221));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4220));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1794_3_lut (.I0(n2641), .I1(n2708_adj_4114), 
            .I2(n2669), .I3(GND_net), .O(n2740_adj_4094));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4219));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_3995), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1341_3_lut (.I0(n382), .I1(n6783), .I2(n1991), .I3(GND_net), 
            .O(n2083));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_mux_3_i31_3_lut (.I0(communication_counter[30]), 
            .I1(n3_adj_3982), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n852));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1704_3_lut_3_lut (.I0(n2558), .I1(n6891), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1551 (.I0(n852), .I1(n749), .I2(n748), .I3(n855), 
            .O(n36607));
    defparam i1_4_lut_adj_1551.LUT_INIT = 16'haaa8;
    SB_LUT4 add_7128_4_lut (.I0(GND_net), .I1(n749), .I2(VCC_net), .I3(n29218), 
            .O(n11517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7128_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7128_4 (.CI(n29218), .I0(n749), .I1(VCC_net), .CO(n29219));
    SB_LUT4 add_3184_25_lut (.I0(GND_net), .I1(n2699_adj_4065), .I2(n78), 
            .I3(n28118), .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_849_7 (.CI(n28549), .I0(n1254), 
            .I1(GND_net), .CO(n28550));
    SB_LUT4 add_3184_24_lut (.I0(GND_net), .I1(n2700_adj_4066), .I2(n79), 
            .I3(n28117), .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_mux_3_i28_3_lut (.I0(communication_counter[27]), 
            .I1(n6_adj_3979), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n855));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i27_3_lut (.I0(communication_counter[26]), 
            .I1(n7_adj_3978), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n958));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1708_3_lut_3_lut (.I0(n2558), .I1(n6895), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_7128_3_lut (.I0(GND_net), .I1(n855), .I2(GND_net), .I3(n29217), 
            .O(n11518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7128_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_24 (.CI(n28117), .I0(n2700_adj_4066), .I1(n79), 
            .CO(n28118));
    SB_LUT4 add_555_12_lut (.I0(duty[10]), .I1(n41708), .I2(n15_adj_3932), 
            .I3(n27577), .O(pwm_setpoint_22__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3184_23_lut (.I0(GND_net), .I1(n2701_adj_4067), .I2(n80), 
            .I3(n28116), .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_7128_3 (.CI(n29217), .I0(n855), .I1(GND_net), .CO(n29218));
    SB_LUT4 div_46_i1408_3_lut (.I0(n2083), .I1(n6800), .I2(n2093), .I3(GND_net), 
            .O(n2182));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1709_3_lut_3_lut (.I0(n2558), .I1(n6896), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3184_23 (.CI(n28116), .I0(n2701_adj_4067), .I1(n80), 
            .CO(n28117));
    SB_CARRY add_7128_2 (.CI(VCC_net), .I0(n958), .I1(VCC_net), .CO(n29217));
    SB_LUT4 add_3184_22_lut (.I0(GND_net), .I1(n2702_adj_4068), .I2(n81), 
            .I3(n28115), .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_849_6_lut (.I0(GND_net), .I1(n1255), 
            .I2(GND_net), .I3(n28548), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_849_6 (.CI(n28548), .I0(n1255), 
            .I1(GND_net), .CO(n28549));
    SB_LUT4 blue_1137_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(blue[7]), 
            .I3(n28312), .O(n38_adj_4147)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_22 (.CI(n28115), .I0(n2702_adj_4068), .I1(n81), 
            .CO(n28116));
    SB_LUT4 blue_1137_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(blue[6]), 
            .I3(n28311), .O(n39_adj_4148)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3184_21_lut (.I0(GND_net), .I1(n2703_adj_4069), .I2(n82), 
            .I3(n28114), .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_12 (.CI(n27577), .I0(n41708), .I1(n15_adj_3932), 
            .CO(n27578));
    SB_LUT4 i1_3_lut_adj_1552 (.I0(n956), .I1(n957), .I2(n958), .I3(GND_net), 
            .O(n34624));
    defparam i1_3_lut_adj_1552.LUT_INIT = 16'hfefe;
    SB_CARRY add_3179_4 (.CI(n27977), .I0(n2279), .I1(n98), .CO(n27978));
    SB_CARRY add_3184_21 (.CI(n28114), .I0(n2703_adj_4069), .I1(n82), 
            .CO(n28115));
    SB_LUT4 communication_counter_31__I_0_add_849_5_lut (.I0(GND_net), .I1(n1256), 
            .I2(VCC_net), .I3(n28547), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1137_add_4_8 (.CI(n28311), .I0(GND_net), .I1(blue[6]), 
            .CO(n28312));
    SB_LUT4 add_3184_20_lut (.I0(GND_net), .I1(n2704_adj_4070), .I2(n83), 
            .I3(n28113), .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_11_lut (.I0(duty[9]), .I1(n41708), .I2(n16), .I3(n27576), 
            .O(pwm_setpoint_22__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 blue_1137_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(blue[5]), 
            .I3(n28310), .O(n40_adj_4149)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_20 (.CI(n28113), .I0(n2704_adj_4070), .I1(n83), 
            .CO(n28114));
    SB_LUT4 add_3179_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n27976), 
            .O(n6839)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3179_3 (.CI(n27976), .I0(n2280), .I1(n99), .CO(n27977));
    SB_LUT4 add_3179_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3179_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21074_4_lut (.I0(n954), .I1(n953), .I2(n34624), .I3(n955), 
            .O(n986));
    defparam i21074_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 add_3184_19_lut (.I0(GND_net), .I1(n2705_adj_4071), .I2(n84), 
            .I3(n28112), .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28123_2_lut (.I0(n36236), .I1(n746), .I2(GND_net), .I3(GND_net), 
            .O(n953));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i28123_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_4568), .I3(n29216), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3179_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n27976));
    SB_LUT4 i13606_3_lut (.I0(Kp[6]), .I1(\data_in_frame[2] [6]), .I2(n35752), 
            .I3(GND_net), .O(n18113));   // verilog/coms.v(126[12] 289[6])
    defparam i13606_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY blue_1137_add_4_7 (.CI(n28310), .I0(GND_net), .I1(blue[5]), 
            .CO(n28311));
    SB_CARRY communication_counter_31__I_0_add_849_5 (.CI(n28547), .I0(n1256), 
            .I1(VCC_net), .CO(n28548));
    SB_LUT4 blue_1137_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(blue[4]), 
            .I3(n28309), .O(n41_adj_4150)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1043_3_lut (.I0(n1533), .I1(n6715), .I2(n1553), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_849_4_lut (.I0(GND_net), .I1(n1257), 
            .I2(VCC_net), .I3(n28546), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1473_3_lut (.I0(n2182), .I1(n6818), .I2(n2192), .I3(GND_net), 
            .O(n2278));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1473_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3184_19 (.CI(n28112), .I0(n2705_adj_4071), .I1(n84), 
            .CO(n28113));
    SB_CARRY communication_counter_31__I_0_add_849_4 (.CI(n28546), .I0(n1257), 
            .I1(VCC_net), .CO(n28547));
    SB_LUT4 add_3184_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n28111), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_849_3_lut (.I0(GND_net), .I1(n1258), 
            .I2(GND_net), .I3(n28545), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1137_add_4_6 (.CI(n28309), .I0(GND_net), .I1(blue[4]), 
            .CO(n28310));
    SB_CARRY add_3184_18 (.CI(n28111), .I0(n2706), .I1(n85), .CO(n28112));
    SB_DFF color_16__59 (.Q(color[16]), .C(LED_c), .D(n17951));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_17__58 (.Q(color[17]), .C(LED_c), .D(n17950));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_18__57 (.Q(color[18]), .C(LED_c), .D(n17949));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_23__52 (.Q(color[23]), .C(LED_c), .D(n17948));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_19__56 (.Q(color[19]), .C(LED_c), .D(n17947));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_20__55 (.Q(color[20]), .C(LED_c), .D(n17946));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_DFF color_21__54 (.Q(color[21]), .C(LED_c), .D(n17945));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_LUT4 add_3184_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n28110), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF color_22__53 (.Q(color[22]), .C(LED_c), .D(n17943));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4569), .I3(n29215), .O(n3_adj_3982)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n27975), 
            .O(n6804)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_32 (.CI(n29215), 
            .I0(GND_net), .I1(n3_adj_4569), .CO(n29216));
    SB_LUT4 div_46_i1536_3_lut (.I0(n2278), .I1(n6837), .I2(n2288), .I3(GND_net), 
            .O(n2371));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1536_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4570), .I3(n29214), .O(n4_adj_3981)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1710_3_lut_3_lut (.I0(n2558), .I1(n6897), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1711_3_lut_3_lut (.I0(n2558), .I1(n6898), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3184_17 (.CI(n28110), .I0(n2707), .I1(n86), .CO(n28111));
    SB_LUT4 blue_1137_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(blue[3]), 
            .I3(n28308), .O(n42_adj_4151)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13607_3_lut (.I0(Kp[7]), .I1(\data_in_frame[2] [7]), .I2(n35752), 
            .I3(GND_net), .O(n18114));   // verilog/coms.v(126[12] 289[6])
    defparam i13607_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_849_3 (.CI(n28545), .I0(n1258), 
            .I1(GND_net), .CO(n28546));
    SB_CARRY communication_counter_31__I_0_add_849_2 (.CI(VCC_net), .I0(n1358), 
            .I1(VCC_net), .CO(n28545));
    SB_LUT4 communication_counter_31__I_0_add_916_12_lut (.I0(n1382), .I1(n1349), 
            .I2(VCC_net), .I3(n28544), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_916_11_lut (.I0(GND_net), .I1(n1350), 
            .I2(VCC_net), .I3(n28543), .O(n1417_adj_4154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n27974), 
            .O(n6805)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_916_11 (.CI(n28543), .I0(n1350), 
            .I1(VCC_net), .CO(n28544));
    SB_CARRY blue_1137_add_4_5 (.CI(n28308), .I0(GND_net), .I1(blue[3]), 
            .CO(n28309));
    SB_LUT4 div_46_i1715_3_lut_3_lut (.I0(n2558), .I1(n6902), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3184_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n28109), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_916_10_lut (.I0(GND_net), .I1(n1351), 
            .I2(VCC_net), .I3(n28542), .O(n1418_adj_4155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4002), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i809_3_lut (.I0(n375), .I1(n6685), .I2(n1193), .I3(GND_net), 
            .O(n1299));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i809_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_add_916_10 (.CI(n28542), .I0(n1351), 
            .I1(VCC_net), .CO(n28543));
    SB_LUT4 blue_1137_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(blue[2]), 
            .I3(n28307), .O(n43_adj_4152)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_916_9_lut (.I0(GND_net), .I1(n1352), 
            .I2(VCC_net), .I3(n28541), .O(n1419_adj_4156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_17 (.CI(n27974), .I0(n2169), .I1(n85), .CO(n27975));
    SB_LUT4 add_3178_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n27973), 
            .O(n6806)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1137_add_4_4 (.CI(n28307), .I0(GND_net), .I1(blue[2]), 
            .CO(n28308));
    SB_CARRY add_555_11 (.CI(n27576), .I0(n41708), .I1(n16), .CO(n27577));
    SB_CARRY add_3184_16 (.CI(n28109), .I0(n2708), .I1(n87), .CO(n28110));
    SB_LUT4 blue_1137_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(blue[1]), 
            .I3(n28306), .O(n44_adj_4153)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_916_9 (.CI(n28541), .I0(n1352), 
            .I1(VCC_net), .CO(n28542));
    SB_LUT4 div_46_i890_3_lut (.I0(n1299), .I1(n6695), .I2(n1316), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i890_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_31 (.CI(n29214), 
            .I0(GND_net), .I1(n4_adj_4570), .CO(n29215));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4571), .I3(n29213), .O(n5_adj_3980)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i969_3_lut (.I0(n1419), .I1(n6706), .I2(n1436), .I3(GND_net), 
            .O(n1536));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3184_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n28108), 
            .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_916_8_lut (.I0(GND_net), .I1(n1353), 
            .I2(VCC_net), .I3(n28540), .O(n1420_adj_4157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1597_3_lut (.I0(n2371), .I1(n6857), .I2(n2381), .I3(GND_net), 
            .O(n2461));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1597_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1046_3_lut (.I0(n1536), .I1(n6718), .I2(n1553), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1121_3_lut (.I0(n1650), .I1(n6731), .I2(n1667), .I3(GND_net), 
            .O(n1761));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1194_3_lut (.I0(n1761), .I1(n6745), .I2(n1778), .I3(GND_net), 
            .O(n1869));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1265_3_lut (.I0(n1869), .I1(n6760), .I2(n1886), .I3(GND_net), 
            .O(n1974));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1334_3_lut (.I0(n1974), .I1(n6776), .I2(n1991), .I3(GND_net), 
            .O(n2076));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1334_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_555_10_lut (.I0(duty[8]), .I1(n41708), .I2(n17), .I3(n27575), 
            .O(pwm_setpoint_22__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1401_3_lut (.I0(n2076), .I1(n6793), .I2(n2093), .I3(GND_net), 
            .O(n2175));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1466_3_lut (.I0(n2175), .I1(n6811), .I2(n2192), .I3(GND_net), 
            .O(n2271));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1529_3_lut (.I0(n2271), .I1(n6830), .I2(n2288), .I3(GND_net), 
            .O(n2364));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1529_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1590_3_lut (.I0(n2364), .I1(n6850), .I2(n2381), .I3(GND_net), 
            .O(n2454));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1118_3_lut (.I0(n1647), .I1(n6728), .I2(n1667), .I3(GND_net), 
            .O(n1758));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13611_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13950), .I3(GND_net), .O(n18118));   // verilog/coms.v(126[12] 289[6])
    defparam i13611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13612_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13950), .I3(GND_net), .O(n18119));   // verilog/coms.v(126[12] 289[6])
    defparam i13612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1191_3_lut (.I0(n1758), .I1(n6742), .I2(n1778), .I3(GND_net), 
            .O(n1866));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1262_3_lut (.I0(n1866), .I1(n6757), .I2(n1886), .I3(GND_net), 
            .O(n1971));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1331_3_lut (.I0(n1971), .I1(n6773), .I2(n1991), .I3(GND_net), 
            .O(n2073));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1398_3_lut (.I0(n2073), .I1(n6790), .I2(n2093), .I3(GND_net), 
            .O(n2172));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13613_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13950), .I3(GND_net), .O(n18120));   // verilog/coms.v(126[12] 289[6])
    defparam i13613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[10]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_46_i1463_3_lut (.I0(n2172), .I1(n6808), .I2(n2192), .I3(GND_net), 
            .O(n2268));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1526_3_lut (.I0(n2268), .I1(n6827), .I2(n2288), .I3(GND_net), 
            .O(n2361));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1526_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1587_3_lut (.I0(n2361), .I1(n6847), .I2(n2381), .I3(GND_net), 
            .O(n2451));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4449));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mux_77_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_107[10]), 
            .I2(n15), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13614_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13950), .I3(GND_net), .O(n18121));   // verilog/coms.v(126[12] 289[6])
    defparam i13614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4004), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i639_3_lut (.I0(n373), .I1(n6666), .I2(n938), .I3(GND_net), 
            .O(n1048));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i724_3_lut (.I0(n1048), .I1(n6674), .I2(n1067), .I3(GND_net), 
            .O(n1174));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i807_3_lut (.I0(n1174), .I1(n6683), .I2(n1193), .I3(GND_net), 
            .O(n1297));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i888_3_lut (.I0(n1297), .I1(n6693), .I2(n1316), .I3(GND_net), 
            .O(n1417));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i967_3_lut (.I0(n1417), .I1(n6704), .I2(n1436), .I3(GND_net), 
            .O(n1534));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13615_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13950), .I3(GND_net), .O(n18122));   // verilog/coms.v(126[12] 289[6])
    defparam i13615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13616_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13950), .I3(GND_net), .O(n18123));   // verilog/coms.v(126[12] 289[6])
    defparam i13616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13617_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13950), .I3(GND_net), .O(n18124));   // verilog/coms.v(126[12] 289[6])
    defparam i13617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1044_3_lut (.I0(n1534), .I1(n6716), .I2(n1553), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1119_3_lut (.I0(n1648), .I1(n6729), .I2(n1667), .I3(GND_net), 
            .O(n1759));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1192_3_lut (.I0(n1759), .I1(n6743), .I2(n1778), .I3(GND_net), 
            .O(n1867));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1263_3_lut (.I0(n1867), .I1(n6758), .I2(n1886), .I3(GND_net), 
            .O(n1972));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1332_3_lut (.I0(n1972), .I1(n6774), .I2(n1991), .I3(GND_net), 
            .O(n2074));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13618_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13950), .I3(GND_net), .O(n18125));   // verilog/coms.v(126[12] 289[6])
    defparam i13618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13619_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13950), .I3(GND_net), .O(n18126));   // verilog/coms.v(126[12] 289[6])
    defparam i13619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13620_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13950), .I3(GND_net), .O(n18127));   // verilog/coms.v(126[12] 289[6])
    defparam i13620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13621_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13950), .I3(GND_net), .O(n18128));   // verilog/coms.v(126[12] 289[6])
    defparam i13621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1399_3_lut (.I0(n2074), .I1(n6791), .I2(n2093), .I3(GND_net), 
            .O(n2173));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1464_3_lut (.I0(n2173), .I1(n6809), .I2(n2192), .I3(GND_net), 
            .O(n2269));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1527_3_lut (.I0(n2269), .I1(n6828), .I2(n2288), .I3(GND_net), 
            .O(n2362));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1527_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1588_3_lut (.I0(n2362), .I1(n6848), .I2(n2381), .I3(GND_net), 
            .O(n2452));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4447));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33374_3_lut (.I0(n369), .I1(n558), .I2(n392), .I3(GND_net), 
            .O(n510));
    defparam i33374_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i13622_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13950), .I3(GND_net), .O(n18129));   // verilog/coms.v(126[12] 289[6])
    defparam i13622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[11]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_107[11]), 
            .I2(n15), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4012), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32988_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n38981));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i32988_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1553 (.I0(n38981), .I1(n16472), .I2(n99), .I3(n5_adj_4553), 
            .O(n392));
    defparam i1_4_lut_adj_1553.LUT_INIT = 16'hefce;
    SB_LUT4 i1_4_lut_adj_1554 (.I0(n224), .I1(n99), .I2(n16472), .I3(n558), 
            .O(n5_adj_4553));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i1_4_lut_adj_1554.LUT_INIT = 16'h555d;
    SB_LUT4 div_46_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(n93), .I1(n16529), .I2(GND_net), .I3(GND_net), 
            .O(n16526));
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_555_10 (.CI(n27575), .I0(n41708), .I1(n17), .CO(n27576));
    SB_LUT4 i13623_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13950), .I3(GND_net), .O(n18130));   // verilog/coms.v(126[12] 289[6])
    defparam i13623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1556 (.I0(n96), .I1(n16520), .I2(GND_net), .I3(GND_net), 
            .O(n16517));
    defparam i1_2_lut_adj_1556.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i22704_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3953));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22704_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_i274_4_lut (.I0(n5_adj_4553), .I1(n2_adj_3953), .I2(n392), 
            .I3(n99), .O(n34342));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i274_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_46_i1716_3_lut_3_lut (.I0(n2558), .I1(n6903), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46_adj_4241));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1557 (.I0(n46_adj_4241), .I1(n16514), .I2(n98), 
            .I3(n34342), .O(n533));
    defparam i1_4_lut_adj_1557.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4007), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22744_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3937));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22744_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33371_3_lut (.I0(n370), .I1(n558), .I2(n533), .I3(GND_net), 
            .O(n649));
    defparam i33371_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_46_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i460_4_lut (.I0(n649), .I1(n2_adj_3937), .I2(n671), 
            .I3(n99), .O(n784));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i460_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_46_i549_4_lut (.I0(n784), .I1(n4_adj_4612), .I2(n806), 
            .I3(n98), .O(n916));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i549_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_46_i636_3_lut (.I0(n916), .I1(n6663), .I2(n938), .I3(GND_net), 
            .O(n1045));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i721_3_lut (.I0(n1045), .I1(n6671), .I2(n1067), .I3(GND_net), 
            .O(n1171));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i804_3_lut (.I0(n1171), .I1(n6680), .I2(n1193), .I3(GND_net), 
            .O(n1294));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i885_3_lut (.I0(n1294), .I1(n6690), .I2(n1316), .I3(GND_net), 
            .O(n1414));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i964_3_lut (.I0(n1414), .I1(n6701), .I2(n1436), .I3(GND_net), 
            .O(n1531));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13624_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13950), .I3(GND_net), .O(n18131));   // verilog/coms.v(126[12] 289[6])
    defparam i13624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13625_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13950), .I3(GND_net), .O(n18132));   // verilog/coms.v(126[12] 289[6])
    defparam i13625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13626_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13950), .I3(GND_net), .O(n18133));   // verilog/coms.v(126[12] 289[6])
    defparam i13626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13627_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13950), .I3(GND_net), .O(n18134));   // verilog/coms.v(126[12] 289[6])
    defparam i13627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13628_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13950), .I3(GND_net), .O(n18135));   // verilog/coms.v(126[12] 289[6])
    defparam i13628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13629_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13950), .I3(GND_net), .O(n18136));   // verilog/coms.v(126[12] 289[6])
    defparam i13629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13630_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13950), .I3(GND_net), .O(n18137));   // verilog/coms.v(126[12] 289[6])
    defparam i13630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13631_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13950), .I3(GND_net), .O(n18138));   // verilog/coms.v(126[12] 289[6])
    defparam i13631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13632_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13950), .I3(GND_net), .O(n18139));   // verilog/coms.v(126[12] 289[6])
    defparam i13632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13633_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13950), .I3(GND_net), .O(n18140));   // verilog/coms.v(126[12] 289[6])
    defparam i13633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1041_3_lut (.I0(n1531), .I1(n6713), .I2(n1553), .I3(GND_net), 
            .O(n1645));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1116_3_lut (.I0(n1645), .I1(n6726), .I2(n1667), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1189_3_lut (.I0(n1756), .I1(n6740), .I2(n1778), .I3(GND_net), 
            .O(n1864));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1260_3_lut (.I0(n1864), .I1(n6755), .I2(n1886), .I3(GND_net), 
            .O(n1969));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1329_3_lut (.I0(n1969), .I1(n6771), .I2(n1991), .I3(GND_net), 
            .O(n2071));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1396_3_lut (.I0(n2071), .I1(n6788), .I2(n2093), .I3(GND_net), 
            .O(n2170));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1461_3_lut (.I0(n2170), .I1(n6806), .I2(n2192), .I3(GND_net), 
            .O(n2266));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1524_3_lut (.I0(n2266), .I1(n6825), .I2(n2288), .I3(GND_net), 
            .O(n2359));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1656_3_lut (.I0(n2461), .I1(n6878), .I2(n2471), .I3(GND_net), 
            .O(n2548));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13634_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13950), .I3(GND_net), .O(n18141));   // verilog/coms.v(126[12] 289[6])
    defparam i13634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13635_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13950), .I3(GND_net), .O(n18142));   // verilog/coms.v(126[12] 289[6])
    defparam i13635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1266_3_lut (.I0(n1857), .I1(n1924), 
            .I2(n1877), .I3(GND_net), .O(n1956));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1333_3_lut (.I0(n1956), .I1(n2023), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1400_3_lut (.I0(n2055), .I1(n2122), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1467_3_lut (.I0(n2154), .I1(n2221), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1265_3_lut (.I0(n1856), .I1(n1923), 
            .I2(n1877), .I3(GND_net), .O(n1955));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1585_3_lut (.I0(n2359), .I1(n6845), .I2(n2381), .I3(GND_net), 
            .O(n2449));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4451));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4438));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_3997), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1199_3_lut (.I0(n380), .I1(n6750), .I2(n1778), .I3(GND_net), 
            .O(n1874));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1270_3_lut (.I0(n1874), .I1(n6765), .I2(n1886), .I3(GND_net), 
            .O(n1979));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1339_3_lut (.I0(n1979), .I1(n6781), .I2(n1991), .I3(GND_net), 
            .O(n2081));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1406_3_lut (.I0(n2081), .I1(n6798), .I2(n2093), .I3(GND_net), 
            .O(n2180));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1332_3_lut (.I0(n1955), .I1(n2022), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1399_3_lut (.I0(n2054), .I1(n2121), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1466_3_lut (.I0(n2153), .I1(n2220), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1264_3_lut (.I0(n1855), .I1(n1922), 
            .I2(n1877), .I3(GND_net), .O(n1954));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1471_3_lut (.I0(n2180), .I1(n6816), .I2(n2192), .I3(GND_net), 
            .O(n2276));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1534_3_lut (.I0(n2276), .I1(n6835), .I2(n2288), .I3(GND_net), 
            .O(n2369));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1534_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44_adj_4243));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34231_3_lut (.I0(n44_adj_4243), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n40553));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34231_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1558 (.I0(n40553), .I1(n16517), .I2(n97), .I3(n34344), 
            .O(n671));
    defparam i1_4_lut_adj_1558.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4006), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4244));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34201_3_lut (.I0(n42_adj_4244), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n40523));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34201_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34202_3_lut (.I0(n40523), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n40524));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34202_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1559 (.I0(n40524), .I1(n16520), .I2(n96), .I3(n34346), 
            .O(n806));
    defparam i1_4_lut_adj_1559.LUT_INIT = 16'hefce;
    SB_LUT4 i22776_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22776_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33368_3_lut (.I0(n371), .I1(n558), .I2(n671), .I3(GND_net), 
            .O(n785));
    defparam i33368_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 communication_counter_31__I_0_i1331_3_lut (.I0(n1954), .I1(n2021), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3178_16 (.CI(n27973), .I0(n2170), .I1(n86), .CO(n27974));
    SB_LUT4 div_46_i1712_3_lut_3_lut (.I0(n2558), .I1(n6899), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34228_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4245), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4246));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_570_i44_3_lut (.I0(n42_adj_4247), .I1(n96), 
            .I2(n45_adj_4249), .I3(GND_net), .O(n44_adj_4248));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34233_4_lut (.I0(n44_adj_4248), .I1(n40_adj_4246), .I2(n45_adj_4249), 
            .I3(n39549), .O(n40555));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34233_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1560 (.I0(n40555), .I1(n16523), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1560.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i550_4_lut (.I0(n785), .I1(n2), .I2(n806), .I3(n99), 
            .O(n917));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i550_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_46_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4250));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_657_i42_3_lut (.I0(n40_adj_4251), .I1(n96), 
            .I2(n43_adj_4253), .I3(GND_net), .O(n42_adj_4252));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34496_4_lut (.I0(n42_adj_4252), .I1(n38_adj_4250), .I2(n43_adj_4253), 
            .I3(n39537), .O(n40818));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34496_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34497_3_lut (.I0(n40818), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n40819));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34497_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1561 (.I0(n40819), .I1(n16526), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1561.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i637_3_lut (.I0(n917), .I1(n6664), .I2(n938), .I3(GND_net), 
            .O(n1046));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36_adj_4255));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3178_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n27972), 
            .O(n6807)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1262_rep_50_3_lut (.I0(n1853), 
            .I1(n1920), .I2(n1877), .I3(GND_net), .O(n1952));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1262_rep_50_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1329_3_lut (.I0(n1952), .I1(n2019), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1396_3_lut (.I0(n2051), .I1(n2118), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2150));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_742_i40_3_lut (.I0(n38_adj_4256), .I1(n96), 
            .I2(n41_adj_4258), .I3(GND_net), .O(n40_adj_4257));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34502_4_lut (.I0(n40_adj_4257), .I1(n36_adj_4255), .I2(n41_adj_4258), 
            .I3(n39527), .O(n40824));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34502_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34503_3_lut (.I0(n40824), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n40825));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34503_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34407_3_lut (.I0(n40825), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n40729));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34407_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1562 (.I0(n40729), .I1(n16529), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1562.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i722_3_lut (.I0(n1046), .I1(n6672), .I2(n1067), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34_adj_4259));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34195_3_lut (.I0(n34_adj_4259), .I1(n95), .I2(n41_adj_4263), 
            .I3(GND_net), .O(n40517));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34195_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34196_3_lut (.I0(n40517), .I1(n94), .I2(n43_adj_4264), .I3(GND_net), 
            .O(n40518));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34196_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33778_4_lut (.I0(n43_adj_4264), .I1(n41_adj_4263), .I2(n39_adj_4262), 
            .I3(n39519), .O(n40100));
    defparam i33778_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_825_i38_3_lut (.I0(n36_adj_4260), .I1(n96), 
            .I2(n39_adj_4262), .I3(GND_net), .O(n38_adj_4261));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33624_3_lut (.I0(n40518), .I1(n93), .I2(n45_adj_4265), .I3(GND_net), 
            .O(n39946));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33624_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34239_4_lut (.I0(n39946), .I1(n38_adj_4261), .I2(n45_adj_4265), 
            .I3(n40100), .O(n40561));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34239_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1563 (.I0(n40561), .I1(n16532), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1563.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i805_3_lut (.I0(n1172), .I1(n6681), .I2(n1193), .I3(GND_net), 
            .O(n1295));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1463_3_lut (.I0(n2150), .I1(n2217), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1261_3_lut (.I0(n1852), .I1(n1919), 
            .I2(n1877), .I3(GND_net), .O(n1951));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1328_3_lut (.I0(n1951), .I1(n2018), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32_adj_4267));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34193_3_lut (.I0(n32_adj_4267), .I1(n95), .I2(n39_adj_4270), 
            .I3(GND_net), .O(n40515));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34193_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34194_3_lut (.I0(n40515), .I1(n94), .I2(n41_adj_4271), .I3(GND_net), 
            .O(n40516));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34194_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33770_4_lut (.I0(n41_adj_4271), .I1(n39_adj_4270), .I2(n37_adj_4269), 
            .I3(n39507), .O(n40092));
    defparam i33770_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34241_3_lut (.I0(n34_adj_4268), .I1(n96), .I2(n37_adj_4269), 
            .I3(GND_net), .O(n40563));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34241_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33626_3_lut (.I0(n40516), .I1(n93), .I2(n43_adj_4272), .I3(GND_net), 
            .O(n39948));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33626_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34404_4_lut (.I0(n39948), .I1(n40563), .I2(n43_adj_4272), 
            .I3(n40092), .O(n40726));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34404_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34405_3_lut (.I0(n40726), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n40727));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34405_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1564 (.I0(n40727), .I1(n16475), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1564.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i886_3_lut (.I0(n1295), .I1(n6691), .I2(n1316), .I3(GND_net), 
            .O(n1415));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4274));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33163_4_lut (.I0(n37_adj_4279), .I1(n35_adj_4278), .I2(n33_adj_4276), 
            .I3(n31_adj_4274), .O(n39485));
    defparam i33163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_985_i42_3_lut (.I0(n34_adj_4277), .I1(n91), 
            .I2(n45_adj_4284), .I3(GND_net), .O(n42_adj_4282));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4273));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34191_3_lut (.I0(n30_adj_4273), .I1(n95), .I2(n37_adj_4279), 
            .I3(GND_net), .O(n40513));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34191_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34192_3_lut (.I0(n40513), .I1(n94), .I2(n39_adj_4280), .I3(GND_net), 
            .O(n40514));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34192_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33157_4_lut (.I0(n43_adj_4283), .I1(n41_adj_4281), .I2(n39_adj_4280), 
            .I3(n39485), .O(n39479));
    defparam i33157_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 communication_counter_31__I_0_i1395_3_lut (.I0(n2050), .I1(n2117), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1462_3_lut (.I0(n2149), .I1(n2216), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13636_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13950), .I3(GND_net), .O(n18143));   // verilog/coms.v(126[12] 289[6])
    defparam i13636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13637_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13950), .I3(GND_net), .O(n18144));   // verilog/coms.v(126[12] 289[6])
    defparam i13637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34243_4_lut (.I0(n42_adj_4282), .I1(n32_adj_4275), .I2(n45_adj_4284), 
            .I3(n39475), .O(n40565));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34243_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33629_3_lut (.I0(n40514), .I1(n93), .I2(n41_adj_4281), .I3(GND_net), 
            .O(n39951));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33629_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34534_4_lut (.I0(n39951), .I1(n40565), .I2(n45_adj_4284), 
            .I3(n39479), .O(n40856));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34534_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(n40856), .I1(n16535), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i965_3_lut (.I0(n1415), .I1(n6702), .I2(n1436), .I3(GND_net), 
            .O(n1532));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4286));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33145_4_lut (.I0(n35_adj_4291), .I1(n33_adj_4290), .I2(n31_adj_4288), 
            .I3(n29_adj_4286), .O(n39467));
    defparam i33145_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1062_i40_3_lut (.I0(n32_adj_4289), .I1(n91), 
            .I2(n43_adj_4296), .I3(GND_net), .O(n40_adj_4294));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4285));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34185_3_lut (.I0(n28_adj_4285), .I1(n95), .I2(n35_adj_4291), 
            .I3(GND_net), .O(n40507));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34185_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34186_3_lut (.I0(n40507), .I1(n94), .I2(n37_adj_4292), .I3(GND_net), 
            .O(n40508));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34186_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33138_4_lut (.I0(n41_adj_4295), .I1(n39_adj_4293), .I2(n37_adj_4292), 
            .I3(n39467), .O(n39460));
    defparam i33138_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34494_4_lut (.I0(n40_adj_4294), .I1(n30_adj_4287), .I2(n43_adj_4296), 
            .I3(n39455), .O(n40816));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34494_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33631_3_lut (.I0(n40508), .I1(n93), .I2(n39_adj_4293), .I3(GND_net), 
            .O(n39953));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33631_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34607_4_lut (.I0(n39953), .I1(n40816), .I2(n43_adj_4296), 
            .I3(n39460), .O(n40929));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34607_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34608_3_lut (.I0(n40929), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n40930));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34608_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(n40930), .I1(n16538), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1042_3_lut (.I0(n1532), .I1(n6714), .I2(n1553), .I3(GND_net), 
            .O(n1646));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3178_15 (.CI(n27972), .I0(n2171), .I1(n87), .CO(n27973));
    SB_LUT4 i13638_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13950), .I3(GND_net), .O(n18145));   // verilog/coms.v(126[12] 289[6])
    defparam i13638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13639_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13950), .I3(GND_net), .O(n18146));   // verilog/coms.v(126[12] 289[6])
    defparam i13639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13640_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13950), .I3(GND_net), .O(n18147));   // verilog/coms.v(126[12] 289[6])
    defparam i13640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4298));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33118_4_lut (.I0(n33_adj_4303), .I1(n31_adj_4302), .I2(n29_adj_4300), 
            .I3(n27_adj_4298), .O(n39440));
    defparam i33118_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1137_i38_3_lut (.I0(n30_adj_4301), .I1(n91), 
            .I2(n41_adj_4308), .I3(GND_net), .O(n38_adj_4306));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_4297));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34183_3_lut (.I0(n26_adj_4297), .I1(n95), .I2(n33_adj_4303), 
            .I3(GND_net), .O(n40505));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34183_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34184_3_lut (.I0(n40505), .I1(n94), .I2(n35_adj_4304), .I3(GND_net), 
            .O(n40506));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34184_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33112_4_lut (.I0(n39_adj_4307), .I1(n37_adj_4305), .I2(n35_adj_4304), 
            .I3(n39440), .O(n39434));
    defparam i33112_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34504_4_lut (.I0(n38_adj_4306), .I1(n28_adj_4299), .I2(n41_adj_4308), 
            .I3(n39432), .O(n40826));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34504_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33633_3_lut (.I0(n40506), .I1(n93), .I2(n37_adj_4305), .I3(GND_net), 
            .O(n39955));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33633_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34613_4_lut (.I0(n39955), .I1(n40826), .I2(n41_adj_4308), 
            .I3(n39434), .O(n40935));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34613_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34614_3_lut (.I0(n40935), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n40936));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34614_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34580_3_lut (.I0(n40936), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n40902));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34580_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(n40902), .I1(n16541), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1117_3_lut (.I0(n1646), .I1(n6727), .I2(n1667), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4310));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33053_4_lut (.I0(n31_adj_4316), .I1(n29_adj_4314), .I2(n27_adj_4312), 
            .I3(n25_adj_4310), .O(n39374));
    defparam i33053_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33045_4_lut (.I0(n37_adj_4321), .I1(n35_adj_4319), .I2(n33_adj_4318), 
            .I3(n39374), .O(n39366));
    defparam i33045_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13641_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13950), .I3(GND_net), .O(n18148));   // verilog/coms.v(126[12] 289[6])
    defparam i13641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1259_3_lut (.I0(n1850), .I1(n1917), 
            .I2(n1877), .I3(GND_net), .O(n1949));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1326_3_lut (.I0(n1949), .I1(n2016), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1393_3_lut (.I0(n2048), .I1(n2115), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1460_3_lut (.I0(n2147), .I1(n2214), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1258_3_lut (.I0(n1849), .I1(n1916), 
            .I2(n1877), .I3(GND_net), .O(n1948));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1325_3_lut (.I0(n1948), .I1(n2015), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1392_3_lut (.I0(n2047), .I1(n2114), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1459_3_lut (.I0(n2146), .I1(n2213), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4309));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1210_i32_3_lut (.I0(n30_adj_4315), .I1(n93), 
            .I2(n35_adj_4319), .I3(GND_net), .O(n32_adj_4317));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1210_i36_3_lut (.I0(n28_adj_4313), .I1(n91), 
            .I2(n39_adj_4322), .I3(GND_net), .O(n36_adj_4320));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34547_4_lut (.I0(n36_adj_4320), .I1(n26_adj_4311), .I2(n39_adj_4322), 
            .I3(n39342), .O(n40869));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34547_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34548_3_lut (.I0(n40869), .I1(n90), .I2(n41_adj_4323), .I3(GND_net), 
            .O(n40870));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34548_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34493_3_lut (.I0(n40870), .I1(n89), .I2(n43_adj_4324), .I3(GND_net), 
            .O(n40815));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34493_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34213_4_lut (.I0(n43_adj_4324), .I1(n41_adj_4323), .I2(n39_adj_4322), 
            .I3(n39366), .O(n40535));
    defparam i34213_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34012_4_lut (.I0(n32_adj_4317), .I1(n24_adj_4309), .I2(n35_adj_4319), 
            .I3(n39372), .O(n40334));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34012_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34425_3_lut (.I0(n40815), .I1(n88), .I2(n45_adj_4326), .I3(GND_net), 
            .O(n44_adj_4325));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34425_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34014_4_lut (.I0(n44_adj_4325), .I1(n40334), .I2(n45_adj_4326), 
            .I3(n40535), .O(n40336));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34014_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1568 (.I0(n40336), .I1(n16485), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1568.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1190_3_lut (.I0(n1757), .I1(n6741), .I2(n1778), .I3(GND_net), 
            .O(n1865));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4328));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i32971_4_lut (.I0(n29_adj_4334), .I1(n27_adj_4332), .I2(n25_adj_4330), 
            .I3(n23_adj_4328), .O(n39291));
    defparam i32971_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32963_4_lut (.I0(n35_adj_4339), .I1(n33_adj_4337), .I2(n31_adj_4336), 
            .I3(n39291), .O(n39283));
    defparam i32963_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4327));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1281_i30_3_lut (.I0(n28_adj_4333), .I1(n93), 
            .I2(n33_adj_4337), .I3(GND_net), .O(n30_adj_4335));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1281_i34_3_lut (.I0(n26_adj_4331), .I1(n91), 
            .I2(n37_adj_4340), .I3(GND_net), .O(n34_adj_4338));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34549_4_lut (.I0(n34_adj_4338), .I1(n24_adj_4329), .I2(n37_adj_4340), 
            .I3(n39281), .O(n40871));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34549_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34550_3_lut (.I0(n40871), .I1(n90), .I2(n39_adj_4341), .I3(GND_net), 
            .O(n40872));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34550_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34491_3_lut (.I0(n40872), .I1(n89), .I2(n41_adj_4342), .I3(GND_net), 
            .O(n40813));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34491_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34179_4_lut (.I0(n41_adj_4342), .I1(n39_adj_4341), .I2(n37_adj_4340), 
            .I3(n39283), .O(n40501));
    defparam i34179_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34360_4_lut (.I0(n30_adj_4335), .I1(n22_adj_4327), .I2(n33_adj_4337), 
            .I3(n39287), .O(n40682));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34360_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34427_3_lut (.I0(n40813), .I1(n88), .I2(n43_adj_4344), .I3(GND_net), 
            .O(n42_adj_4343));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34427_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34526_4_lut (.I0(n42_adj_4343), .I1(n40682), .I2(n43_adj_4344), 
            .I3(n40501), .O(n40848));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34526_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34527_3_lut (.I0(n40848), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n40849));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34527_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(n40849), .I1(n16544), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1261_3_lut (.I0(n1865), .I1(n6756), .I2(n1886), .I3(GND_net), 
            .O(n1970));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4350));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i32912_4_lut (.I0(n27_adj_4356), .I1(n25_adj_4354), .I2(n23_adj_4352), 
            .I3(n21_adj_4350), .O(n39232));
    defparam i32912_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32900_4_lut (.I0(n33_adj_4361), .I1(n31_adj_4359), .I2(n29_adj_4358), 
            .I3(n39232), .O(n39220));
    defparam i32900_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4349));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1350_i28_3_lut (.I0(n26_adj_4355), .I1(n93), 
            .I2(n31_adj_4359), .I3(GND_net), .O(n28_adj_4357));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1350_i32_3_lut (.I0(n24_adj_4353), .I1(n91), 
            .I2(n35_adj_4362), .I3(GND_net), .O(n32_adj_4360));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34551_4_lut (.I0(n32_adj_4360), .I1(n22_adj_4351), .I2(n35_adj_4362), 
            .I3(n39216), .O(n40873));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34551_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34552_3_lut (.I0(n40873), .I1(n90), .I2(n37_adj_4363), .I3(GND_net), 
            .O(n40874));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34552_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34489_3_lut (.I0(n40874), .I1(n89), .I2(n39_adj_4364), .I3(GND_net), 
            .O(n40811));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34489_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34161_4_lut (.I0(n39_adj_4364), .I1(n37_adj_4363), .I2(n35_adj_4362), 
            .I3(n39220), .O(n40483));
    defparam i34161_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34553_4_lut (.I0(n28_adj_4357), .I1(n20_adj_4349), .I2(n31_adj_4359), 
            .I3(n39230), .O(n40875));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34553_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34429_3_lut (.I0(n40811), .I1(n88), .I2(n41_adj_4365), .I3(GND_net), 
            .O(n40751));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34429_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34624_4_lut (.I0(n40751), .I1(n40875), .I2(n41_adj_4365), 
            .I3(n40483), .O(n40946));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34624_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34625_3_lut (.I0(n40946), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n40947));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34625_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i34566_3_lut (.I0(n40947), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n40888));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34566_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1570 (.I0(n40888), .I1(n16491), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1570.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1330_3_lut (.I0(n1970), .I1(n6772), .I2(n1991), .I3(GND_net), 
            .O(n2072));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4369));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i32863_4_lut (.I0(n25_adj_4375), .I1(n23_adj_4373), .I2(n21_adj_4371), 
            .I3(n19_adj_4369), .O(n39183));
    defparam i32863_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32851_4_lut (.I0(n31_adj_4380), .I1(n29_adj_4378), .I2(n27_adj_4377), 
            .I3(n39183), .O(n39171));
    defparam i32851_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34145_4_lut (.I0(n37_adj_4383), .I1(n35_adj_4382), .I2(n33_adj_4381), 
            .I3(n39171), .O(n40467));
    defparam i34145_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4368));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34352_3_lut (.I0(n18_adj_4368), .I1(n87), .I2(n41_adj_4385), 
            .I3(GND_net), .O(n40674));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34352_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34353_3_lut (.I0(n40674), .I1(n86), .I2(n43_adj_4387), .I3(GND_net), 
            .O(n40675));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34353_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33486_4_lut (.I0(n43_adj_4387), .I1(n41_adj_4385), .I2(n29_adj_4378), 
            .I3(n39181), .O(n39808));
    defparam i33486_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1417_i26_3_lut (.I0(n24_adj_4374), .I1(n93), 
            .I2(n29_adj_4378), .I3(GND_net), .O(n26_adj_4376));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34262_3_lut (.I0(n40675), .I1(n85), .I2(n45_adj_4388), .I3(GND_net), 
            .O(n42_adj_4386));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34262_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1718_3_lut_3_lut (.I0(n2558), .I1(n6905), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13642_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13950), .I3(GND_net), .O(n18149));   // verilog/coms.v(126[12] 289[6])
    defparam i13642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13643_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13950), .I3(GND_net), .O(n18150));   // verilog/coms.v(126[12] 289[6])
    defparam i13643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13644_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13950), .I3(GND_net), .O(n18151));   // verilog/coms.v(126[12] 289[6])
    defparam i13644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i30_3_lut (.I0(n22_adj_4372), .I1(n91), 
            .I2(n33_adj_4381), .I3(GND_net), .O(n30_adj_4379));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34555_4_lut (.I0(n30_adj_4379), .I1(n20_adj_4370), .I2(n33_adj_4381), 
            .I3(n39168), .O(n40877));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34555_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34556_3_lut (.I0(n40877), .I1(n90), .I2(n35_adj_4382), .I3(GND_net), 
            .O(n40878));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34556_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34485_3_lut (.I0(n40878), .I1(n89), .I2(n37_adj_4383), .I3(GND_net), 
            .O(n40807));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34485_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33490_4_lut (.I0(n43_adj_4387), .I1(n41_adj_4385), .I2(n39_adj_4384), 
            .I3(n40467), .O(n39812));
    defparam i33490_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34018_4_lut (.I0(n42_adj_4386), .I1(n26_adj_4376), .I2(n45_adj_4388), 
            .I3(n39808), .O(n40340));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34018_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34435_3_lut (.I0(n40807), .I1(n88), .I2(n39_adj_4384), .I3(GND_net), 
            .O(n40757));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34435_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34020_4_lut (.I0(n40757), .I1(n40340), .I2(n45_adj_4388), 
            .I3(n39812), .O(n40342));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34020_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n40342), .I1(n16495), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1397_3_lut (.I0(n2072), .I1(n6789), .I2(n2093), .I3(GND_net), 
            .O(n2171));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4390));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i32813_4_lut (.I0(n23_adj_4396), .I1(n21_adj_4394), .I2(n19_adj_4392), 
            .I3(n17_adj_4390), .O(n39133));
    defparam i32813_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32807_4_lut (.I0(n29_adj_4400), .I1(n27_adj_4398), .I2(n25_adj_4397), 
            .I3(n39133), .O(n39127));
    defparam i32807_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34141_4_lut (.I0(n35_adj_4403), .I1(n33_adj_4402), .I2(n31_adj_4401), 
            .I3(n39127), .O(n40463));
    defparam i34141_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4389));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34348_3_lut (.I0(n16_adj_4389), .I1(n87), .I2(n39_adj_4405), 
            .I3(GND_net), .O(n40670));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34348_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34349_3_lut (.I0(n40670), .I1(n86), .I2(n41_adj_4406), .I3(GND_net), 
            .O(n40671));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34349_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33458_4_lut (.I0(n41_adj_4406), .I1(n39_adj_4405), .I2(n27_adj_4398), 
            .I3(n39131), .O(n39780));
    defparam i33458_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34267_3_lut (.I0(n22_adj_4395), .I1(n93), .I2(n27_adj_4398), 
            .I3(GND_net), .O(n40589));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34267_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34266_3_lut (.I0(n40671), .I1(n85), .I2(n43_adj_4407), .I3(GND_net), 
            .O(n40588));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34266_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13645_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13950), .I3(GND_net), .O(n18152));   // verilog/coms.v(126[12] 289[6])
    defparam i13645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13646_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13950), .I3(GND_net), .O(n18153));   // verilog/coms.v(126[12] 289[6])
    defparam i13646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13647_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13950), .I3(GND_net), .O(n18154));   // verilog/coms.v(126[12] 289[6])
    defparam i13647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13648_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13950), .I3(GND_net), .O(n18155));   // verilog/coms.v(126[12] 289[6])
    defparam i13648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13649_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13950), .I3(GND_net), .O(n18156));   // verilog/coms.v(126[12] 289[6])
    defparam i13649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13650_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13950), .I3(GND_net), .O(n18157));   // verilog/coms.v(126[12] 289[6])
    defparam i13650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i28_3_lut (.I0(n20_adj_4393), .I1(n91), 
            .I2(n31_adj_4401), .I3(GND_net), .O(n28_adj_4399));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34559_4_lut (.I0(n28_adj_4399), .I1(n18_adj_4391), .I2(n31_adj_4401), 
            .I3(n39125), .O(n40881));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34559_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34560_3_lut (.I0(n40881), .I1(n90), .I2(n33_adj_4402), .I3(GND_net), 
            .O(n40882));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34560_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34481_3_lut (.I0(n40882), .I1(n89), .I2(n35_adj_4403), .I3(GND_net), 
            .O(n40803));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34481_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33460_4_lut (.I0(n41_adj_4406), .I1(n39_adj_4405), .I2(n37_adj_4404), 
            .I3(n40463), .O(n39782));
    defparam i33460_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34346_4_lut (.I0(n40588), .I1(n40589), .I2(n43_adj_4407), 
            .I3(n39780), .O(n40668));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34346_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34437_3_lut (.I0(n40803), .I1(n88), .I2(n37_adj_4404), .I3(GND_net), 
            .O(n40759));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34437_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34571_4_lut (.I0(n40759), .I1(n40668), .I2(n43_adj_4407), 
            .I3(n39782), .O(n40893));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34571_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34572_3_lut (.I0(n40893), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n40894));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34572_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n40894), .I1(n16547), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i1462_3_lut (.I0(n2171), .I1(n6807), .I2(n2192), .I3(GND_net), 
            .O(n2267));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33400_4_lut (.I0(n37_adj_4424), .I1(n25_adj_4417), .I2(n23_adj_4416), 
            .I3(n21_adj_4414), .O(n39722));
    defparam i33400_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33932_4_lut (.I0(n19_adj_4412), .I1(n17_adj_4410), .I2(n2373), 
            .I3(n98), .O(n40254));
    defparam i33932_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34135_4_lut (.I0(n25_adj_4417), .I1(n23_adj_4416), .I2(n21_adj_4414), 
            .I3(n40254), .O(n40457));
    defparam i34135_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34133_4_lut (.I0(n31_adj_4421), .I1(n29_adj_4420), .I2(n27_adj_4419), 
            .I3(n40457), .O(n40455));
    defparam i34133_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33404_4_lut (.I0(n37_adj_4424), .I1(n35_adj_4423), .I2(n33_adj_4422), 
            .I3(n40455), .O(n39726));
    defparam i33404_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4408));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34175_3_lut (.I0(n14_adj_4408), .I1(n87), .I2(n37_adj_4424), 
            .I3(GND_net), .O(n40497));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34175_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34176_3_lut (.I0(n40497), .I1(n86), .I2(n39_adj_4425), .I3(GND_net), 
            .O(n40498));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34176_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1545_i40_3_lut (.I0(n22_adj_4415), .I1(n83), 
            .I2(n45_adj_4429), .I3(GND_net), .O(n40_adj_4426));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33391_4_lut (.I0(n43_adj_4428), .I1(n41_adj_4427), .I2(n39_adj_4425), 
            .I3(n39722), .O(n39713));
    defparam i33391_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34272_4_lut (.I0(n40_adj_4426), .I1(n20_adj_4413), .I2(n45_adj_4429), 
            .I3(n39709), .O(n40594));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34272_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33647_3_lut (.I0(n40498), .I1(n85), .I2(n41_adj_4427), .I3(GND_net), 
            .O(n39969));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33647_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13651_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13950), .I3(GND_net), .O(n18158));   // verilog/coms.v(126[12] 289[6])
    defparam i13651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13652_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13950), .I3(GND_net), .O(n18159));   // verilog/coms.v(126[12] 289[6])
    defparam i13652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13653_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13950), .I3(GND_net), .O(n18160));   // verilog/coms.v(126[12] 289[6])
    defparam i13653_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_30 (.CI(n29213), 
            .I0(GND_net), .I1(n5_adj_4571), .CO(n29214));
    SB_CARRY communication_counter_31__I_0_add_916_8 (.CI(n28540), .I0(n1353), 
            .I1(VCC_net), .CO(n28541));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4572), .I3(n29212), .O(n6_adj_3979)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_78_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[12]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_107[12]), 
            .I2(n15), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY blue_1137_add_4_3 (.CI(n28306), .I0(GND_net), .I1(blue[1]), 
            .CO(n28307));
    SB_LUT4 blue_1137_add_4_2_lut (.I0(GND_net), .I1(color_23__N_34), .I2(blue[0]), 
            .I3(GND_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam blue_1137_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_29 (.CI(n29212), 
            .I0(GND_net), .I1(n6_adj_4572), .CO(n29213));
    SB_LUT4 communication_counter_31__I_0_add_916_7_lut (.I0(GND_net), .I1(n1354), 
            .I2(GND_net), .I3(n28539), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY blue_1137_add_4_2 (.CI(GND_net), .I0(color_23__N_34), .I1(blue[0]), 
            .CO(n28306));
    SB_CARRY add_3184_15 (.CI(n28108), .I0(n2709), .I1(n88), .CO(n28109));
    SB_CARRY communication_counter_31__I_0_add_916_7 (.CI(n28539), .I0(n1354), 
            .I1(GND_net), .CO(n28540));
    SB_LUT4 communication_counter_31__I_0_add_1586_22_lut (.I0(n2372_adj_4237), 
            .I1(n2339), .I2(VCC_net), .I3(n28305), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4573), .I3(n29211), .O(n7_adj_3978)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_916_6_lut (.I0(GND_net), .I1(n1355), 
            .I2(GND_net), .I3(n28538), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_21_lut (.I0(GND_net), .I1(n2340), 
            .I2(VCC_net), .I3(n28304), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3184_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n28107), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_9_lut (.I0(duty[7]), .I1(n41708), .I2(n18), .I3(n27574), 
            .O(pwm_setpoint_22__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_916_6 (.CI(n28538), .I0(n1355), 
            .I1(GND_net), .CO(n28539));
    SB_CARRY communication_counter_31__I_0_add_1586_21 (.CI(n28304), .I0(n2340), 
            .I1(VCC_net), .CO(n28305));
    SB_CARRY add_3184_14 (.CI(n28107), .I0(n2710), .I1(n89), .CO(n28108));
    SB_CARRY add_555_9 (.CI(n27574), .I0(n41708), .I1(n18), .CO(n27575));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_28 (.CI(n29211), 
            .I0(GND_net), .I1(n7_adj_4573), .CO(n29212));
    SB_LUT4 communication_counter_31__I_0_add_916_5_lut (.I0(GND_net), .I1(n1356), 
            .I2(VCC_net), .I3(n28537), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n27971), 
            .O(n6808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13861_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n33775), .I3(GND_net), .O(n18368));   // verilog/coms.v(126[12] 289[6])
    defparam i13861_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3178_14 (.CI(n27971), .I0(n2172), .I1(n88), .CO(n27972));
    SB_CARRY communication_counter_31__I_0_add_916_5 (.CI(n28537), .I0(n1356), 
            .I1(VCC_net), .CO(n28538));
    SB_LUT4 communication_counter_31__I_0_add_1586_20_lut (.I0(GND_net), .I1(n2341), 
            .I2(VCC_net), .I3(n28303), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_916_4_lut (.I0(GND_net), .I1(n1357), 
            .I2(VCC_net), .I3(n28536), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_4574), .I3(n29210), .O(n8_adj_3977)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_916_4 (.CI(n28536), .I0(n1357), 
            .I1(VCC_net), .CO(n28537));
    SB_LUT4 communication_counter_31__I_0_add_916_3_lut (.I0(GND_net), .I1(n1358), 
            .I2(GND_net), .I3(n28535), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_20 (.CI(n28303), .I0(n2341), 
            .I1(VCC_net), .CO(n28304));
    SB_LUT4 add_3184_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n28106), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_19_lut (.I0(GND_net), .I1(n2342), 
            .I2(VCC_net), .I3(n28302), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_13 (.CI(n28106), .I0(n2711), .I1(n90), .CO(n28107));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_27 (.CI(n29210), 
            .I0(GND_net), .I1(n8_adj_4574), .CO(n29211));
    SB_CARRY communication_counter_31__I_0_add_916_3 (.CI(n28535), .I0(n1358), 
            .I1(GND_net), .CO(n28536));
    SB_CARRY communication_counter_31__I_0_add_1586_19 (.CI(n28302), .I0(n2342), 
            .I1(VCC_net), .CO(n28303));
    SB_LUT4 add_3184_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n28105), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_8_lut (.I0(duty[6]), .I1(n41708), .I2(n19), .I3(n27573), 
            .O(pwm_setpoint_22__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3178_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n27970), 
            .O(n6809)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_916_2 (.CI(VCC_net), .I0(n1458), 
            .I1(VCC_net), .CO(n28535));
    SB_CARRY add_3184_12 (.CI(n28105), .I0(n2712), .I1(n91), .CO(n28106));
    SB_LUT4 communication_counter_31__I_0_add_983_13_lut (.I0(n1481), .I1(n1448), 
            .I2(VCC_net), .I3(n28534), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_4575), .I3(n29209), .O(n9_adj_3976)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_26 (.CI(n29209), 
            .I0(GND_net), .I1(n9_adj_4575), .CO(n29210));
    SB_CARRY add_3178_13 (.CI(n27970), .I0(n2173), .I1(n89), .CO(n27971));
    SB_CARRY add_555_8 (.CI(n27573), .I0(n41708), .I1(n19), .CO(n27574));
    SB_LUT4 add_3184_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n28104), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_4576), .I3(n29208), .O(n10_adj_3975)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_18_lut (.I0(GND_net), .I1(n2343), 
            .I2(VCC_net), .I3(n28301), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_25 (.CI(n29208), 
            .I0(GND_net), .I1(n10_adj_4576), .CO(n29209));
    SB_LUT4 communication_counter_31__I_0_add_983_12_lut (.I0(GND_net), .I1(n1449), 
            .I2(VCC_net), .I3(n28533), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_18 (.CI(n28301), .I0(n2343), 
            .I1(VCC_net), .CO(n28302));
    SB_CARRY add_3184_11 (.CI(n28104), .I0(n2713), .I1(n92), .CO(n28105));
    SB_LUT4 communication_counter_31__I_0_add_1586_17_lut (.I0(GND_net), .I1(n2344), 
            .I2(VCC_net), .I3(n28300), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_4577), .I3(n29207), .O(n11_adj_3974)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_12 (.CI(n28533), .I0(n1449), 
            .I1(VCC_net), .CO(n28534));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_24 (.CI(n29207), 
            .I0(GND_net), .I1(n11_adj_4577), .CO(n29208));
    SB_CARRY communication_counter_31__I_0_add_1586_17 (.CI(n28300), .I0(n2344), 
            .I1(VCC_net), .CO(n28301));
    SB_LUT4 communication_counter_31__I_0_add_1586_16_lut (.I0(GND_net), .I1(n2345), 
            .I2(VCC_net), .I3(n28299), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_983_11_lut (.I0(GND_net), .I1(n1450), 
            .I2(VCC_net), .I3(n28532), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n27969), 
            .O(n6810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_11 (.CI(n28532), .I0(n1450), 
            .I1(VCC_net), .CO(n28533));
    SB_CARRY add_3178_12 (.CI(n27969), .I0(n2174), .I1(n90), .CO(n27970));
    SB_LUT4 communication_counter_31__I_0_add_983_10_lut (.I0(GND_net), .I1(n1451), 
            .I2(VCC_net), .I3(n28531), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_16 (.CI(n28299), .I0(n2345), 
            .I1(VCC_net), .CO(n28300));
    SB_LUT4 add_3178_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n27968), 
            .O(n6811)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_15_lut (.I0(GND_net), .I1(n2346_adj_4240), 
            .I2(VCC_net), .I3(n28298), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_10 (.CI(n28531), .I0(n1451), 
            .I1(VCC_net), .CO(n28532));
    SB_LUT4 add_555_7_lut (.I0(duty[5]), .I1(n41708), .I2(n20), .I3(n27572), 
            .O(pwm_setpoint_22__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3184_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n28103), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_15 (.CI(n28298), .I0(n2346_adj_4240), 
            .I1(VCC_net), .CO(n28299));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_4578), .I3(n29206), .O(n12_adj_3973)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_983_9_lut (.I0(GND_net), .I1(n1452), 
            .I2(VCC_net), .I3(n28530), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_14_lut (.I0(GND_net), .I1(n2347), 
            .I2(VCC_net), .I3(n28297), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_9 (.CI(n28530), .I0(n1452), 
            .I1(VCC_net), .CO(n28531));
    SB_CARRY communication_counter_31__I_0_add_1586_14 (.CI(n28297), .I0(n2347), 
            .I1(VCC_net), .CO(n28298));
    SB_CARRY add_3184_10 (.CI(n28103), .I0(n2714), .I1(n93), .CO(n28104));
    SB_LUT4 add_3184_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n28102), 
            .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_7 (.CI(n27572), .I0(n41708), .I1(n20), .CO(n27573));
    SB_CARRY add_3178_11 (.CI(n27968), .I0(n2175), .I1(n91), .CO(n27969));
    SB_LUT4 add_3178_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n27967), 
            .O(n6812)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_10 (.CI(n27967), .I0(n2176), .I1(n92), .CO(n27968));
    SB_LUT4 add_3178_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n27966), 
            .O(n6813)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_9 (.CI(n28102), .I0(n2715), .I1(n94), .CO(n28103));
    SB_CARRY add_3178_9 (.CI(n27966), .I0(n2177), .I1(n93), .CO(n27967));
    SB_LUT4 add_3178_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n27965), 
            .O(n6814)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_8 (.CI(n27965), .I0(n2178), .I1(n94), .CO(n27966));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_23 (.CI(n29206), 
            .I0(GND_net), .I1(n12_adj_4578), .CO(n29207));
    SB_LUT4 communication_counter_31__I_0_add_983_8_lut (.I0(GND_net), .I1(n1453), 
            .I2(VCC_net), .I3(n28529), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_13_lut (.I0(GND_net), .I1(n2348), 
            .I2(VCC_net), .I3(n28296), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_4579), .I3(n29205), .O(n13_adj_3972)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_8 (.CI(n28529), .I0(n1453), 
            .I1(VCC_net), .CO(n28530));
    SB_CARRY communication_counter_31__I_0_add_1586_13 (.CI(n28296), .I0(n2348), 
            .I1(VCC_net), .CO(n28297));
    SB_LUT4 add_3184_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n28101), 
            .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_12_lut (.I0(GND_net), .I1(n2349), 
            .I2(VCC_net), .I3(n28295), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_983_7_lut (.I0(GND_net), .I1(n1454), 
            .I2(GND_net), .I3(n28528), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_22 (.CI(n29205), 
            .I0(GND_net), .I1(n13_adj_4579), .CO(n29206));
    SB_CARRY communication_counter_31__I_0_add_983_7 (.CI(n28528), .I0(n1454), 
            .I1(GND_net), .CO(n28529));
    SB_CARRY communication_counter_31__I_0_add_1586_12 (.CI(n28295), .I0(n2349), 
            .I1(VCC_net), .CO(n28296));
    SB_LUT4 communication_counter_31__I_0_add_983_6_lut (.I0(GND_net), .I1(n1455), 
            .I2(GND_net), .I3(n28527), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_4580), .I3(n29204), .O(n14_adj_3971)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_6 (.CI(n28527), .I0(n1455), 
            .I1(GND_net), .CO(n28528));
    SB_LUT4 communication_counter_31__I_0_add_1586_11_lut (.I0(GND_net), .I1(n2350), 
            .I2(VCC_net), .I3(n28294), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_8 (.CI(n28101), .I0(n2716), .I1(n95), .CO(n28102));
    SB_CARRY communication_counter_31__I_0_add_1586_11 (.CI(n28294), .I0(n2350), 
            .I1(VCC_net), .CO(n28295));
    SB_LUT4 communication_counter_31__I_0_add_983_5_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n28526), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_21 (.CI(n29204), 
            .I0(GND_net), .I1(n14_adj_4580), .CO(n29205));
    SB_CARRY communication_counter_31__I_0_add_983_5 (.CI(n28526), .I0(n1456), 
            .I1(VCC_net), .CO(n28527));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_4581), .I3(n29203), .O(n15_adj_3970)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_983_4_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n28525), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_10_lut (.I0(GND_net), .I1(n2351), 
            .I2(VCC_net), .I3(n28293), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_20 (.CI(n29203), 
            .I0(GND_net), .I1(n15_adj_4581), .CO(n29204));
    SB_CARRY communication_counter_31__I_0_add_983_4 (.CI(n28525), .I0(n1457), 
            .I1(VCC_net), .CO(n28526));
    SB_CARRY communication_counter_31__I_0_add_1586_10 (.CI(n28293), .I0(n2351), 
            .I1(VCC_net), .CO(n28294));
    SB_LUT4 add_3184_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n28100), 
            .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_4582), .I3(n29202), .O(n16_adj_3969)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_983_3_lut (.I0(GND_net), .I1(n1458), 
            .I2(GND_net), .I3(n28524), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_9_lut (.I0(GND_net), .I1(n2352), 
            .I2(VCC_net), .I3(n28292), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_983_3 (.CI(n28524), .I0(n1458), 
            .I1(GND_net), .CO(n28525));
    SB_CARRY add_3184_7 (.CI(n28100), .I0(n2717), .I1(n96), .CO(n28101));
    SB_LUT4 add_555_6_lut (.I0(duty[4]), .I1(n41708), .I2(n21), .I3(n27571), 
            .O(pwm_setpoint_22__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_1586_9 (.CI(n28292), .I0(n2352), 
            .I1(VCC_net), .CO(n28293));
    SB_LUT4 add_3184_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n28099), 
            .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_19 (.CI(n29202), 
            .I0(GND_net), .I1(n16_adj_4582), .CO(n29203));
    SB_CARRY communication_counter_31__I_0_add_983_2 (.CI(VCC_net), .I0(n1558), 
            .I1(VCC_net), .CO(n28524));
    SB_LUT4 communication_counter_31__I_0_add_1586_8_lut (.I0(GND_net), .I1(n2353), 
            .I2(VCC_net), .I3(n28291), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_4583), .I3(n29201), .O(n17_adj_3968)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_14_lut (.I0(n1580), .I1(n1547), 
            .I2(VCC_net), .I3(n28523), .O(n1646_adj_4121)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_1050_13_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n28522), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_8 (.CI(n28291), .I0(n2353), 
            .I1(VCC_net), .CO(n28292));
    SB_CARRY add_3184_6 (.CI(n28099), .I0(n2718), .I1(n97), .CO(n28100));
    SB_LUT4 communication_counter_31__I_0_add_1586_7_lut (.I0(GND_net), .I1(n2354), 
            .I2(GND_net), .I3(n28290), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3184_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n28098), 
            .O(n6953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_5 (.CI(n28098), .I0(n2719), .I1(n98), .CO(n28099));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_18 (.CI(n29201), 
            .I0(GND_net), .I1(n17_adj_4583), .CO(n29202));
    SB_CARRY communication_counter_31__I_0_add_1050_13 (.CI(n28522), .I0(n1548), 
            .I1(VCC_net), .CO(n28523));
    SB_CARRY communication_counter_31__I_0_add_1586_7 (.CI(n28290), .I0(n2354), 
            .I1(GND_net), .CO(n28291));
    SB_LUT4 communication_counter_31__I_0_add_1050_12_lut (.I0(GND_net), .I1(n1549), 
            .I2(VCC_net), .I3(n28521), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_4584), .I3(n29200), .O(n18_adj_3967)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_12 (.CI(n28521), .I0(n1549), 
            .I1(VCC_net), .CO(n28522));
    SB_LUT4 communication_counter_31__I_0_add_1586_6_lut (.I0(GND_net), .I1(n2355), 
            .I2(GND_net), .I3(n28289), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3184_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n28097), 
            .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_6 (.CI(n28289), .I0(n2355), 
            .I1(GND_net), .CO(n28290));
    SB_LUT4 communication_counter_31__I_0_add_1050_11_lut (.I0(GND_net), .I1(n1550), 
            .I2(VCC_net), .I3(n28520), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_5_lut (.I0(GND_net), .I1(n2356), 
            .I2(VCC_net), .I3(n28288), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3184_4 (.CI(n28097), .I0(n2720), .I1(n99), .CO(n28098));
    SB_CARRY communication_counter_31__I_0_add_1586_5 (.CI(n28288), .I0(n2356), 
            .I1(VCC_net), .CO(n28289));
    SB_CARRY communication_counter_31__I_0_add_1050_11 (.CI(n28520), .I0(n1550), 
            .I1(VCC_net), .CO(n28521));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_17 (.CI(n29200), 
            .I0(GND_net), .I1(n18_adj_4584), .CO(n29201));
    SB_LUT4 communication_counter_31__I_0_add_1050_10_lut (.I0(GND_net), .I1(n1551), 
            .I2(VCC_net), .I3(n28519), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_4585), .I3(n29199), .O(n19_adj_3966)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1717_3_lut_3_lut (.I0(n2558), .I1(n6904), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3178_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n27964), 
            .O(n6815)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_7 (.CI(n27964), .I0(n2179), .I1(n95), .CO(n27965));
    SB_CARRY communication_counter_31__I_0_add_1050_10 (.CI(n28519), .I0(n1551), 
            .I1(VCC_net), .CO(n28520));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_16 (.CI(n29199), 
            .I0(GND_net), .I1(n19_adj_4585), .CO(n29200));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_4586), .I3(n29198), .O(n20_adj_3965)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_15 (.CI(n29198), 
            .I0(GND_net), .I1(n20_adj_4586), .CO(n29199));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_4587), .I3(n29197), .O(n21_adj_3964)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_14 (.CI(n29197), 
            .I0(GND_net), .I1(n21_adj_4587), .CO(n29198));
    SB_CARRY add_555_6 (.CI(n27571), .I0(n41708), .I1(n21), .CO(n27572));
    SB_LUT4 communication_counter_31__I_0_add_1050_9_lut (.I0(GND_net), .I1(n1552), 
            .I2(VCC_net), .I3(n28518), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4239), 
            .I2(VCC_net), .I3(n28287), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n27963), 
            .O(n6816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_9 (.CI(n28518), .I0(n1552), 
            .I1(VCC_net), .CO(n28519));
    SB_LUT4 add_3184_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n28096), 
            .O(n6955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3184_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_4 (.CI(n28287), .I0(n2357_adj_4239), 
            .I1(VCC_net), .CO(n28288));
    SB_LUT4 communication_counter_31__I_0_add_1050_8_lut (.I0(GND_net), .I1(n1553_adj_4130), 
            .I2(VCC_net), .I3(n28517), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_6 (.CI(n27963), .I0(n2180), .I1(n96), .CO(n27964));
    SB_LUT4 add_555_5_lut (.I0(duty[3]), .I1(n41708), .I2(n22), .I3(n27570), 
            .O(pwm_setpoint_22__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3184_3 (.CI(n28096), .I0(n390), .I1(n558), .CO(n28097));
    SB_LUT4 add_3178_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n27962), 
            .O(n6817)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4238), 
            .I2(GND_net), .I3(n28286), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1586_3 (.CI(n28286), .I0(n2358_adj_4238), 
            .I1(GND_net), .CO(n28287));
    SB_CARRY communication_counter_31__I_0_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4225), 
            .I1(VCC_net), .CO(n28286));
    SB_LUT4 communication_counter_1136_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n28285), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_8 (.CI(n28517), .I0(n1553_adj_4130), 
            .I1(VCC_net), .CO(n28518));
    SB_CARRY add_3184_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n28096));
    SB_CARRY add_3178_5 (.CI(n27962), .I0(n2181), .I1(n97), .CO(n27963));
    SB_LUT4 communication_counter_1136_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n28284), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_7_lut (.I0(GND_net), .I1(n1554_adj_4131), 
            .I2(GND_net), .I3(n28516), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13654_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13950), .I3(GND_net), .O(n18161));   // verilog/coms.v(126[12] 289[6])
    defparam i13654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13655_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13950), .I3(GND_net), .O(n18162));   // verilog/coms.v(126[12] 289[6])
    defparam i13655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1714_3_lut_3_lut (.I0(n2558), .I1(n6901), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4218));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_78_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[13]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_107[13]), 
            .I2(n15), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3931));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4199));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_78_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[14]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_107[14]), 
            .I2(n15), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13656_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13950), .I3(GND_net), .O(n18163));   // verilog/coms.v(126[12] 289[6])
    defparam i13656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13657_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13950), .I3(GND_net), .O(n18164));   // verilog/coms.v(126[12] 289[6])
    defparam i13657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13658_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13950), .I3(GND_net), .O(n18165));   // verilog/coms.v(126[12] 289[6])
    defparam i13658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13659_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13950), .I3(GND_net), .O(n18166));   // verilog/coms.v(126[12] 289[6])
    defparam i13659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4198));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_78_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[15]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_107[15]), 
            .I2(n15), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4197));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13660_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13950), .I3(GND_net), .O(n18167));   // verilog/coms.v(126[12] 289[6])
    defparam i13660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13661_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13950), .I3(GND_net), .O(n18168));   // verilog/coms.v(126[12] 289[6])
    defparam i13661_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1136_add_4_32 (.CI(n28284), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n28285));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_4588), .I3(n29196), .O(n22_adj_3963)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13662_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13950), .I3(GND_net), .O(n18169));   // verilog/coms.v(126[12] 289[6])
    defparam i13662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4196));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13663_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13950), .I3(GND_net), .O(n18170));   // verilog/coms.v(126[12] 289[6])
    defparam i13663_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_13 (.CI(n29196), 
            .I0(GND_net), .I1(n22_adj_4588), .CO(n29197));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_4589), .I3(n29195), .O(n23_adj_3962)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_12 (.CI(n29195), 
            .I0(GND_net), .I1(n23_adj_4589), .CO(n29196));
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_1050_7 (.CI(n28516), .I0(n1554_adj_4131), 
            .I1(GND_net), .CO(n28517));
    SB_LUT4 mux_78_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[16]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_107[16]), 
            .I2(n15), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_4590), .I3(n29194), .O(n24_adj_3961)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1589_3_lut (.I0(n2363), .I1(n6849), .I2(n2381), .I3(GND_net), 
            .O(n2453));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_11 (.CI(n29194), 
            .I0(GND_net), .I1(n24_adj_4590), .CO(n29195));
    SB_LUT4 add_3178_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n27961), 
            .O(n6818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_78_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[17]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3178_4 (.CI(n27961), .I0(n2182), .I1(n98), .CO(n27962));
    SB_LUT4 mux_77_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_107[17]), 
            .I2(n15), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3178_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n27960), 
            .O(n6819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_3 (.CI(n27960), .I0(n2183), .I1(n99), .CO(n27961));
    SB_LUT4 add_3178_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n27960));
    SB_LUT4 add_3177_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n27959), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3177_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n27958), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_16 (.CI(n27958), .I0(n2070), .I1(n86), .CO(n27959));
    SB_LUT4 add_3177_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n27957), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_6_lut (.I0(GND_net), .I1(n1555), 
            .I2(GND_net), .I3(n28515), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n28283), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n28095), 
            .O(n6909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_4591), .I3(n29193), .O(n25_adj_3960)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_6 (.CI(n28515), .I0(n1555), 
            .I1(GND_net), .CO(n28516));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_10 (.CI(n29193), 
            .I0(GND_net), .I1(n25_adj_4591), .CO(n29194));
    SB_CARRY communication_counter_1136_add_4_31 (.CI(n28283), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n28284));
    SB_LUT4 div_46_i1707_3_lut_3_lut (.I0(n2558), .I1(n6894), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_78_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[18]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3177_15 (.CI(n27957), .I0(n2071), .I1(n87), .CO(n27958));
    SB_LUT4 mux_77_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_107[18]), 
            .I2(n15), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1136_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n28282), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n28094), 
            .O(n6910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3177_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n27956), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_14 (.CI(n27956), .I0(n2072), .I1(n88), .CO(n27957));
    SB_LUT4 add_3177_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n27955), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_13 (.CI(n27955), .I0(n2073), .I1(n89), .CO(n27956));
    SB_LUT4 add_3177_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n27954), 
            .O(n6791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_12 (.CI(n27954), .I0(n2074), .I1(n90), .CO(n27955));
    SB_LUT4 add_3177_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n27953), 
            .O(n6792)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_11 (.CI(n27953), .I0(n2075), .I1(n91), .CO(n27954));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_4592), .I3(n29192), .O(n26_adj_3959)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_22 (.CI(n28094), .I0(n2619), .I1(n80), .CO(n28095));
    SB_CARRY communication_counter_1136_add_4_30 (.CI(n28282), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n28283));
    SB_LUT4 add_3177_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n27952), 
            .O(n6793)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n28093), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n28281), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_5_lut (.I0(GND_net), .I1(n1556), 
            .I2(VCC_net), .I3(n28514), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_5 (.CI(n28514), .I0(n1556), 
            .I1(VCC_net), .CO(n28515));
    SB_CARRY add_3177_10 (.CI(n27952), .I0(n2076), .I1(n92), .CO(n27953));
    SB_CARRY add_3183_21 (.CI(n28093), .I0(n2620), .I1(n81), .CO(n28094));
    SB_CARRY communication_counter_1136_add_4_29 (.CI(n28281), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n28282));
    SB_LUT4 add_3177_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n27951), 
            .O(n6794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_9 (.CI(n27951), .I0(n2077), .I1(n93), .CO(n27952));
    SB_LUT4 add_3183_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n28092), 
            .O(n6912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n28280), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_4_lut (.I0(GND_net), .I1(n1557), 
            .I2(VCC_net), .I3(n28513), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_9 (.CI(n29192), 
            .I0(GND_net), .I1(n26_adj_4592), .CO(n29193));
    SB_CARRY communication_counter_31__I_0_add_1050_4 (.CI(n28513), .I0(n1557), 
            .I1(VCC_net), .CO(n28514));
    SB_LUT4 add_3177_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n27950), 
            .O(n6795)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_8 (.CI(n27950), .I0(n2078), .I1(n94), .CO(n27951));
    SB_LUT4 add_3177_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n27949), 
            .O(n6796)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_7 (.CI(n27949), .I0(n2079), .I1(n95), .CO(n27950));
    SB_LUT4 add_3177_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n27948), 
            .O(n6797)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_6 (.CI(n27948), .I0(n2080), .I1(n96), .CO(n27949));
    SB_LUT4 add_3177_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n27947), 
            .O(n6798)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_5 (.CI(n27947), .I0(n2081), .I1(n97), .CO(n27948));
    SB_LUT4 add_3177_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n27946), 
            .O(n6799)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_4 (.CI(n27946), .I0(n2082), .I1(n98), .CO(n27947));
    SB_LUT4 add_3177_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n27945), 
            .O(n6800)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_3 (.CI(n27945), .I0(n2083), .I1(n99), .CO(n27946));
    SB_LUT4 add_3177_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6801)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3177_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3177_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n27945));
    SB_LUT4 communication_counter_31__I_0_add_2055_28_lut (.I0(n3065), .I1(n3032), 
            .I2(VCC_net), .I3(n27944), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_2055_27_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n27943), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_27 (.CI(n27943), .I0(n3033), 
            .I1(VCC_net), .CO(n27944));
    SB_LUT4 communication_counter_31__I_0_add_2055_26_lut (.I0(GND_net), .I1(n3034), 
            .I2(VCC_net), .I3(n27942), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_26 (.CI(n27942), .I0(n3034), 
            .I1(VCC_net), .CO(n27943));
    SB_LUT4 communication_counter_31__I_0_add_2055_25_lut (.I0(GND_net), .I1(n3035), 
            .I2(VCC_net), .I3(n27941), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_25 (.CI(n27941), .I0(n3035), 
            .I1(VCC_net), .CO(n27942));
    SB_LUT4 communication_counter_31__I_0_add_2055_24_lut (.I0(GND_net), .I1(n3036), 
            .I2(VCC_net), .I3(n27940), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_24 (.CI(n27940), .I0(n3036), 
            .I1(VCC_net), .CO(n27941));
    SB_LUT4 communication_counter_31__I_0_add_2055_23_lut (.I0(GND_net), .I1(n3037), 
            .I2(VCC_net), .I3(n27939), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_23 (.CI(n27939), .I0(n3037), 
            .I1(VCC_net), .CO(n27940));
    SB_LUT4 communication_counter_31__I_0_add_2055_22_lut (.I0(GND_net), .I1(n3038), 
            .I2(VCC_net), .I3(n27938), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_22 (.CI(n27938), .I0(n3038), 
            .I1(VCC_net), .CO(n27939));
    SB_LUT4 communication_counter_31__I_0_add_2055_21_lut (.I0(GND_net), .I1(n3039), 
            .I2(VCC_net), .I3(n27937), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_21 (.CI(n27937), .I0(n3039), 
            .I1(VCC_net), .CO(n27938));
    SB_LUT4 communication_counter_31__I_0_add_2055_20_lut (.I0(GND_net), .I1(n3040), 
            .I2(VCC_net), .I3(n27936), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_20 (.CI(n27936), .I0(n3040), 
            .I1(VCC_net), .CO(n27937));
    SB_LUT4 mux_78_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[19]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_107[19]), 
            .I2(n15), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_4593), .I3(n29191), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_28 (.CI(n28280), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n28281));
    SB_CARRY add_555_5 (.CI(n27570), .I0(n41708), .I1(n22), .CO(n27571));
    SB_LUT4 communication_counter_31__I_0_add_2055_19_lut (.I0(GND_net), .I1(n3041), 
            .I2(VCC_net), .I3(n27935), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_20 (.CI(n28092), .I0(n2621), .I1(n82), .CO(n28093));
    SB_LUT4 communication_counter_1136_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n28279), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1050_3_lut (.I0(GND_net), .I1(n1558), 
            .I2(GND_net), .I3(n28512), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_19 (.CI(n27935), .I0(n3041), 
            .I1(VCC_net), .CO(n27936));
    SB_LUT4 communication_counter_31__I_0_add_2055_18_lut (.I0(GND_net), .I1(n3042), 
            .I2(VCC_net), .I3(n27934), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1050_3 (.CI(n28512), .I0(n1558), 
            .I1(GND_net), .CO(n28513));
    SB_CARRY communication_counter_31__I_0_add_1050_2 (.CI(VCC_net), .I0(n1658), 
            .I1(VCC_net), .CO(n28512));
    SB_LUT4 communication_counter_31__I_0_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4121), 
            .I2(VCC_net), .I3(n28511), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_DFF communication_counter_1136__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_LUT4 div_46_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_3992), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1539_3_lut (.I0(n385), .I1(n6840), .I2(n2288), .I3(GND_net), 
            .O(n2374));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1539_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13664_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13950), .I3(GND_net), .O(n18171));   // verilog/coms.v(126[12] 289[6])
    defparam i13664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[20]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_107[20]), 
            .I2(n15), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4195));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_2055_18 (.CI(n27934), .I0(n3042), 
            .I1(VCC_net), .CO(n27935));
    SB_LUT4 i13665_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13950), .I3(GND_net), .O(n18172));   // verilog/coms.v(126[12] 289[6])
    defparam i13665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13666_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13950), .I3(GND_net), .O(n18173));   // verilog/coms.v(126[12] 289[6])
    defparam i13666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[21]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_107[21]), 
            .I2(n15), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13667_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13950), .I3(GND_net), .O(n18174));   // verilog/coms.v(126[12] 289[6])
    defparam i13667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_2055_17_lut (.I0(GND_net), .I1(n3043), 
            .I2(VCC_net), .I3(n27933), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_17 (.CI(n27933), .I0(n3043), 
            .I1(VCC_net), .CO(n27934));
    SB_LUT4 communication_counter_31__I_0_add_2055_16_lut (.I0(GND_net), .I1(n3044), 
            .I2(VCC_net), .I3(n27932), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_16 (.CI(n27932), .I0(n3044), 
            .I1(VCC_net), .CO(n27933));
    SB_LUT4 communication_counter_31__I_0_add_2055_15_lut (.I0(GND_net), .I1(n3045), 
            .I2(VCC_net), .I3(n27931), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_15 (.CI(n27931), .I0(n3045), 
            .I1(VCC_net), .CO(n27932));
    SB_LUT4 communication_counter_31__I_0_add_2055_14_lut (.I0(GND_net), .I1(n3046), 
            .I2(VCC_net), .I3(n27930), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_14 (.CI(n27930), .I0(n3046), 
            .I1(VCC_net), .CO(n27931));
    SB_LUT4 communication_counter_31__I_0_add_2055_13_lut (.I0(GND_net), .I1(n3047), 
            .I2(VCC_net), .I3(n27929), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_13 (.CI(n27929), .I0(n3047), 
            .I1(VCC_net), .CO(n27930));
    SB_LUT4 communication_counter_31__I_0_add_2055_12_lut (.I0(GND_net), .I1(n3048), 
            .I2(VCC_net), .I3(n27928), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_12 (.CI(n27928), .I0(n3048), 
            .I1(VCC_net), .CO(n27929));
    SB_LUT4 communication_counter_31__I_0_add_2055_11_lut (.I0(GND_net), .I1(n3049), 
            .I2(VCC_net), .I3(n27927), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_11 (.CI(n27927), .I0(n3049), 
            .I1(VCC_net), .CO(n27928));
    SB_LUT4 communication_counter_31__I_0_add_2055_10_lut (.I0(GND_net), .I1(n3050), 
            .I2(VCC_net), .I3(n27926), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_10 (.CI(n27926), .I0(n3050), 
            .I1(VCC_net), .CO(n27927));
    SB_LUT4 communication_counter_31__I_0_add_2055_9_lut (.I0(GND_net), .I1(n3051), 
            .I2(VCC_net), .I3(n27925), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_9 (.CI(n27925), .I0(n3051), 
            .I1(VCC_net), .CO(n27926));
    SB_LUT4 communication_counter_31__I_0_add_2055_8_lut (.I0(GND_net), .I1(n3052), 
            .I2(VCC_net), .I3(n27924), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_8 (.CI(n27924), .I0(n3052), 
            .I1(VCC_net), .CO(n27925));
    SB_LUT4 communication_counter_31__I_0_add_2055_7_lut (.I0(GND_net), .I1(n3053), 
            .I2(VCC_net), .I3(n27923), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_7 (.CI(n27923), .I0(n3053), 
            .I1(VCC_net), .CO(n27924));
    SB_LUT4 communication_counter_31__I_0_add_2055_6_lut (.I0(GND_net), .I1(n3054), 
            .I2(GND_net), .I3(n27922), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_27 (.CI(n28279), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n28280));
    SB_LUT4 i13668_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13950), .I3(GND_net), .O(n18175));   // verilog/coms.v(126[12] 289[6])
    defparam i13668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3183_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n28091), 
            .O(n6913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_6 (.CI(n27922), .I0(n3054), 
            .I1(GND_net), .CO(n27923));
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3183_19 (.CI(n28091), .I0(n2622), .I1(n83), .CO(n28092));
    SB_LUT4 i13669_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13950), .I3(GND_net), .O(n18176));   // verilog/coms.v(126[12] 289[6])
    defparam i13669_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_8 (.CI(n29191), 
            .I0(GND_net), .I1(n27_adj_4593), .CO(n29192));
    SB_LUT4 communication_counter_31__I_0_add_2055_5_lut (.I0(GND_net), .I1(n3055), 
            .I2(GND_net), .I3(n27921), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4122), 
            .I2(VCC_net), .I3(n28510), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_5 (.CI(n27921), .I0(n3055), 
            .I1(GND_net), .CO(n27922));
    SB_LUT4 communication_counter_31__I_0_add_2055_4_lut (.I0(GND_net), .I1(n3056), 
            .I2(VCC_net), .I3(n27920), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_4 (.CI(n27920), .I0(n3056), 
            .I1(VCC_net), .CO(n27921));
    SB_LUT4 communication_counter_31__I_0_add_2055_3_lut (.I0(GND_net), .I1(n3057), 
            .I2(VCC_net), .I3(n27919), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_3 (.CI(n27919), .I0(n3057), 
            .I1(VCC_net), .CO(n27920));
    SB_LUT4 communication_counter_31__I_0_add_2055_2_lut (.I0(GND_net), .I1(n3058), 
            .I2(GND_net), .I3(VCC_net), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2055_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2055_2 (.CI(VCC_net), .I0(n3058), 
            .I1(GND_net), .CO(n27919));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_4594), .I3(n29190), .O(n28_adj_3958)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13670_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13950), .I3(GND_net), .O(n18177));   // verilog/coms.v(126[12] 289[6])
    defparam i13670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4194));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13671_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13950), .I3(GND_net), .O(n18178));   // verilog/coms.v(126[12] 289[6])
    defparam i13671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4193));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3176_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n27918), 
            .O(n6769)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n27917), 
            .O(n6770)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_15 (.CI(n27917), .I0(n1968), .I1(n87), .CO(n27918));
    SB_LUT4 add_3176_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n27916), 
            .O(n6771)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_14 (.CI(n27916), .I0(n1969), .I1(n88), .CO(n27917));
    SB_LUT4 add_3176_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n27915), 
            .O(n6772)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_13 (.CI(n27915), .I0(n1970), .I1(n89), .CO(n27916));
    SB_LUT4 add_3176_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n27914), 
            .O(n6773)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_12 (.CI(n27914), .I0(n1971), .I1(n90), .CO(n27915));
    SB_LUT4 add_3176_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n27913), 
            .O(n6774)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_11 (.CI(n27913), .I0(n1972), .I1(n91), .CO(n27914));
    SB_LUT4 add_3176_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n27912), 
            .O(n6775)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_10 (.CI(n27912), .I0(n1973), .I1(n92), .CO(n27913));
    SB_LUT4 add_3176_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n27911), 
            .O(n6776)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_9 (.CI(n27911), .I0(n1974), .I1(n93), .CO(n27912));
    SB_LUT4 add_3176_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n27910), 
            .O(n6777)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_8 (.CI(n27910), .I0(n1975), .I1(n94), .CO(n27911));
    SB_LUT4 add_3176_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n27909), 
            .O(n6778)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_7 (.CI(n27909), .I0(n1976), .I1(n95), .CO(n27910));
    SB_LUT4 add_3176_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n27908), 
            .O(n6779)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_6 (.CI(n27908), .I0(n1977), .I1(n96), .CO(n27909));
    SB_LUT4 add_3176_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n27907), 
            .O(n6780)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_5 (.CI(n27907), .I0(n1978), .I1(n97), .CO(n27908));
    SB_LUT4 add_3176_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n27906), 
            .O(n6781)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_4 (.CI(n27906), .I0(n1979), .I1(n98), .CO(n27907));
    SB_LUT4 add_3176_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n27905), 
            .O(n6782)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_3 (.CI(n27905), .I0(n1980), .I1(n99), .CO(n27906));
    SB_LUT4 add_3176_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6783)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n27905));
    SB_LUT4 add_3175_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n27904), 
            .O(n6753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3175_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n27903), 
            .O(n6754)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_14 (.CI(n27903), .I0(n1863), .I1(n88), .CO(n27904));
    SB_LUT4 add_3175_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n27902), 
            .O(n6755)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_13 (.CI(n27902), .I0(n1864), .I1(n89), .CO(n27903));
    SB_LUT4 add_3175_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n27901), 
            .O(n6756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_12 (.CI(n27901), .I0(n1865), .I1(n90), .CO(n27902));
    SB_LUT4 add_3175_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n27900), 
            .O(n6757)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_11 (.CI(n27900), .I0(n1866), .I1(n91), .CO(n27901));
    SB_LUT4 add_3175_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n27899), 
            .O(n6758)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_10 (.CI(n27899), .I0(n1867), .I1(n92), .CO(n27900));
    SB_LUT4 add_3175_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n27898), 
            .O(n6759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_9 (.CI(n27898), .I0(n1868), .I1(n93), .CO(n27899));
    SB_LUT4 add_3175_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n27897), 
            .O(n6760)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_8 (.CI(n27897), .I0(n1869), .I1(n94), .CO(n27898));
    SB_LUT4 add_3175_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n27896), 
            .O(n6761)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_7 (.CI(n27896), .I0(n1870), .I1(n95), .CO(n27897));
    SB_LUT4 add_3175_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n27895), 
            .O(n6762)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_6 (.CI(n27895), .I0(n1871), .I1(n96), .CO(n27896));
    SB_LUT4 add_3175_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n27894), 
            .O(n6763)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_5 (.CI(n27894), .I0(n1872), .I1(n97), .CO(n27895));
    SB_LUT4 add_3175_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n27893), 
            .O(n6764)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_4 (.CI(n27893), .I0(n1873), .I1(n98), .CO(n27894));
    SB_LUT4 add_3175_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n27892), 
            .O(n6765)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_3 (.CI(n27892), .I0(n1874), .I1(n99), .CO(n27893));
    SB_LUT4 add_3175_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6766)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3175_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3175_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n27892));
    SB_LUT4 communication_counter_31__I_0_add_2122_29_lut (.I0(n3164), .I1(n3131), 
            .I2(VCC_net), .I3(n27891), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_2122_28_lut (.I0(GND_net), .I1(n3132), 
            .I2(VCC_net), .I3(n27890), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_28 (.CI(n27890), .I0(n3132), 
            .I1(VCC_net), .CO(n27891));
    SB_LUT4 communication_counter_31__I_0_add_2122_27_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n27889), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_27 (.CI(n27889), .I0(n3133), 
            .I1(VCC_net), .CO(n27890));
    SB_LUT4 communication_counter_31__I_0_add_2122_26_lut (.I0(GND_net), .I1(n3134), 
            .I2(VCC_net), .I3(n27888), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_26 (.CI(n27888), .I0(n3134), 
            .I1(VCC_net), .CO(n27889));
    SB_LUT4 communication_counter_31__I_0_add_2122_25_lut (.I0(GND_net), .I1(n3135), 
            .I2(VCC_net), .I3(n27887), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_25 (.CI(n27887), .I0(n3135), 
            .I1(VCC_net), .CO(n27888));
    SB_LUT4 communication_counter_31__I_0_add_2122_24_lut (.I0(GND_net), .I1(n3136), 
            .I2(VCC_net), .I3(n27886), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_24 (.CI(n27886), .I0(n3136), 
            .I1(VCC_net), .CO(n27887));
    SB_LUT4 communication_counter_31__I_0_add_2122_23_lut (.I0(GND_net), .I1(n3137), 
            .I2(VCC_net), .I3(n27885), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_23 (.CI(n27885), .I0(n3137), 
            .I1(VCC_net), .CO(n27886));
    SB_LUT4 communication_counter_31__I_0_add_2122_22_lut (.I0(GND_net), .I1(n3138), 
            .I2(VCC_net), .I3(n27884), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_22 (.CI(n27884), .I0(n3138), 
            .I1(VCC_net), .CO(n27885));
    SB_LUT4 communication_counter_31__I_0_add_2122_21_lut (.I0(GND_net), .I1(n3139), 
            .I2(VCC_net), .I3(n27883), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_21 (.CI(n27883), .I0(n3139), 
            .I1(VCC_net), .CO(n27884));
    SB_LUT4 communication_counter_31__I_0_add_2122_20_lut (.I0(GND_net), .I1(n3140), 
            .I2(VCC_net), .I3(n27882), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_20 (.CI(n27882), .I0(n3140), 
            .I1(VCC_net), .CO(n27883));
    SB_LUT4 communication_counter_31__I_0_add_2122_19_lut (.I0(GND_net), .I1(n3141), 
            .I2(VCC_net), .I3(n27881), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_19 (.CI(n27881), .I0(n3141), 
            .I1(VCC_net), .CO(n27882));
    SB_LUT4 communication_counter_31__I_0_add_2122_18_lut (.I0(GND_net), .I1(n3142), 
            .I2(VCC_net), .I3(n27880), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_18 (.CI(n27880), .I0(n3142), 
            .I1(VCC_net), .CO(n27881));
    SB_LUT4 communication_counter_31__I_0_add_2122_17_lut (.I0(GND_net), .I1(n3143), 
            .I2(VCC_net), .I3(n27879), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_17 (.CI(n27879), .I0(n3143), 
            .I1(VCC_net), .CO(n27880));
    SB_LUT4 communication_counter_31__I_0_add_2122_16_lut (.I0(GND_net), .I1(n3144), 
            .I2(VCC_net), .I3(n27878), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_16 (.CI(n27878), .I0(n3144), 
            .I1(VCC_net), .CO(n27879));
    SB_LUT4 communication_counter_31__I_0_add_2122_15_lut (.I0(GND_net), .I1(n3145), 
            .I2(VCC_net), .I3(n27877), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_15 (.CI(n27877), .I0(n3145), 
            .I1(VCC_net), .CO(n27878));
    SB_LUT4 communication_counter_31__I_0_add_2122_14_lut (.I0(GND_net), .I1(n3146), 
            .I2(VCC_net), .I3(n27876), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_14 (.CI(n27876), .I0(n3146), 
            .I1(VCC_net), .CO(n27877));
    SB_LUT4 communication_counter_31__I_0_add_2122_13_lut (.I0(GND_net), .I1(n3147), 
            .I2(VCC_net), .I3(n27875), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_13 (.CI(n27875), .I0(n3147), 
            .I1(VCC_net), .CO(n27876));
    SB_LUT4 communication_counter_31__I_0_add_2122_12_lut (.I0(GND_net), .I1(n3148), 
            .I2(VCC_net), .I3(n27874), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_12 (.CI(n27874), .I0(n3148), 
            .I1(VCC_net), .CO(n27875));
    SB_LUT4 communication_counter_31__I_0_add_2122_11_lut (.I0(GND_net), .I1(n3149), 
            .I2(VCC_net), .I3(n27873), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_11 (.CI(n27873), .I0(n3149), 
            .I1(VCC_net), .CO(n27874));
    SB_LUT4 communication_counter_31__I_0_add_2122_10_lut (.I0(GND_net), .I1(n3150), 
            .I2(VCC_net), .I3(n27872), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_10 (.CI(n27872), .I0(n3150), 
            .I1(VCC_net), .CO(n27873));
    SB_LUT4 communication_counter_31__I_0_add_2122_9_lut (.I0(GND_net), .I1(n3151), 
            .I2(VCC_net), .I3(n27871), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_9 (.CI(n27871), .I0(n3151), 
            .I1(VCC_net), .CO(n27872));
    SB_LUT4 communication_counter_31__I_0_add_2122_8_lut (.I0(GND_net), .I1(n3152), 
            .I2(VCC_net), .I3(n27870), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_8 (.CI(n27870), .I0(n3152), 
            .I1(VCC_net), .CO(n27871));
    SB_LUT4 communication_counter_31__I_0_add_2122_7_lut (.I0(GND_net), .I1(n3153), 
            .I2(VCC_net), .I3(n27869), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_7 (.CI(n27869), .I0(n3153), 
            .I1(VCC_net), .CO(n27870));
    SB_LUT4 communication_counter_31__I_0_add_2122_6_lut (.I0(GND_net), .I1(n3154), 
            .I2(GND_net), .I3(n27868), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_6 (.CI(n27868), .I0(n3154), 
            .I1(GND_net), .CO(n27869));
    SB_LUT4 communication_counter_31__I_0_add_2122_5_lut (.I0(GND_net), .I1(n3155), 
            .I2(GND_net), .I3(n27867), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_5 (.CI(n27867), .I0(n3155), 
            .I1(GND_net), .CO(n27868));
    SB_LUT4 communication_counter_31__I_0_add_2122_4_lut (.I0(GND_net), .I1(n3156), 
            .I2(VCC_net), .I3(n27866), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_4 (.CI(n27866), .I0(n3156), 
            .I1(VCC_net), .CO(n27867));
    SB_LUT4 communication_counter_31__I_0_add_2122_3_lut (.I0(GND_net), .I1(n3157), 
            .I2(VCC_net), .I3(n27865), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_3 (.CI(n27865), .I0(n3157), 
            .I1(VCC_net), .CO(n27866));
    SB_LUT4 communication_counter_31__I_0_add_2122_2_lut (.I0(GND_net), .I1(n3158), 
            .I2(GND_net), .I3(VCC_net), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2122_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2122_2 (.CI(VCC_net), .I0(n3158), 
            .I1(GND_net), .CO(n27865));
    SB_LUT4 add_3174_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n27864), 
            .O(n6738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3174_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n27863), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_13 (.CI(n27863), .I0(n1755), .I1(n89), .CO(n27864));
    SB_LUT4 add_3174_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n27862), 
            .O(n6740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_12 (.CI(n27862), .I0(n1756), .I1(n90), .CO(n27863));
    SB_LUT4 add_3174_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n27861), 
            .O(n6741)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_11 (.CI(n27861), .I0(n1757), .I1(n91), .CO(n27862));
    SB_LUT4 add_3174_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n27860), 
            .O(n6742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_10 (.CI(n27860), .I0(n1758), .I1(n92), .CO(n27861));
    SB_LUT4 add_3174_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n27859), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_9 (.CI(n27859), .I0(n1759), .I1(n93), .CO(n27860));
    SB_LUT4 add_3174_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n27858), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_8 (.CI(n27858), .I0(n1760), .I1(n94), .CO(n27859));
    SB_LUT4 add_3174_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n27857), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_7 (.CI(n27857), .I0(n1761), .I1(n95), .CO(n27858));
    SB_LUT4 add_3174_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n27856), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_6 (.CI(n27856), .I0(n1762), .I1(n96), .CO(n27857));
    SB_LUT4 add_3174_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n27855), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_5 (.CI(n27855), .I0(n1763), .I1(n97), .CO(n27856));
    SB_LUT4 add_3174_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n27854), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_4 (.CI(n27854), .I0(n1764), .I1(n98), .CO(n27855));
    SB_LUT4 add_3174_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n27853), 
            .O(n6749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_3 (.CI(n27853), .I0(n1765), .I1(n99), .CO(n27854));
    SB_LUT4 add_3174_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3174_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3174_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n27853));
    SB_LUT4 communication_counter_31__I_0_add_2189_30_lut (.I0(n3263), .I1(n3230), 
            .I2(VCC_net), .I3(n27852), .O(n37078)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_2189_29_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n27851), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_29 (.CI(n27851), .I0(n3231), 
            .I1(VCC_net), .CO(n27852));
    SB_LUT4 communication_counter_31__I_0_add_2189_28_lut (.I0(GND_net), .I1(n3232), 
            .I2(VCC_net), .I3(n27850), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_28 (.CI(n27850), .I0(n3232), 
            .I1(VCC_net), .CO(n27851));
    SB_LUT4 communication_counter_31__I_0_add_2189_27_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n27849), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_27 (.CI(n27849), .I0(n3233), 
            .I1(VCC_net), .CO(n27850));
    SB_LUT4 communication_counter_31__I_0_add_2189_26_lut (.I0(GND_net), .I1(n3234), 
            .I2(VCC_net), .I3(n27848), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_26 (.CI(n27848), .I0(n3234), 
            .I1(VCC_net), .CO(n27849));
    SB_LUT4 communication_counter_31__I_0_add_2189_25_lut (.I0(GND_net), .I1(n3235), 
            .I2(VCC_net), .I3(n27847), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_25 (.CI(n27847), .I0(n3235), 
            .I1(VCC_net), .CO(n27848));
    SB_LUT4 communication_counter_31__I_0_add_2189_24_lut (.I0(GND_net), .I1(n3236), 
            .I2(VCC_net), .I3(n27846), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_24 (.CI(n27846), .I0(n3236), 
            .I1(VCC_net), .CO(n27847));
    SB_LUT4 communication_counter_31__I_0_add_2189_23_lut (.I0(GND_net), .I1(n3237), 
            .I2(VCC_net), .I3(n27845), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_23 (.CI(n27845), .I0(n3237), 
            .I1(VCC_net), .CO(n27846));
    SB_LUT4 communication_counter_31__I_0_add_2189_22_lut (.I0(GND_net), .I1(n3238), 
            .I2(VCC_net), .I3(n27844), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_22 (.CI(n27844), .I0(n3238), 
            .I1(VCC_net), .CO(n27845));
    SB_LUT4 communication_counter_31__I_0_add_2189_21_lut (.I0(GND_net), .I1(n3239), 
            .I2(VCC_net), .I3(n27843), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_21 (.CI(n27843), .I0(n3239), 
            .I1(VCC_net), .CO(n27844));
    SB_LUT4 communication_counter_31__I_0_add_2189_20_lut (.I0(GND_net), .I1(n3240), 
            .I2(VCC_net), .I3(n27842), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_20 (.CI(n27842), .I0(n3240), 
            .I1(VCC_net), .CO(n27843));
    SB_LUT4 communication_counter_31__I_0_add_2189_19_lut (.I0(GND_net), .I1(n3241), 
            .I2(VCC_net), .I3(n27841), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_19 (.CI(n27841), .I0(n3241), 
            .I1(VCC_net), .CO(n27842));
    SB_LUT4 communication_counter_31__I_0_add_2189_18_lut (.I0(GND_net), .I1(n3242), 
            .I2(VCC_net), .I3(n27840), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_18 (.CI(n27840), .I0(n3242), 
            .I1(VCC_net), .CO(n27841));
    SB_LUT4 communication_counter_31__I_0_add_2189_17_lut (.I0(GND_net), .I1(n3243), 
            .I2(VCC_net), .I3(n27839), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_17 (.CI(n27839), .I0(n3243), 
            .I1(VCC_net), .CO(n27840));
    SB_LUT4 communication_counter_31__I_0_add_2189_16_lut (.I0(GND_net), .I1(n3244), 
            .I2(VCC_net), .I3(n27838), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_16 (.CI(n27838), .I0(n3244), 
            .I1(VCC_net), .CO(n27839));
    SB_LUT4 communication_counter_31__I_0_add_2189_15_lut (.I0(GND_net), .I1(n3245), 
            .I2(VCC_net), .I3(n27837), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_15 (.CI(n27837), .I0(n3245), 
            .I1(VCC_net), .CO(n27838));
    SB_LUT4 communication_counter_31__I_0_add_2189_14_lut (.I0(GND_net), .I1(n3246), 
            .I2(VCC_net), .I3(n27836), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_14 (.CI(n27836), .I0(n3246), 
            .I1(VCC_net), .CO(n27837));
    SB_LUT4 communication_counter_31__I_0_add_2189_13_lut (.I0(GND_net), .I1(n3247), 
            .I2(VCC_net), .I3(n27835), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_13 (.CI(n27835), .I0(n3247), 
            .I1(VCC_net), .CO(n27836));
    SB_LUT4 communication_counter_31__I_0_add_2189_12_lut (.I0(GND_net), .I1(n3248), 
            .I2(VCC_net), .I3(n27834), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_12 (.CI(n27834), .I0(n3248), 
            .I1(VCC_net), .CO(n27835));
    SB_LUT4 communication_counter_31__I_0_add_2189_11_lut (.I0(GND_net), .I1(n3249), 
            .I2(VCC_net), .I3(n27833), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_11 (.CI(n27833), .I0(n3249), 
            .I1(VCC_net), .CO(n27834));
    SB_LUT4 communication_counter_31__I_0_add_2189_10_lut (.I0(GND_net), .I1(n3250), 
            .I2(VCC_net), .I3(n27832), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_10 (.CI(n27832), .I0(n3250), 
            .I1(VCC_net), .CO(n27833));
    SB_LUT4 communication_counter_31__I_0_add_2189_9_lut (.I0(GND_net), .I1(n3251), 
            .I2(VCC_net), .I3(n27831), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_9 (.CI(n27831), .I0(n3251), 
            .I1(VCC_net), .CO(n27832));
    SB_LUT4 communication_counter_31__I_0_add_2189_8_lut (.I0(GND_net), .I1(n3252), 
            .I2(VCC_net), .I3(n27830), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_8 (.CI(n27830), .I0(n3252), 
            .I1(VCC_net), .CO(n27831));
    SB_LUT4 communication_counter_31__I_0_add_2189_7_lut (.I0(GND_net), .I1(n3253), 
            .I2(VCC_net), .I3(n27829), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_7 (.CI(n27829), .I0(n3253), 
            .I1(VCC_net), .CO(n27830));
    SB_LUT4 communication_counter_31__I_0_add_2189_6_lut (.I0(GND_net), .I1(n3254), 
            .I2(GND_net), .I3(n27828), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_6 (.CI(n27828), .I0(n3254), 
            .I1(GND_net), .CO(n27829));
    SB_LUT4 communication_counter_31__I_0_add_2189_5_lut (.I0(GND_net), .I1(n3255), 
            .I2(GND_net), .I3(n27827), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_5 (.CI(n27827), .I0(n3255), 
            .I1(GND_net), .CO(n27828));
    SB_LUT4 i13672_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13950), .I3(GND_net), .O(n18179));   // verilog/coms.v(126[12] 289[6])
    defparam i13672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3930));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1600_3_lut (.I0(n2374), .I1(n6860), .I2(n2381), .I3(GND_net), 
            .O(n2464));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1600_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1654_3_lut (.I0(n2459), .I1(n6876), .I2(n2471), .I3(GND_net), 
            .O(n2546));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4192));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13673_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13950), .I3(GND_net), .O(n18180));   // verilog/coms.v(126[12] 289[6])
    defparam i13673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13674_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13950), .I3(GND_net), .O(n18181));   // verilog/coms.v(126[12] 289[6])
    defparam i13674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13675_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13950), .I3(GND_net), .O(n18182));   // verilog/coms.v(126[12] 289[6])
    defparam i13675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1940_3_lut (.I0(n2851), .I1(n2918), 
            .I2(n2867), .I3(GND_net), .O(n2950));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1939_3_lut (.I0(n2850), .I1(n2917), 
            .I2(n2867), .I3(GND_net), .O(n2949));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34206_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), .I3(GND_net), 
            .O(n2947));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1942_3_lut (.I0(n2853), .I1(n2920), 
            .I2(n2867), .I3(GND_net), .O(n2952));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1934_3_lut (.I0(n2845), .I1(n2912), 
            .I2(n2867), .I3(GND_net), .O(n2944));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1933_3_lut (.I0(n2844), .I1(n2911), 
            .I2(n2867), .I3(GND_net), .O(n2943));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1935_3_lut (.I0(n2846), .I1(n2913), 
            .I2(n2867), .I3(GND_net), .O(n2945));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1136_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n28278), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_2189_4_lut (.I0(GND_net), .I1(n3256), 
            .I2(VCC_net), .I3(n27826), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_4 (.CI(n27826), .I0(n3256), 
            .I1(VCC_net), .CO(n27827));
    SB_LUT4 div_46_i1659_3_lut (.I0(n2464), .I1(n6881), .I2(n2471), .I3(GND_net), 
            .O(n2551));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1936_3_lut (.I0(n2847), .I1(n2914), 
            .I2(n2867), .I3(GND_net), .O(n2946));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1938_3_lut (.I0(n2849), .I1(n2916), 
            .I2(n2867), .I3(GND_net), .O(n2948));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_2189_3_lut (.I0(GND_net), .I1(n3257), 
            .I2(VCC_net), .I3(n27825), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_2189_3 (.CI(n27825), .I0(n3257), 
            .I1(VCC_net), .CO(n27826));
    SB_LUT4 communication_counter_31__I_0_i1941_3_lut (.I0(n2852), .I1(n2919), 
            .I2(n2867), .I3(GND_net), .O(n2951));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1926_3_lut (.I0(n2837), .I1(n2904), 
            .I2(n2867), .I3(GND_net), .O(n2936));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1925_3_lut (.I0(n2836), .I1(n2903), 
            .I2(n2867), .I3(GND_net), .O(n2935));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1924_3_lut (.I0(n2835), .I1(n2902), 
            .I2(n2867), .I3(GND_net), .O(n2934));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1136_add_4_26 (.CI(n28278), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n28279));
    SB_LUT4 communication_counter_1136_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n28277), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1932_3_lut (.I0(n2843), .I1(n2910), 
            .I2(n2867), .I3(GND_net), .O(n2942));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_2189_2_lut (.I0(GND_net), .I1(n3258), 
            .I2(GND_net), .I3(VCC_net), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2189_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n28090), 
            .O(n6914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_25 (.CI(n28277), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n28278));
    SB_CARRY communication_counter_31__I_0_add_2189_2 (.CI(VCC_net), .I0(n3258), 
            .I1(GND_net), .CO(n27825));
    SB_LUT4 communication_counter_31__I_0_i1931_3_lut (.I0(n2842), .I1(n2909), 
            .I2(n2867), .I3(GND_net), .O(n2941));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1117_14 (.CI(n28510), .I0(n1647_adj_4122), 
            .I1(VCC_net), .CO(n28511));
    SB_LUT4 add_3173_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n27824), 
            .O(n6724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_18 (.CI(n28090), .I0(n2623), .I1(n84), .CO(n28091));
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_7 (.CI(n29190), 
            .I0(GND_net), .I1(n28_adj_4594), .CO(n29191));
    SB_LUT4 add_3173_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n27823), 
            .O(n6725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1945_3_lut (.I0(n2856), .I1(n2923), 
            .I2(n2867), .I3(GND_net), .O(n2955));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3173_12 (.CI(n27823), .I0(n1644), .I1(n90), .CO(n27824));
    SB_LUT4 communication_counter_31__I_0_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4123), 
            .I2(VCC_net), .I3(n28509), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n28276), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_4595), .I3(n29189), .O(n29_adj_3957)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_6 (.CI(n29189), 
            .I0(GND_net), .I1(n29_adj_4595), .CO(n29190));
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_4596), .I3(n29188), .O(n30_adj_3956)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_5 (.CI(n29188), 
            .I0(GND_net), .I1(n30_adj_4596), .CO(n29189));
    SB_LUT4 add_3173_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n27822), 
            .O(n6726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n28089), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_4597), .I3(n29187), .O(n31_adj_3955)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_11 (.CI(n27822), .I0(n1645), .I1(n91), .CO(n27823));
    SB_LUT4 communication_counter_31__I_0_i1943_3_lut (.I0(n2854), .I1(n2921), 
            .I2(n2867), .I3(GND_net), .O(n2953));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3183_17 (.CI(n28089), .I0(n2624), .I1(n85), .CO(n28090));
    SB_CARRY communication_counter_1136_add_4_24 (.CI(n28276), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n28277));
    SB_LUT4 add_3173_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n27821), 
            .O(n6727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_13 (.CI(n28509), .I0(n1648_adj_4123), 
            .I1(VCC_net), .CO(n28510));
    SB_LUT4 communication_counter_31__I_0_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4124), 
            .I2(VCC_net), .I3(n28508), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_4 (.CI(n29187), 
            .I0(GND_net), .I1(n31_adj_4597), .CO(n29188));
    SB_LUT4 communication_counter_31__I_0_i1944_3_lut (.I0(n2855), .I1(n2922), 
            .I2(n2867), .I3(GND_net), .O(n2954));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1117_12 (.CI(n28508), .I0(n1649_adj_4124), 
            .I1(VCC_net), .CO(n28509));
    SB_CARRY add_3173_10 (.CI(n27821), .I0(n1646), .I1(n92), .CO(n27822));
    SB_LUT4 communication_counter_31__I_0_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4125), 
            .I2(VCC_net), .I3(n28507), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_mux_3_i7_3_lut (.I0(communication_counter[6]), 
            .I1(n27), .I2(communication_counter[31]), .I3(GND_net), .O(n2958));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1947_3_lut (.I0(n2858), .I1(n2925), 
            .I2(n2867), .I3(GND_net), .O(n2957));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3183_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n28088), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_11 (.CI(n28507), .I0(n1650_adj_4125), 
            .I1(VCC_net), .CO(n28508));
    SB_LUT4 communication_counter_31__I_0_i1946_3_lut (.I0(n2857_adj_4078), 
            .I1(n2924), .I2(n2867), .I3(GND_net), .O(n2956));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1136_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n28275), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1869_3_lut (.I0(n2748_adj_4086), 
            .I1(n2815), .I2(n2768), .I3(GND_net), .O(n2847));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1870_3_lut (.I0(n2749_adj_4085), 
            .I1(n2816), .I2(n2768), .I3(GND_net), .O(n2848));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4126), 
            .I2(VCC_net), .I3(n28506), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3173_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n27820), 
            .O(n6728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i1866_3_lut (.I0(n2745_adj_4089), 
            .I1(n2812), .I2(n2768), .I3(GND_net), .O(n2844));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3173_9 (.CI(n27820), .I0(n1647), .I1(n93), .CO(n27821));
    SB_LUT4 add_3173_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n27819), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_3990), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1865_3_lut (.I0(n2744_adj_4090), 
            .I1(n2811), .I2(n2768), .I3(GND_net), .O(n2843));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3173_8 (.CI(n27819), .I0(n1648), .I1(n94), .CO(n27820));
    SB_LUT4 communication_counter_31__I_0_i1868_3_lut (.I0(n2747_adj_4087), 
            .I1(n2814), .I2(n2768), .I3(GND_net), .O(n2846));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_3_lut_adj_1573 (.I0(bit_ctr[4]), .I1(n39063), .I2(n17536), 
            .I3(GND_net), .O(n32678));   // verilog/neopixel.v(35[12] 117[6])
    defparam i21_3_lut_adj_1573.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1871_3_lut (.I0(n2750_adj_4084), 
            .I1(n2817), .I2(n2768), .I3(GND_net), .O(n2849));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1136_add_4_23 (.CI(n28275), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n28276));
    SB_LUT4 div_46_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4444));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3173_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n27818), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4445));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3173_7 (.CI(n27818), .I0(n1649), .I1(n95), .CO(n27819));
    SB_LUT4 communication_counter_31__I_0_i1875_3_lut (.I0(n2754_adj_4080), 
            .I1(n2821), .I2(n2768), .I3(GND_net), .O(n2853));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3173_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n27817), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_6 (.CI(n27817), .I0(n1650), .I1(n96), .CO(n27818));
    SB_LUT4 div_46_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4446));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3173_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n27816), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1874_3_lut (.I0(n2753_adj_4081), 
            .I1(n2820), .I2(n2768), .I3(GND_net), .O(n2852));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1867_3_lut (.I0(n2746_adj_4088), 
            .I1(n2813), .I2(n2768), .I3(GND_net), .O(n2845));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1873_3_lut (.I0(n2752_adj_4082), 
            .I1(n2819), .I2(n2768), .I3(GND_net), .O(n2851));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4055), .I3(n29186), .O(n32_adj_3954)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1872_3_lut (.I0(n2751_adj_4083), 
            .I1(n2818), .I2(n2768), .I3(GND_net), .O(n2850));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3173_5 (.CI(n27816), .I0(n1651), .I1(n97), .CO(n27817));
    SB_LUT4 communication_counter_31__I_0_i1862_3_lut (.I0(n2741_adj_4093), 
            .I1(n2808), .I2(n2768), .I3(GND_net), .O(n2840));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3173_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n27815), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33347_4_lut (.I0(n35_adj_4446), .I1(n23_adj_4439), .I2(n21_adj_4438), 
            .I3(n19_adj_4436), .O(n39669));
    defparam i33347_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3173_4 (.CI(n27815), .I0(n1652), .I1(n98), .CO(n27816));
    SB_CARRY add_3183_16 (.CI(n28088), .I0(n2625), .I1(n86), .CO(n28089));
    SB_LUT4 add_3173_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n27814), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3173_3 (.CI(n27814), .I0(n1653), .I1(n99), .CO(n27815));
    SB_LUT4 add_3173_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3173_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33890_4_lut (.I0(n17_adj_4434), .I1(n15_adj_4432), .I2(n2464), 
            .I3(n98), .O(n40212));
    defparam i33890_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY add_3173_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n27814));
    SB_LUT4 communication_counter_31__I_0_i1857_3_lut (.I0(n2736_adj_4098), 
            .I1(n2803), .I2(n2768), .I3(GND_net), .O(n2835));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1877_3_lut (.I0(n2756), .I1(n2823), 
            .I2(n2768), .I3(GND_net), .O(n2855));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1876_3_lut (.I0(n2755_adj_4079), 
            .I1(n2822), .I2(n2768), .I3(GND_net), .O(n2854));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3172_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n27813), 
            .O(n6711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1864_3_lut (.I0(n2743_adj_4091), 
            .I1(n2810), .I2(n2768), .I3(GND_net), .O(n2842));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i8_3_lut (.I0(communication_counter[7]), 
            .I1(n26_adj_3959), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2858));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1117_10 (.CI(n28506), .I0(n1651_adj_4126), 
            .I1(VCC_net), .CO(n28507));
    SB_LUT4 add_3172_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n27812), 
            .O(n6712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4127), 
            .I2(VCC_net), .I3(n28505), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_3 (.CI(n29186), 
            .I0(GND_net), .I1(n7_adj_4055), .CO(n29187));
    SB_CARRY communication_counter_31__I_0_add_1117_9 (.CI(n28505), .I0(n1652_adj_4127), 
            .I1(VCC_net), .CO(n28506));
    SB_LUT4 communication_counter_31__I_0_i1879_3_lut (.I0(n2758), .I1(n2825), 
            .I2(n2768), .I3(GND_net), .O(n2857_adj_4078));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3172_11 (.CI(n27812), .I0(n1530), .I1(n91), .CO(n27813));
    SB_LUT4 communication_counter_31__I_0_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4128), 
            .I2(VCC_net), .I3(n28504), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_8 (.CI(n28504), .I0(n1653_adj_4128), 
            .I1(VCC_net), .CO(n28505));
    SB_LUT4 communication_counter_31__I_0_i1878_3_lut (.I0(n2757), .I1(n2824), 
            .I2(n2768), .I3(GND_net), .O(n2856));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1807_3_lut (.I0(n2654), .I1(n2721), 
            .I2(n2669), .I3(GND_net), .O(n2753_adj_4081));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1117_7_lut (.I0(GND_net), .I1(n1654), 
            .I2(GND_net), .I3(n28503), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n28274), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13687_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13950), .I3(GND_net), .O(n18194));   // verilog/coms.v(126[12] 289[6])
    defparam i13687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3172_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n27811), 
            .O(n6713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_7 (.CI(n28503), .I0(n1654), 
            .I1(GND_net), .CO(n28504));
    SB_CARRY communication_counter_1136_add_4_22 (.CI(n28274), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n28275));
    SB_LUT4 communication_counter_1136_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n28273), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1792_3_lut (.I0(n2639), .I1(n2706_adj_4116), 
            .I2(n2669), .I3(GND_net), .O(n2738_adj_4096));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1791_3_lut (.I0(n2638_adj_4136), 
            .I1(n2705_adj_4117), .I2(n2669), .I3(GND_net), .O(n2737_adj_4097));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1790_3_lut (.I0(n2637_adj_4137), 
            .I1(n2704_adj_4118), .I2(n2669), .I3(GND_net), .O(n2736_adj_4098));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1809_3_lut (.I0(n2656), .I1(n2723_adj_4101), 
            .I2(n2669), .I3(GND_net), .O(n2755_adj_4079));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1808_3_lut (.I0(n2655), .I1(n2722), 
            .I2(n2669), .I3(GND_net), .O(n2754_adj_4080));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i9_3_lut (.I0(communication_counter[8]), 
            .I1(n25_adj_3960), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2758));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3172_10 (.CI(n27811), .I0(n1531), .I1(n92), .CO(n27812));
    SB_CARRY communication_counter_1136_add_4_21 (.CI(n28273), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n28274));
    SB_LUT4 communication_counter_31__I_0_i1811_3_lut (.I0(n2658), .I1(n2725), 
            .I2(n2669), .I3(GND_net), .O(n2757));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1117_6_lut (.I0(GND_net), .I1(n1655), 
            .I2(GND_net), .I3(n28502), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1810_3_lut (.I0(n2657), .I1(n2724_adj_4100), 
            .I2(n2669), .I3(GND_net), .O(n2756));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_4598), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_4598), .CO(n29186));
    SB_LUT4 communication_counter_1136_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n28272), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_4_lut (.I0(duty[2]), .I1(n41708), .I2(n23), .I3(n27569), 
            .O(pwm_setpoint_22__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_3_lut_adj_1574 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n34698));
    defparam i1_3_lut_adj_1574.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut (.I0(n2750_adj_4084), .I1(n2745_adj_4089), .I2(n2746_adj_4088), 
            .I3(n2749_adj_4085), .O(n34));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(n2743_adj_4091), .I1(n2754_adj_4080), .I2(n34698), 
            .I3(n2755_adj_4079), .O(n25_adj_3933));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut (.I0(n2739_adj_4095), .I1(n2741_adj_4093), .I2(n2740_adj_4094), 
            .I3(n2742_adj_4092), .O(n32));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2736_adj_4098), .I1(n2737_adj_4097), .I2(n2735_adj_4099), 
            .I3(n2738_adj_4096), .O(n31));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1575 (.I0(n2753_adj_4081), .I1(n2752_adj_4082), 
            .I2(n2751_adj_4083), .I3(n2748_adj_4086), .O(n35));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n25_adj_3933), .I1(n34), .I2(n2747_adj_4087), 
            .I3(n2744_adj_4090), .O(n37));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13688_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13950), .I3(GND_net), .O(n18195));   // verilog/coms.v(126[12] 289[6])
    defparam i13688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3172_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n27810), 
            .O(n6714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_20 (.CI(n28272), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n28273));
    SB_CARRY add_3172_9 (.CI(n27810), .I0(n1532), .I1(n93), .CO(n27811));
    SB_LUT4 add_3172_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n27809), 
            .O(n6715)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n28271), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_6 (.CI(n28502), .I0(n1655), 
            .I1(GND_net), .CO(n28503));
    SB_LUT4 i13689_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13950), .I3(GND_net), .O(n18196));   // verilog/coms.v(126[12] 289[6])
    defparam i13689_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3172_8 (.CI(n27809), .I0(n1533), .I1(n94), .CO(n27810));
    SB_LUT4 add_3183_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n28087), 
            .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_19 (.CI(n28271), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n28272));
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31), .I3(n32), .O(n2768));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_add_1117_5_lut (.I0(GND_net), .I1(n1656), 
            .I2(VCC_net), .I3(n28501), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3172_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n27808), 
            .O(n6716)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1861_3_lut (.I0(n2740_adj_4094), 
            .I1(n2807), .I2(n2768), .I3(GND_net), .O(n2839));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1117_5 (.CI(n28501), .I0(n1656), 
            .I1(VCC_net), .CO(n28502));
    SB_LUT4 communication_counter_1136_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n28270), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1859_3_lut (.I0(n2738_adj_4096), 
            .I1(n2805), .I2(n2768), .I3(GND_net), .O(n2837));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3172_7 (.CI(n27808), .I0(n1534), .I1(n95), .CO(n27809));
    SB_LUT4 communication_counter_31__I_0_i1860_3_lut (.I0(n2739_adj_4095), 
            .I1(n2806), .I2(n2768), .I3(GND_net), .O(n2838));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1136_add_4_18 (.CI(n28270), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n28271));
    SB_LUT4 communication_counter_31__I_0_i1858_3_lut (.I0(n2737_adj_4097), 
            .I1(n2804), .I2(n2768), .I3(GND_net), .O(n2836));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1576 (.I0(n2856), .I1(n2857_adj_4078), .I2(n2858), 
            .I3(GND_net), .O(n34769));
    defparam i1_3_lut_adj_1576.LUT_INIT = 16'hfefe;
    SB_LUT4 i13690_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13950), .I3(GND_net), .O(n18197));   // verilog/coms.v(126[12] 289[6])
    defparam i13690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1577 (.I0(n2842), .I1(n2854), .I2(n34769), .I3(n2855), 
            .O(n26_adj_4049));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_4_lut_adj_1577.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut_adj_1578 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33_adj_4048));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1579 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4050));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i1_2_lut_adj_1579.LUT_INIT = 16'heeee;
    SB_LUT4 i13691_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13950), 
            .I3(GND_net), .O(n18198));   // verilog/coms.v(126[12] 289[6])
    defparam i13691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_4_lut_adj_1580 (.I0(n33_adj_4048), .I1(n2840), .I2(n26_adj_4049), 
            .I3(n2841), .O(n38_adj_4044));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1581 (.I0(n2850), .I1(n2851), .I2(n2845), .I3(n2852), 
            .O(n36_adj_4046));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2853), .I1(n2849), .I2(n2846), .I3(n22_adj_4050), 
            .O(n37_adj_4045));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3172_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n27807), 
            .O(n6717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_6 (.CI(n27807), .I0(n1535), .I1(n96), .CO(n27808));
    SB_LUT4 communication_counter_1136_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n28269), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1117_4_lut (.I0(GND_net), .I1(n1657), 
            .I2(VCC_net), .I3(n28500), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_17 (.CI(n28269), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n28270));
    SB_CARRY add_3183_15 (.CI(n28087), .I0(n2626), .I1(n87), .CO(n28088));
    SB_CARRY communication_counter_31__I_0_add_1117_4 (.CI(n28500), .I0(n1657), 
            .I1(VCC_net), .CO(n28501));
    SB_LUT4 add_3183_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n28086), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1117_3_lut (.I0(GND_net), .I1(n1658), 
            .I2(GND_net), .I3(n28499), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_3 (.CI(n28499), .I0(n1658), 
            .I1(GND_net), .CO(n28500));
    SB_LUT4 add_3172_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n27806), 
            .O(n6718)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_14 (.CI(n28086), .I0(n2627), .I1(n88), .CO(n28087));
    SB_LUT4 i14_4_lut_adj_1582 (.I0(n2843), .I1(n2844), .I2(n2848), .I3(n2847), 
            .O(n35_adj_4047));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_1136_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n28268), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4346), 
            .I1(VCC_net), .CO(n28499));
    SB_CARRY add_3172_5 (.CI(n27806), .I0(n1536), .I1(n97), .CO(n27807));
    SB_LUT4 i20_4_lut (.I0(n35_adj_4047), .I1(n37_adj_4045), .I2(n36_adj_4046), 
            .I3(n38_adj_4044), .O(n2867));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3172_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n27805), 
            .O(n6719)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1863_3_lut (.I0(n2742_adj_4092), 
            .I1(n2809), .I2(n2768), .I3(GND_net), .O(n2841));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1930_3_lut (.I0(n2841), .I1(n2908), 
            .I2(n2867), .I3(GND_net), .O(n2940));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1184_16_lut (.I0(n1745), .I1(n1745), 
            .I2(n1778_adj_4345), .I3(n28498), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 communication_counter_31__I_0_add_1184_15_lut (.I0(n1746), .I1(n1746), 
            .I2(n1778_adj_4345), .I3(n28497), .O(n1845)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_1545_i26_3_lut (.I0(n18_adj_4411), .I1(n91), 
            .I2(n29_adj_4420), .I3(GND_net), .O(n26_adj_4418));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3172_4 (.CI(n27805), .I0(n1537), .I1(n98), .CO(n27806));
    SB_DFF communication_counter_1136__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_LUT4 i34506_4_lut (.I0(n26_adj_4418), .I1(n16_adj_4409), .I2(n29_adj_4420), 
            .I3(n39736), .O(n40828));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34506_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3172_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n27804), 
            .O(n6720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34507_3_lut (.I0(n40828), .I1(n90), .I2(n31_adj_4421), .I3(GND_net), 
            .O(n40829));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34507_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_i1928_3_lut (.I0(n2839), .I1(n2906), 
            .I2(n2867), .I3(GND_net), .O(n2938));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34397_3_lut (.I0(n40829), .I1(n89), .I2(n33_adj_4422), .I3(GND_net), 
            .O(n40719));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34397_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_i1929_3_lut (.I0(n2840), .I1(n2907), 
            .I2(n2867), .I3(GND_net), .O(n2939));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1927_3_lut (.I0(n2838), .I1(n2905), 
            .I2(n2867), .I3(GND_net), .O(n2937));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34326_4_lut (.I0(n43_adj_4428), .I1(n41_adj_4427), .I2(n39_adj_4425), 
            .I3(n39726), .O(n40648));
    defparam i34326_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34536_4_lut (.I0(n39969), .I1(n40594), .I2(n45_adj_4429), 
            .I3(n39713), .O(n40858));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34536_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33645_3_lut (.I0(n40719), .I1(n88), .I2(n35_adj_4423), .I3(GND_net), 
            .O(n39967));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33645_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_3_lut_adj_1583 (.I0(n2956), .I1(n2957), .I2(n2958), .I3(GND_net), 
            .O(n34715));
    defparam i1_3_lut_adj_1583.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(n2954), .I1(n2953), .I2(n34715), .I3(n2955), 
            .O(n28_adj_4554));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i6_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i34538_4_lut (.I0(n39967), .I1(n40858), .I2(n45_adj_4429), 
            .I3(n40648), .O(n40860));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34538_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY communication_counter_31__I_0_add_1184_15 (.CI(n28497), .I0(n1746), 
            .I1(n1778_adj_4345), .CO(n28498));
    SB_LUT4 i1_4_lut_adj_1584 (.I0(n40860), .I1(n16498), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'hceef;
    SB_LUT4 communication_counter_31__I_0_i1804_3_lut (.I0(n2651), .I1(n2718_adj_4104), 
            .I2(n2669), .I3(GND_net), .O(n2750_adj_4084));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35_adj_4551));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1585 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_4552));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1586 (.I0(n35_adj_4551), .I1(n2941), .I2(n28_adj_4554), 
            .I3(n2942), .O(n40_adj_4547));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i18_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1658_3_lut (.I0(n2463), .I1(n6880), .I2(n2471), .I3(GND_net), 
            .O(n2550));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_add_1184_14_lut (.I0(n1747), .I1(n1747), 
            .I2(n1778_adj_4345), .I3(n28496), .O(n1846)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY communication_counter_1136_add_4_16 (.CI(n28268), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n28269));
    SB_LUT4 i13692_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13950), 
            .I3(GND_net), .O(n18199));   // verilog/coms.v(126[12] 289[6])
    defparam i13692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3183_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n28085), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4187));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_1184_14 (.CI(n28496), .I0(n1747), 
            .I1(n1778_adj_4345), .CO(n28497));
    SB_LUT4 communication_counter_1136_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n28267), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4186));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3183_13 (.CI(n28085), .I0(n2628), .I1(n89), .CO(n28086));
    SB_LUT4 communication_counter_31__I_0_i1803_3_lut (.I0(n2650), .I1(n2717_adj_4105), 
            .I2(n2669), .I3(GND_net), .O(n2749_adj_4085));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4249));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4253));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4258));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3183_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n28084), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1184_13_lut (.I0(n1748), .I1(n1748), 
            .I2(n1778_adj_4345), .I3(n28495), .O(n1847)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4263));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4264));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1525_3_lut (.I0(n2267), .I1(n6826), .I2(n2288), .I3(GND_net), 
            .O(n2360));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4262));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4265));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3172_3 (.CI(n27804), .I0(n1538), .I1(n99), .CO(n27805));
    SB_CARRY communication_counter_31__I_0_add_1184_13 (.CI(n28495), .I0(n1748), 
            .I1(n1778_adj_4345), .CO(n28496));
    SB_CARRY add_3183_12 (.CI(n28084), .I0(n2629), .I1(n90), .CO(n28085));
    SB_LUT4 add_3183_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n28083), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4270));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1184_12_lut (.I0(n1749), .I1(n1749), 
            .I2(n1778_adj_4345), .I3(n28494), .O(n1848)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4271));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3172_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3172_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3172_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n27804));
    SB_LUT4 add_3171_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n27803), 
            .O(n6699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_15 (.CI(n28267), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n28268));
    SB_LUT4 communication_counter_1136_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n28266), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4269));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4272));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4278));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4276));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1136_add_4_14 (.CI(n28266), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n28267));
    SB_LUT4 add_3171_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n27802), 
            .O(n6700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1184_12 (.CI(n28494), .I0(n1749), 
            .I1(n1778_adj_4345), .CO(n28495));
    SB_LUT4 communication_counter_31__I_0_add_1184_11_lut (.I0(n1750), .I1(n1750), 
            .I2(n1778_adj_4345), .I3(n28493), .O(n1849)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 communication_counter_1136_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n28265), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_10 (.CI(n27802), .I0(n1413), .I1(n92), .CO(n27803));
    SB_LUT4 div_46_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4279));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4280));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1184_11 (.CI(n28493), .I0(n1750), 
            .I1(n1778_adj_4345), .CO(n28494));
    SB_LUT4 div_46_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4283));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1136_add_4_13 (.CI(n28265), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n28266));
    SB_LUT4 div_46_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4281));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1184_10_lut (.I0(n1751), .I1(n1751), 
            .I2(n1778_adj_4345), .I3(n28492), .O(n1850)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4284));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_1136_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n28264), .O(n155_adj_4129)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_11 (.CI(n28083), .I0(n2630), .I1(n91), .CO(n28084));
    SB_LUT4 add_3171_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n27801), 
            .O(n6701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_9 (.CI(n27801), .I0(n1414), .I1(n93), .CO(n27802));
    SB_CARRY communication_counter_31__I_0_add_1184_10 (.CI(n28492), .I0(n1751), 
            .I1(n1778_adj_4345), .CO(n28493));
    SB_LUT4 communication_counter_31__I_0_add_1184_9_lut (.I0(n1752), .I1(n1752), 
            .I2(n1778_adj_4345), .I3(n28491), .O(n1851)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_3183_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n28082), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3171_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n27800), 
            .O(n6702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_8 (.CI(n27800), .I0(n1415), .I1(n94), .CO(n27801));
    SB_CARRY communication_counter_31__I_0_add_1184_9 (.CI(n28491), .I0(n1752), 
            .I1(n1778_adj_4345), .CO(n28492));
    SB_LUT4 communication_counter_31__I_0_add_1184_8_lut (.I0(n1753), .I1(n1753), 
            .I2(n1778_adj_4345), .I3(n28490), .O(n1852)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4290));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1136_add_4_12 (.CI(n28264), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n28265));
    SB_LUT4 div_46_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4288));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1184_8 (.CI(n28490), .I0(n1753), 
            .I1(n1778_adj_4345), .CO(n28491));
    SB_LUT4 communication_counter_1136_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n28263), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_11 (.CI(n28263), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n28264));
    SB_LUT4 add_3171_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n27799), 
            .O(n6703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4291));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3183_10 (.CI(n28082), .I0(n2631), .I1(n92), .CO(n28083));
    SB_LUT4 add_3183_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n28081), 
            .O(n6923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_9 (.CI(n28081), .I0(n2632), .I1(n93), .CO(n28082));
    SB_LUT4 communication_counter_31__I_0_add_1184_7_lut (.I0(n1754_adj_4367), 
            .I1(n1754_adj_4367), .I2(n41718), .I3(n28489), .O(n1853)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_3171_7 (.CI(n27799), .I0(n1416), .I1(n95), .CO(n27800));
    SB_LUT4 add_3171_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n27798), 
            .O(n6704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n28262), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_6 (.CI(n27798), .I0(n1417), .I1(n96), .CO(n27799));
    SB_LUT4 add_3171_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n27797), 
            .O(n6705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_5 (.CI(n27797), .I0(n1418), .I1(n97), .CO(n27798));
    SB_LUT4 div_46_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4292));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1184_7 (.CI(n28489), .I0(n1754_adj_4367), 
            .I1(n41718), .CO(n28490));
    SB_LUT4 add_3171_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n27796), 
            .O(n6706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4295));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4293));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4296));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_DFF communication_counter_1136__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155_adj_4129));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF communication_counter_1136__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(48[28:51])
    SB_DFF blue_1137__i1 (.Q(blue[1]), .C(LED_c), .D(n44_adj_4153));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_DFF blue_1137__i2 (.Q(blue[2]), .C(LED_c), .D(n43_adj_4152));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_LUT4 communication_counter_31__I_0_add_1184_6_lut (.I0(n1755_adj_4366), 
            .I1(n1755_adj_4366), .I2(n41718), .I3(n28488), .O(n1854)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY communication_counter_31__I_0_add_1184_6 (.CI(n28488), .I0(n1755_adj_4366), 
            .I1(n41718), .CO(n28489));
    SB_CARRY communication_counter_1136_add_4_10 (.CI(n28262), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n28263));
    SB_LUT4 communication_counter_1136_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n28261), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n28080), 
            .O(n6924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_8 (.CI(n28080), .I0(n2633), .I1(n94), .CO(n28081));
    SB_CARRY add_3171_4 (.CI(n27796), .I0(n1419), .I1(n98), .CO(n27797));
    SB_LUT4 add_3171_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n27795), 
            .O(n6707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3171_3 (.CI(n27795), .I0(n1420), .I1(n99), .CO(n27796));
    SB_LUT4 div_46_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4302));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3171_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6708)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3171_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_9 (.CI(n28261), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n28262));
    SB_LUT4 div_46_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4300));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4303));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1184_5_lut (.I0(n1756_adj_4348), 
            .I1(n1756_adj_4348), .I2(n1778_adj_4345), .I3(n28487), .O(n1855)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 div_46_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4304));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3171_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n27795));
    SB_LUT4 communication_counter_1136_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n28260), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n28079), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_2298_9_lut (.I0(n39039), .I1(GND_net), 
            .I2(n3452), .I3(n27794), .O(n39038)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3183_7 (.CI(n28079), .I0(n2634), .I1(n95), .CO(n28080));
    SB_CARRY communication_counter_31__I_0_add_1184_5 (.CI(n28487), .I0(n1756_adj_4348), 
            .I1(n1778_adj_4345), .CO(n28488));
    SB_CARRY communication_counter_1136_add_4_8 (.CI(n28260), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n28261));
    SB_LUT4 communication_counter_31__I_0_add_1184_4_lut (.I0(n1757_adj_4347), 
            .I1(n1757_adj_4347), .I2(n1778_adj_4345), .I3(n28486), .O(n1856)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFF blue_1137__i3 (.Q(blue[3]), .C(LED_c), .D(n42_adj_4151));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_DFF blue_1137__i4 (.Q(blue[4]), .C(LED_c), .D(n41_adj_4150));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_DFF blue_1137__i5 (.Q(blue[5]), .C(LED_c), .D(n40_adj_4149));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_DFF blue_1137__i6 (.Q(blue[6]), .C(LED_c), .D(n39_adj_4148));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_DFF blue_1137__i7 (.Q(blue[7]), .C(LED_c), .D(n38_adj_4147));   // verilog/TinyFPGA_B.v(53[13:19])
    SB_LUT4 communication_counter_31__I_0_add_2298_8_lut (.I0(n36485), .I1(GND_net), 
            .I2(n3453), .I3(n27793), .O(n39039)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY communication_counter_31__I_0_add_2298_8 (.CI(n27793), .I0(GND_net), 
            .I1(n3453), .CO(n27794));
    SB_LUT4 communication_counter_31__I_0_add_2298_7_lut (.I0(n36483), .I1(GND_net), 
            .I2(n3454), .I3(n27792), .O(n36485)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY communication_counter_31__I_0_add_2298_7 (.CI(n27792), .I0(GND_net), 
            .I1(n3454), .CO(n27793));
    SB_LUT4 communication_counter_31__I_0_add_2298_6_lut (.I0(n36481), .I1(GND_net), 
            .I2(n3455), .I3(n27791), .O(n36483)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY communication_counter_31__I_0_add_2298_6 (.CI(n27791), .I0(GND_net), 
            .I1(n3455), .CO(n27792));
    SB_LUT4 communication_counter_1136_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n28259), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1184_4 (.CI(n28486), .I0(n1757_adj_4347), 
            .I1(n1778_adj_4345), .CO(n28487));
    SB_CARRY communication_counter_1136_add_4_7 (.CI(n28259), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n28260));
    SB_LUT4 add_3183_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n28078), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_6 (.CI(n28078), .I0(n2635), .I1(n96), .CO(n28079));
    SB_LUT4 communication_counter_31__I_0_add_2298_5_lut (.I0(n36479), .I1(GND_net), 
            .I2(n3456), .I3(n27790), .O(n36481)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_5_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_46_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4307));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_2298_5 (.CI(n27790), .I0(GND_net), 
            .I1(n3456), .CO(n27791));
    SB_LUT4 communication_counter_31__I_0_add_1184_3_lut (.I0(n1758_adj_4346), 
            .I1(n1758_adj_4346), .I2(n41718), .I3(n28485), .O(n1857)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1184_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 communication_counter_31__I_0_add_2298_4_lut (.I0(n36477), .I1(GND_net), 
            .I2(n3457), .I3(n27789), .O(n36479)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_4_lut.LUT_INIT = 16'hebbe;
    SB_CARRY communication_counter_31__I_0_add_2298_4 (.CI(n27789), .I0(GND_net), 
            .I1(n3457), .CO(n27790));
    SB_LUT4 communication_counter_31__I_0_add_2298_3_lut (.I0(n3477), .I1(GND_net), 
            .I2(n3458), .I3(n27788), .O(n36477)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_46_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4305));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1184_3 (.CI(n28485), .I0(n1758_adj_4346), 
            .I1(n41718), .CO(n28486));
    SB_CARRY communication_counter_31__I_0_add_2298_3 (.CI(n27788), .I0(GND_net), 
            .I1(n3458), .CO(n27789));
    SB_CARRY communication_counter_31__I_0_add_1184_2 (.CI(VCC_net), .I0(n1858), 
            .I1(VCC_net), .CO(n28485));
    SB_LUT4 communication_counter_31__I_0_add_1251_17_lut (.I0(n1877), .I1(n1844), 
            .I2(VCC_net), .I3(n28484), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4308));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_2298_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3459), .I3(VCC_net), .O(n3477)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_2298_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1251_16_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n28483), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n28258), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n28077), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_16 (.CI(n28483), .I0(n1845), 
            .I1(VCC_net), .CO(n28484));
    SB_LUT4 div_46_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4316));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_2298_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n3459), .CO(n27788));
    SB_LUT4 div_46_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4318));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4314));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1251_15_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n28482), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_6 (.CI(n28258), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n28259));
    SB_LUT4 div_46_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4321));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1251_15 (.CI(n28482), .I0(n1846), 
            .I1(VCC_net), .CO(n28483));
    SB_LUT4 add_3170_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n27787), 
            .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1136_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n28257), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_5 (.CI(n28077), .I0(n2636), .I1(n97), .CO(n28078));
    SB_CARRY communication_counter_1136_add_4_5 (.CI(n28257), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n28258));
    SB_LUT4 communication_counter_31__I_0_add_1251_14_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n28481), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3183_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n28076), 
            .O(n6928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n27786), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_9 (.CI(n27786), .I0(n1293), .I1(n93), .CO(n27787));
    SB_LUT4 add_3170_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n27785), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_4 (.CI(n27569), .I0(n41708), .I1(n23), .CO(n27570));
    SB_CARRY communication_counter_31__I_0_add_1251_14 (.CI(n28481), .I0(n1847), 
            .I1(VCC_net), .CO(n28482));
    SB_LUT4 div_46_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4312));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4322));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4323));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1251_13_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n28480), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4324));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_1136_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n28256), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_4 (.CI(n28076), .I0(n2637), .I1(n98), .CO(n28077));
    SB_CARRY add_3170_8 (.CI(n27785), .I0(n1294), .I1(n94), .CO(n27786));
    SB_LUT4 add_3183_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n28075), 
            .O(n6929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4319));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4326));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3170_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n27784), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_13 (.CI(n28480), .I0(n1848), 
            .I1(VCC_net), .CO(n28481));
    SB_CARRY communication_counter_1136_add_4_4 (.CI(n28256), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n28257));
    SB_LUT4 communication_counter_1136_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n28255), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4334));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1251_12_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n28479), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3183_3 (.CI(n28075), .I0(n2638), .I1(n99), .CO(n28076));
    SB_CARRY communication_counter_31__I_0_add_1251_12 (.CI(n28479), .I0(n1849), 
            .I1(VCC_net), .CO(n28480));
    SB_LUT4 communication_counter_31__I_0_add_1251_11_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n28478), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_7 (.CI(n27784), .I0(n1295), .I1(n95), .CO(n27785));
    SB_LUT4 add_3183_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3183_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1136_add_4_3 (.CI(n28255), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n28256));
    SB_LUT4 div_46_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4336));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4332));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4339));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3183_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n28075));
    SB_LUT4 add_3182_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n28074), 
            .O(n6886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n27783), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_11 (.CI(n28478), .I0(n1850), 
            .I1(VCC_net), .CO(n28479));
    SB_LUT4 communication_counter_1136_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1136_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3182_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n28073), 
            .O(n6887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1251_10_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n28477), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4330));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4340));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3170_6 (.CI(n27783), .I0(n1296), .I1(n96), .CO(n27784));
    SB_LUT4 div_46_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4341));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_1136_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n28255));
    SB_CARRY communication_counter_31__I_0_add_1251_10 (.CI(n28477), .I0(n1851), 
            .I1(VCC_net), .CO(n28478));
    SB_LUT4 communication_counter_31__I_0_add_1251_9_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n28476), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_9 (.CI(n28476), .I0(n1852), 
            .I1(VCC_net), .CO(n28477));
    SB_LUT4 communication_counter_31__I_0_add_1251_8_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n28475), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_8 (.CI(n28475), .I0(n1853), 
            .I1(VCC_net), .CO(n28476));
    SB_LUT4 communication_counter_31__I_0_add_1653_23_lut (.I0(n2471_adj_4224), 
            .I1(n2438), .I2(VCC_net), .I3(n28254), .O(n2537_adj_4175)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3182_21 (.CI(n28073), .I0(n2535), .I1(n81), .CO(n28074));
    SB_LUT4 add_3170_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n27782), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4342));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1251_7_lut (.I0(GND_net), .I1(n1854), 
            .I2(GND_net), .I3(n28474), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1251_7 (.CI(n28474), .I0(n1854), 
            .I1(GND_net), .CO(n28475));
    SB_CARRY add_3170_5 (.CI(n27782), .I0(n1297), .I1(n97), .CO(n27783));
    SB_LUT4 communication_counter_31__I_0_add_1653_22_lut (.I0(GND_net), .I1(n2439), 
            .I2(VCC_net), .I3(n28253), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_555_3_lut (.I0(duty[1]), .I1(n41708), .I2(n24), .I3(n27568), 
            .O(pwm_setpoint_22__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY communication_counter_31__I_0_add_1653_22 (.CI(n28253), .I0(n2439), 
            .I1(VCC_net), .CO(n28254));
    SB_LUT4 communication_counter_31__I_0_add_1653_21_lut (.I0(GND_net), .I1(n2440), 
            .I2(VCC_net), .I3(n28252), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n27781), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1251_6_lut (.I0(GND_net), .I1(n1855), 
            .I2(GND_net), .I3(n28473), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_21 (.CI(n28252), .I0(n2440), 
            .I1(VCC_net), .CO(n28253));
    SB_LUT4 div_46_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4337));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3182_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n28072), 
            .O(n6888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_4 (.CI(n27781), .I0(n1298), .I1(n98), .CO(n27782));
    SB_LUT4 div_46_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4344));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1251_6 (.CI(n28473), .I0(n1855), 
            .I1(GND_net), .CO(n28474));
    SB_LUT4 communication_counter_31__I_0_add_1653_20_lut (.I0(GND_net), .I1(n2441), 
            .I2(VCC_net), .I3(n28251), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_20 (.CI(n28072), .I0(n2536), .I1(n82), .CO(n28073));
    SB_LUT4 add_3182_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n28071), 
            .O(n6889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1251_5_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n28472), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4356));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1251_5 (.CI(n28472), .I0(n1856), 
            .I1(VCC_net), .CO(n28473));
    SB_CARRY communication_counter_31__I_0_add_1653_20 (.CI(n28251), .I0(n2441), 
            .I1(VCC_net), .CO(n28252));
    SB_CARRY add_3182_19 (.CI(n28071), .I0(n2537), .I1(n83), .CO(n28072));
    SB_LUT4 div_46_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4358));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34117_4_lut (.I0(n23_adj_4439), .I1(n21_adj_4438), .I2(n19_adj_4436), 
            .I3(n40212), .O(n40439));
    defparam i34117_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 communication_counter_31__I_0_add_1251_4_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n28471), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_19_lut (.I0(GND_net), .I1(n2442), 
            .I2(VCC_net), .I3(n28250), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3182_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n28070), 
            .O(n6890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_19 (.CI(n28250), .I0(n2442), 
            .I1(VCC_net), .CO(n28251));
    SB_LUT4 div_46_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4354));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4361));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3170_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n27780), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_3 (.CI(n27780), .I0(n1299), .I1(n99), .CO(n27781));
    SB_CARRY communication_counter_31__I_0_add_1251_4 (.CI(n28471), .I0(n1857), 
            .I1(VCC_net), .CO(n28472));
    SB_LUT4 div_46_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4352));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1653_18_lut (.I0(GND_net), .I1(n2443), 
            .I2(VCC_net), .I3(n28249), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1251_3_lut (.I0(GND_net), .I1(n1858), 
            .I2(GND_net), .I3(n28470), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4362));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4363));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1251_3 (.CI(n28470), .I0(n1858), 
            .I1(GND_net), .CO(n28471));
    SB_CARRY communication_counter_31__I_0_add_1251_2 (.CI(VCC_net), .I0(n1958), 
            .I1(VCC_net), .CO(n28470));
    SB_LUT4 communication_counter_31__I_0_add_1318_18_lut (.I0(n1976_adj_4266), 
            .I1(n1943), .I2(VCC_net), .I3(n28469), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY communication_counter_31__I_0_add_1653_18 (.CI(n28249), .I0(n2443), 
            .I1(VCC_net), .CO(n28250));
    SB_LUT4 add_3170_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_17_lut (.I0(GND_net), .I1(n2444), 
            .I2(VCC_net), .I3(n28248), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_17_lut (.I0(GND_net), .I1(n1944), 
            .I2(VCC_net), .I3(n28468), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_17 (.CI(n28468), .I0(n1944), 
            .I1(VCC_net), .CO(n28469));
    SB_CARRY communication_counter_31__I_0_add_1653_17 (.CI(n28248), .I0(n2444), 
            .I1(VCC_net), .CO(n28249));
    SB_LUT4 div_46_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4364));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3182_18 (.CI(n28070), .I0(n2538), .I1(n84), .CO(n28071));
    SB_CARRY add_3170_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n27780));
    SB_LUT4 communication_counter_31__I_0_add_1653_16_lut (.I0(GND_net), .I1(n2445), 
            .I2(VCC_net), .I3(n28247), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_3 (.CI(n27568), .I0(n41708), .I1(n24), .CO(n27569));
    SB_LUT4 div_46_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4359));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1653_16 (.CI(n28247), .I0(n2445), 
            .I1(VCC_net), .CO(n28248));
    SB_LUT4 add_3182_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n28069), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_16_lut (.I0(GND_net), .I1(n1945), 
            .I2(VCC_net), .I3(n28467), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3182_17 (.CI(n28069), .I0(n2539), .I1(n85), .CO(n28070));
    SB_LUT4 div_46_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4365));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_16 (.CI(n28467), .I0(n1945), 
            .I1(VCC_net), .CO(n28468));
    SB_LUT4 communication_counter_31__I_0_add_1653_15_lut (.I0(GND_net), .I1(n2446), 
            .I2(VCC_net), .I3(n28246), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3169_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n27779), 
            .O(n6678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3169_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n27778), 
            .O(n6679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY communication_counter_31__I_0_add_1653_15 (.CI(n28246), .I0(n2446), 
            .I1(VCC_net), .CO(n28247));
    SB_LUT4 communication_counter_31__I_0_add_1653_14_lut (.I0(GND_net), .I1(n2447_adj_4236), 
            .I2(VCC_net), .I3(n28245), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4375));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_555_2_lut (.I0(duty[0]), .I1(n41708), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_555_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3169_8 (.CI(n27778), .I0(n1170), .I1(n94), .CO(n27779));
    SB_LUT4 div_46_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4377));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_15_lut (.I0(GND_net), .I1(n1946), 
            .I2(VCC_net), .I3(n28466), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_555_2 (.CI(VCC_net), .I0(n41708), .I1(n25), .CO(n27568));
    SB_CARRY communication_counter_31__I_0_add_1653_14 (.CI(n28245), .I0(n2447_adj_4236), 
            .I1(VCC_net), .CO(n28246));
    SB_LUT4 add_3182_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n28068), 
            .O(n6892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4378));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4373));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_15 (.CI(n28466), .I0(n1946), 
            .I1(VCC_net), .CO(n28467));
    SB_LUT4 div_46_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4380));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3169_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n27777), 
            .O(n6680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_14_lut (.I0(GND_net), .I1(n1947), 
            .I2(VCC_net), .I3(n28465), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_14 (.CI(n28465), .I0(n1947), 
            .I1(VCC_net), .CO(n28466));
    SB_LUT4 communication_counter_31__I_0_add_1653_13_lut (.I0(GND_net), .I1(n2448_adj_4235), 
            .I2(VCC_net), .I3(n28244), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4371));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3182_16 (.CI(n28068), .I0(n2540), .I1(n86), .CO(n28069));
    SB_LUT4 div_46_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4381));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4382));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1653_13 (.CI(n28244), .I0(n2448_adj_4235), 
            .I1(VCC_net), .CO(n28245));
    SB_LUT4 add_3182_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n28067), 
            .O(n6893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3182_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4383));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_13_lut (.I0(GND_net), .I1(n1948), 
            .I2(VCC_net), .I3(n28464), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4385));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4387));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_13 (.CI(n28464), .I0(n1948), 
            .I1(VCC_net), .CO(n28465));
    SB_LUT4 communication_counter_31__I_0_add_1653_12_lut (.I0(GND_net), .I1(n2449_adj_4234), 
            .I2(VCC_net), .I3(n28243), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_7 (.CI(n27777), .I0(n1171), .I1(n95), .CO(n27778));
    SB_LUT4 add_3169_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n27776), 
            .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4384));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3182_10 (.CI(n28062), .I0(n2546), .I1(n92), .CO(n28063));
    SB_CARRY add_3169_6 (.CI(n27776), .I0(n1172), .I1(n96), .CO(n27777));
    SB_CARRY communication_counter_31__I_0_add_1653_12 (.CI(n28243), .I0(n2449_adj_4234), 
            .I1(VCC_net), .CO(n28244));
    SB_LUT4 add_3169_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n27775), 
            .O(n6682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_12_lut (.I0(GND_net), .I1(n1949), 
            .I2(VCC_net), .I3(n28463), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_12 (.CI(n28463), .I0(n1949), 
            .I1(VCC_net), .CO(n28464));
    SB_LUT4 div_46_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4388));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_11_lut (.I0(GND_net), .I1(n1950), 
            .I2(VCC_net), .I3(n28462), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_11_lut (.I0(GND_net), .I1(n2450_adj_4233), 
            .I2(VCC_net), .I3(n28242), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_11 (.CI(n28242), .I0(n2450_adj_4233), 
            .I1(VCC_net), .CO(n28243));
    SB_CARRY add_3169_5 (.CI(n27775), .I0(n1173), .I1(n97), .CO(n27776));
    SB_LUT4 add_3169_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n27774), 
            .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_4 (.CI(n27774), .I0(n1174), .I1(n98), .CO(n27775));
    SB_LUT4 communication_counter_31__I_0_add_1653_10_lut (.I0(GND_net), .I1(n2451_adj_4232), 
            .I2(VCC_net), .I3(n28241), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3169_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n27773), 
            .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34115_4_lut (.I0(n29_adj_4443), .I1(n27_adj_4442), .I2(n25_adj_4441), 
            .I3(n40439), .O(n40437));
    defparam i34115_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_46_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4396));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_11 (.CI(n28462), .I0(n1950), 
            .I1(VCC_net), .CO(n28463));
    SB_LUT4 communication_counter_31__I_0_add_1318_10_lut (.I0(GND_net), .I1(n1951), 
            .I2(VCC_net), .I3(n28461), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_10 (.CI(n28241), .I0(n2451_adj_4232), 
            .I1(VCC_net), .CO(n28242));
    SB_LUT4 div_46_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4397));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3169_3 (.CI(n27773), .I0(n1175), .I1(n99), .CO(n27774));
    SB_LUT4 communication_counter_31__I_0_add_1653_9_lut (.I0(GND_net), .I1(n2452_adj_4231), 
            .I2(VCC_net), .I3(n28240), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3169_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3169_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3169_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n27773));
    SB_LUT4 div_46_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4398));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1653_9 (.CI(n28240), .I0(n2452_adj_4231), 
            .I1(VCC_net), .CO(n28241));
    SB_LUT4 div_46_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4394));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3168_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n27772), 
            .O(n6669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_10 (.CI(n28461), .I0(n1951), 
            .I1(VCC_net), .CO(n28462));
    SB_LUT4 communication_counter_31__I_0_add_1653_8_lut (.I0(GND_net), .I1(n2453_adj_4230), 
            .I2(VCC_net), .I3(n28239), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n27771), 
            .O(n6670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4400));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_9_lut (.I0(GND_net), .I1(n1952), 
            .I2(VCC_net), .I3(n28460), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4392));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4401));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_9 (.CI(n28460), .I0(n1952), 
            .I1(VCC_net), .CO(n28461));
    SB_CARRY communication_counter_31__I_0_add_1653_8 (.CI(n28239), .I0(n2453_adj_4230), 
            .I1(VCC_net), .CO(n28240));
    SB_LUT4 div_46_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4402));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_8_lut (.I0(GND_net), .I1(n1953), 
            .I2(VCC_net), .I3(n28459), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_8 (.CI(n28459), .I0(n1953), 
            .I1(VCC_net), .CO(n28460));
    SB_LUT4 div_46_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4403));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_7 (.CI(n27771), .I0(n1044), .I1(n95), .CO(n27772));
    SB_LUT4 communication_counter_31__I_0_add_1653_7_lut (.I0(GND_net), .I1(n2454_adj_4229), 
            .I2(GND_net), .I3(n28238), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n27770), 
            .O(n6671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_7 (.CI(n28238), .I0(n2454_adj_4229), 
            .I1(GND_net), .CO(n28239));
    SB_CARRY add_3168_6 (.CI(n27770), .I0(n1045), .I1(n96), .CO(n27771));
    SB_LUT4 add_3168_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n27769), 
            .O(n6672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_5 (.CI(n27769), .I0(n1046), .I1(n97), .CO(n27770));
    SB_LUT4 add_3168_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n27768), 
            .O(n6673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_6_lut (.I0(GND_net), .I1(n2455_adj_4228), 
            .I2(GND_net), .I3(n28237), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_7_lut (.I0(GND_net), .I1(n1954), 
            .I2(GND_net), .I3(n28458), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4405));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3168_4 (.CI(n27768), .I0(n1047), .I1(n98), .CO(n27769));
    SB_LUT4 div_46_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4406));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4404));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3182_15 (.CI(n28067), .I0(n2541), .I1(n87), .CO(n28068));
    SB_LUT4 add_3168_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n27767), 
            .O(n6674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_3 (.CI(n27767), .I0(n1048), .I1(n99), .CO(n27768));
    SB_LUT4 div_46_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4407));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_7 (.CI(n28458), .I0(n1954), 
            .I1(GND_net), .CO(n28459));
    SB_LUT4 div_46_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4414));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1653_6 (.CI(n28237), .I0(n2455_adj_4228), 
            .I1(GND_net), .CO(n28238));
    SB_LUT4 communication_counter_31__I_0_add_1318_6_lut (.I0(GND_net), .I1(n1955), 
            .I2(GND_net), .I3(n28457), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4424));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1653_5_lut (.I0(GND_net), .I1(n2456_adj_4227), 
            .I2(VCC_net), .I3(n28236), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n27767));
    SB_LUT4 add_3167_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n27766), 
            .O(n6661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n27765), 
            .O(n6662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4417));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1653_5 (.CI(n28236), .I0(n2456_adj_4227), 
            .I1(VCC_net), .CO(n28237));
    SB_CARRY add_3167_6 (.CI(n27765), .I0(n915), .I1(n96), .CO(n27766));
    SB_CARRY communication_counter_31__I_0_add_1318_6 (.CI(n28457), .I0(n1955), 
            .I1(GND_net), .CO(n28458));
    SB_LUT4 div_46_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4416));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4412));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_5_lut (.I0(GND_net), .I1(n1956), 
            .I2(VCC_net), .I3(n28456), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_4_lut (.I0(GND_net), .I1(n2457_adj_4226), 
            .I2(VCC_net), .I3(n28235), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n27764), 
            .O(n6663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4419));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4410));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_5 (.CI(n28456), .I0(n1956), 
            .I1(VCC_net), .CO(n28457));
    SB_CARRY add_3167_5 (.CI(n27764), .I0(n916), .I1(n97), .CO(n27765));
    SB_CARRY communication_counter_31__I_0_add_1653_4 (.CI(n28235), .I0(n2457_adj_4226), 
            .I1(VCC_net), .CO(n28236));
    SB_LUT4 div_46_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4420));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3167_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n27763), 
            .O(n6664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1653_3_lut (.I0(GND_net), .I1(n2458_adj_4225), 
            .I2(GND_net), .I3(n28234), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_4 (.CI(n27763), .I0(n917), .I1(n98), .CO(n27764));
    SB_LUT4 add_3167_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n27762), 
            .O(n6665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4421));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4422));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3167_3 (.CI(n27762), .I0(n918), .I1(n99), .CO(n27763));
    SB_LUT4 div_46_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4425));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_add_1318_4_lut (.I0(GND_net), .I1(n1957), 
            .I2(VCC_net), .I3(n28455), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1653_3 (.CI(n28234), .I0(n2458_adj_4225), 
            .I1(GND_net), .CO(n28235));
    SB_CARRY communication_counter_31__I_0_add_1318_4 (.CI(n28455), .I0(n1957), 
            .I1(VCC_net), .CO(n28456));
    SB_CARRY communication_counter_31__I_0_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4158), 
            .I1(VCC_net), .CO(n28234));
    SB_LUT4 add_3167_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n6666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n27762));
    SB_LUT4 add_6419_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n27761), 
            .O(n10705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4427));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4428));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_6419_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n27760), 
            .O(n10706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1318_3_lut (.I0(GND_net), .I1(n1958), 
            .I2(GND_net), .I3(n28454), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4175), 
            .I2(VCC_net), .I3(n28233), .O(n2636_adj_4138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4423));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_6419_6 (.CI(n27760), .I0(n3354), .I1(GND_net), .CO(n27761));
    SB_LUT4 add_6419_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n27759), 
            .O(n10707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1318_3 (.CI(n28454), .I0(n1958), 
            .I1(GND_net), .CO(n28455));
    SB_LUT4 communication_counter_31__I_0_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4174), 
            .I2(VCC_net), .I3(n28232), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_5 (.CI(n27759), .I0(n3355), .I1(GND_net), .CO(n27760));
    SB_LUT4 div_46_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4429));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY communication_counter_31__I_0_add_1318_2 (.CI(VCC_net), .I0(n2058), 
            .I1(VCC_net), .CO(n28454));
    SB_CARRY communication_counter_31__I_0_add_1720_23 (.CI(n28232), .I0(n2538_adj_4174), 
            .I1(VCC_net), .CO(n28233));
    SB_LUT4 add_6419_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n27758), 
            .O(n10708)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_4 (.CI(n27758), .I0(n3356), .I1(VCC_net), .CO(n27759));
    SB_LUT4 add_6419_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n27757), 
            .O(n10709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4436));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 communication_counter_31__I_0_i1730_3_lut (.I0(n2545_adj_4167), 
            .I1(n2612), .I2(n2570), .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1586_3_lut (.I0(n2360), .I1(n6846), .I2(n2381), .I3(GND_net), 
            .O(n2450));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1729_3_lut (.I0(n2544_adj_4168), 
            .I1(n2611), .I2(n2570), .I3(GND_net), .O(n2643_adj_4120));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6419_3 (.CI(n27757), .I0(n3357), .I1(VCC_net), .CO(n27758));
    SB_LUT4 add_6419_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10710)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6419_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6419_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n27757));
    SB_LUT4 communication_counter_31__I_0_add_1385_19_lut (.I0(n2075_adj_4254), 
            .I1(n2042), .I2(VCC_net), .I3(n28453), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4173), 
            .I2(VCC_net), .I3(n28231), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1385_18_lut (.I0(GND_net), .I1(n2043), 
            .I2(VCC_net), .I3(n28452), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_22 (.CI(n28231), .I0(n2539_adj_4173), 
            .I1(VCC_net), .CO(n28232));
    SB_CARRY communication_counter_31__I_0_add_1385_18 (.CI(n28452), .I0(n2043), 
            .I1(VCC_net), .CO(n28453));
    SB_LUT4 communication_counter_31__I_0_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4172), 
            .I2(VCC_net), .I3(n28230), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1385_17_lut (.I0(GND_net), .I1(n2044), 
            .I2(VCC_net), .I3(n28451), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1385_17 (.CI(n28451), .I0(n2044), 
            .I1(VCC_net), .CO(n28452));
    SB_LUT4 communication_counter_31__I_0_i1728_3_lut (.I0(n2543_adj_4169), 
            .I1(n2610), .I2(n2570), .I3(GND_net), .O(n2642_adj_4134));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1720_21 (.CI(n28230), .I0(n2540_adj_4172), 
            .I1(VCC_net), .CO(n28231));
    SB_LUT4 communication_counter_31__I_0_add_1385_16_lut (.I0(GND_net), .I1(n2045), 
            .I2(VCC_net), .I3(n28450), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1385_16 (.CI(n28450), .I0(n2045), 
            .I1(VCC_net), .CO(n28451));
    SB_LUT4 communication_counter_31__I_0_add_1385_15_lut (.I0(GND_net), .I1(n2046), 
            .I2(VCC_net), .I3(n28449), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4171), 
            .I2(VCC_net), .I3(n28229), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1385_15 (.CI(n28449), .I0(n2046), 
            .I1(VCC_net), .CO(n28450));
    SB_CARRY communication_counter_31__I_0_add_1720_20 (.CI(n28229), .I0(n2541_adj_4171), 
            .I1(VCC_net), .CO(n28230));
    SB_LUT4 communication_counter_31__I_0_add_1385_14_lut (.I0(GND_net), .I1(n2047), 
            .I2(VCC_net), .I3(n28448), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1735_3_lut (.I0(n2550_adj_4162), 
            .I1(n2617), .I2(n2570), .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1385_14 (.CI(n28448), .I0(n2047), 
            .I1(VCC_net), .CO(n28449));
    SB_LUT4 communication_counter_31__I_0_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4170), 
            .I2(VCC_net), .I3(n28228), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_19 (.CI(n28228), .I0(n2542_adj_4170), 
            .I1(VCC_net), .CO(n28229));
    SB_LUT4 communication_counter_31__I_0_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4169), 
            .I2(VCC_net), .I3(n28227), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1385_13_lut (.I0(GND_net), .I1(n2048), 
            .I2(VCC_net), .I3(n28447), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1732_3_lut (.I0(n2547_adj_4165), 
            .I1(n2614), .I2(n2570), .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1385_13 (.CI(n28447), .I0(n2048), 
            .I1(VCC_net), .CO(n28448));
    SB_LUT4 communication_counter_31__I_0_add_1385_12_lut (.I0(GND_net), .I1(n2049), 
            .I2(VCC_net), .I3(n28446), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_18 (.CI(n28227), .I0(n2543_adj_4169), 
            .I1(VCC_net), .CO(n28228));
    SB_CARRY communication_counter_31__I_0_add_1385_12 (.CI(n28446), .I0(n2049), 
            .I1(VCC_net), .CO(n28447));
    SB_LUT4 i33351_4_lut (.I0(n35_adj_4446), .I1(n33_adj_4445), .I2(n31_adj_4444), 
            .I3(n40437), .O(n39673));
    defparam i33351_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 communication_counter_31__I_0_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4168), 
            .I2(VCC_net), .I3(n28226), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1385_11_lut (.I0(GND_net), .I1(n2050), 
            .I2(VCC_net), .I3(n28445), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_17 (.CI(n28226), .I0(n2544_adj_4168), 
            .I1(VCC_net), .CO(n28227));
    SB_CARRY communication_counter_31__I_0_add_1385_11 (.CI(n28445), .I0(n2050), 
            .I1(VCC_net), .CO(n28446));
    SB_LUT4 communication_counter_31__I_0_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4167), 
            .I2(VCC_net), .I3(n28225), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1606_i12_4_lut (.I0(n387), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4430));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_i1769_3_lut_3_lut (.I0(n2642), .I1(n6924), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_add_1385_10_lut (.I0(GND_net), .I1(n2051), 
            .I2(VCC_net), .I3(n28444), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_16 (.CI(n28225), .I0(n2545_adj_4167), 
            .I1(VCC_net), .CO(n28226));
    SB_LUT4 div_46_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4217));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_1385_10 (.CI(n28444), .I0(n2051), 
            .I1(VCC_net), .CO(n28445));
    SB_LUT4 communication_counter_31__I_0_add_1385_9_lut (.I0(GND_net), .I1(n2052), 
            .I2(VCC_net), .I3(n28443), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4166), 
            .I2(VCC_net), .I3(n28224), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_15 (.CI(n28224), .I0(n2546_adj_4166), 
            .I1(VCC_net), .CO(n28225));
    SB_LUT4 communication_counter_31__I_0_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4165), 
            .I2(VCC_net), .I3(n28223), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13330_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n24632), 
            .I3(n16424), .O(n17837));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13330_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY communication_counter_31__I_0_add_1720_14 (.CI(n28223), .I0(n2547_adj_4165), 
            .I1(VCC_net), .CO(n28224));
    SB_CARRY communication_counter_31__I_0_add_1385_9 (.CI(n28443), .I0(n2052), 
            .I1(VCC_net), .CO(n28444));
    SB_LUT4 communication_counter_31__I_0_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4164), 
            .I2(VCC_net), .I3(n28222), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_13 (.CI(n28222), .I0(n2548_adj_4164), 
            .I1(VCC_net), .CO(n28223));
    SB_LUT4 communication_counter_31__I_0_add_1385_8_lut (.I0(GND_net), .I1(n2053), 
            .I2(VCC_net), .I3(n28442), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13331_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n24632), 
            .I3(n16429), .O(n17838));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13331_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY communication_counter_31__I_0_add_1385_8 (.CI(n28442), .I0(n2053), 
            .I1(VCC_net), .CO(n28443));
    SB_LUT4 communication_counter_31__I_0_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4163), 
            .I2(VCC_net), .I3(n28221), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_12 (.CI(n28221), .I0(n2549_adj_4163), 
            .I1(VCC_net), .CO(n28222));
    SB_LUT4 communication_counter_31__I_0_add_1385_7_lut (.I0(GND_net), .I1(n2054), 
            .I2(GND_net), .I3(n28441), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4162), 
            .I2(VCC_net), .I3(n28220), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_11 (.CI(n28220), .I0(n2550_adj_4162), 
            .I1(VCC_net), .CO(n28221));
    SB_CARRY communication_counter_31__I_0_add_1385_7 (.CI(n28441), .I0(n2054), 
            .I1(GND_net), .CO(n28442));
    SB_LUT4 div_46_i1754_3_lut_3_lut (.I0(n2642), .I1(n6909), .I2(n2618), 
            .I3(GND_net), .O(n2699_adj_4065));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4216));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_1385_6_lut (.I0(GND_net), .I1(n2055), 
            .I2(GND_net), .I3(n28440), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13332_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n16424), 
            .O(n17839));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13332_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY communication_counter_31__I_0_add_1385_6 (.CI(n28440), .I0(n2055), 
            .I1(GND_net), .CO(n28441));
    SB_LUT4 communication_counter_31__I_0_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4161), 
            .I2(VCC_net), .I3(n28219), .O(n2618_adj_4146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1737_3_lut (.I0(n2552_adj_4160), 
            .I1(n2619_adj_4145), .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13333_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n16429), 
            .O(n17840));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13333_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 communication_counter_31__I_0_add_1385_5_lut (.I0(GND_net), .I1(n2056), 
            .I2(VCC_net), .I3(n28439), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13334_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4022), 
            .I3(n16424), .O(n17841));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13334_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY communication_counter_31__I_0_add_1720_10 (.CI(n28219), .I0(n2551_adj_4161), 
            .I1(VCC_net), .CO(n28220));
    SB_CARRY communication_counter_31__I_0_add_1385_5 (.CI(n28439), .I0(n2056), 
            .I1(VCC_net), .CO(n28440));
    SB_LUT4 communication_counter_31__I_0_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4160), 
            .I2(VCC_net), .I3(n28218), .O(n2619_adj_4145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_9 (.CI(n28218), .I0(n2552_adj_4160), 
            .I1(VCC_net), .CO(n28219));
    SB_LUT4 div_46_i1755_3_lut_3_lut (.I0(n2642), .I1(n6910), .I2(n2619), 
            .I3(GND_net), .O(n2700_adj_4066));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1731_3_lut (.I0(n2546_adj_4166), 
            .I1(n2613), .I2(n2570), .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13335_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4022), 
            .I3(n16429), .O(n17842));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13335_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 communication_counter_31__I_0_add_1385_4_lut (.I0(GND_net), .I1(n2057), 
            .I2(VCC_net), .I3(n28438), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4159), 
            .I2(VCC_net), .I3(n28217), .O(n2620_adj_4144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1723_3_lut (.I0(n2538_adj_4174), 
            .I1(n2605), .I2(n2570), .I3(GND_net), .O(n2637_adj_4137));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1385_4 (.CI(n28438), .I0(n2057), 
            .I1(VCC_net), .CO(n28439));
    SB_CARRY communication_counter_31__I_0_add_1720_8 (.CI(n28217), .I0(n2553_adj_4159), 
            .I1(VCC_net), .CO(n28218));
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_205[23]), 
            .I2(n3_adj_3984), .I3(n27713), .O(displacement_23__N_81[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4215));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_205[22]), 
            .I2(n3_adj_3984), .I3(n27712), .O(displacement_23__N_81[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n27712), .I0(displacement_23__N_205[22]), 
            .I1(n3_adj_3984), .CO(n27713));
    SB_LUT4 communication_counter_31__I_0_add_1385_3_lut (.I0(GND_net), .I1(n2058), 
            .I2(GND_net), .I3(n28437), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_7_lut (.I0(GND_net), .I1(n2554), 
            .I2(GND_net), .I3(n28216), .O(n2621_adj_4143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1736_3_lut (.I0(n2551_adj_4161), 
            .I1(n2618_adj_4146), .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1385_3 (.CI(n28437), .I0(n2058), 
            .I1(GND_net), .CO(n28438));
    SB_LUT4 communication_counter_31__I_0_i1743_3_lut (.I0(n2558_adj_4158), 
            .I1(n2625_adj_4139), .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4141), 
            .I2(n2570), .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1720_7 (.CI(n28216), .I0(n2554), 
            .I1(GND_net), .CO(n28217));
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_205[21]), 
            .I2(n3_adj_3984), .I3(n27711), .O(displacement_23__N_81[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4142), 
            .I2(n2570), .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n27711), .I0(displacement_23__N_205[21]), 
            .I1(n3_adj_3984), .CO(n27712));
    SB_CARRY communication_counter_31__I_0_add_1385_2 (.CI(VCC_net), .I0(n2158), 
            .I1(VCC_net), .CO(n28437));
    SB_LUT4 communication_counter_31__I_0_i1733_3_lut (.I0(n2548_adj_4164), 
            .I1(n2615), .I2(n2570), .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1720_6_lut (.I0(GND_net), .I1(n2555), 
            .I2(GND_net), .I3(n28215), .O(n2622_adj_4142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1452_20_lut (.I0(n2174_adj_4245), 
            .I1(n2141), .I2(VCC_net), .I3(n28436), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_205[20]), 
            .I2(n3_adj_3984), .I3(n27710), .O(displacement_23__N_81[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_6 (.CI(n28215), .I0(n2555), 
            .I1(GND_net), .CO(n28216));
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n27710), .I0(displacement_23__N_205[20]), 
            .I1(n3_adj_3984), .CO(n27711));
    SB_LUT4 communication_counter_31__I_0_add_1452_19_lut (.I0(GND_net), .I1(n2142), 
            .I2(VCC_net), .I3(n28435), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_205[19]), 
            .I2(n6_adj_3934), .I3(n27709), .O(displacement_23__N_81[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1452_19 (.CI(n28435), .I0(n2142), 
            .I1(VCC_net), .CO(n28436));
    SB_LUT4 communication_counter_31__I_0_add_1720_5_lut (.I0(GND_net), .I1(n2556), 
            .I2(VCC_net), .I3(n28214), .O(n2623_adj_4141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n27709), .I0(displacement_23__N_205[19]), 
            .I1(n6_adj_3934), .CO(n27710));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_205[18]), 
            .I2(n7), .I3(n27708), .O(displacement_23__N_81[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n27708), .I0(displacement_23__N_205[18]), 
            .I1(n7), .CO(n27709));
    SB_LUT4 communication_counter_31__I_0_add_1452_18_lut (.I0(GND_net), .I1(n2143), 
            .I2(VCC_net), .I3(n28434), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_5 (.CI(n28214), .I0(n2556), 
            .I1(VCC_net), .CO(n28215));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_205[17]), 
            .I2(n8_adj_4024), .I3(n27707), .O(displacement_23__N_81[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n27707), .I0(displacement_23__N_205[17]), 
            .I1(n8_adj_4024), .CO(n27708));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_205[16]), 
            .I2(n9_adj_4025), .I3(n27706), .O(displacement_23__N_81[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n27706), .I0(displacement_23__N_205[16]), 
            .I1(n9_adj_4025), .CO(n27707));
    SB_LUT4 div_46_i1756_3_lut_3_lut (.I0(n2642), .I1(n6911), .I2(n2620), 
            .I3(GND_net), .O(n2701_adj_4067));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1757_3_lut_3_lut (.I0(n2642), .I1(n6912), .I2(n2621), 
            .I3(GND_net), .O(n2702_adj_4068));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_31__I_0_add_1452_18 (.CI(n28434), .I0(n2143), 
            .I1(VCC_net), .CO(n28435));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_205[15]), 
            .I2(n10_adj_4026), .I3(n27705), .O(displacement_23__N_81[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1452_17_lut (.I0(GND_net), .I1(n2144), 
            .I2(VCC_net), .I3(n28433), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_4_lut (.I0(GND_net), .I1(n2557), 
            .I2(VCC_net), .I3(n28213), .O(n2624_adj_4140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4214));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n27705), .I0(displacement_23__N_205[15]), 
            .I1(n10_adj_4026), .CO(n27706));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_205[14]), 
            .I2(n11_adj_4027), .I3(n27704), .O(displacement_23__N_81[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_4 (.CI(n28213), .I0(n2557), 
            .I1(VCC_net), .CO(n28214));
    SB_CARRY communication_counter_31__I_0_add_1452_17 (.CI(n28433), .I0(n2144), 
            .I1(VCC_net), .CO(n28434));
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n27704), .I0(displacement_23__N_205[14]), 
            .I1(n11_adj_4027), .CO(n27705));
    SB_LUT4 communication_counter_31__I_0_add_1452_16_lut (.I0(GND_net), .I1(n2145), 
            .I2(VCC_net), .I3(n28432), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4158), 
            .I2(GND_net), .I3(n28212), .O(n2625_adj_4139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1720_3 (.CI(n28212), .I0(n2558_adj_4158), 
            .I1(GND_net), .CO(n28213));
    SB_LUT4 i13336_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4023), 
            .I3(n16424), .O(n17843));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13336_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY communication_counter_31__I_0_add_1452_16 (.CI(n28432), .I0(n2145), 
            .I1(VCC_net), .CO(n28433));
    SB_CARRY communication_counter_31__I_0_add_1720_2 (.CI(VCC_net), .I0(n2658), 
            .I1(VCC_net), .CO(n28212));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_205[13]), 
            .I2(n12_adj_4028), .I3(n27703), .O(displacement_23__N_81[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n27703), .I0(displacement_23__N_205[13]), 
            .I1(n12_adj_4028), .CO(n27704));
    SB_LUT4 communication_counter_31__I_0_add_1452_15_lut (.I0(GND_net), .I1(n2146), 
            .I2(VCC_net), .I3(n28431), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_25_lut (.I0(n2669), .I1(n2636_adj_4138), 
            .I2(VCC_net), .I3(n28211), .O(n2735_adj_4099)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_i1739_3_lut (.I0(n2554), .I1(n2621_adj_4143), 
            .I2(n2570), .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1452_15 (.CI(n28431), .I0(n2146), 
            .I1(VCC_net), .CO(n28432));
    SB_LUT4 communication_counter_31__I_0_i1734_3_lut (.I0(n2549_adj_4163), 
            .I1(n2616), .I2(n2570), .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1787_24_lut (.I0(GND_net), .I1(n2637_adj_4137), 
            .I2(VCC_net), .I3(n28210), .O(n2704_adj_4118)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_205[12]), 
            .I2(n13_adj_4029), .I3(n27702), .O(displacement_23__N_81[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n27702), .I0(displacement_23__N_205[12]), 
            .I1(n13_adj_4029), .CO(n27703));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_205[11]), 
            .I2(n14_adj_4030), .I3(n27701), .O(displacement_23__N_81[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1452_14_lut (.I0(GND_net), .I1(n2147), 
            .I2(VCC_net), .I3(n28430), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_24 (.CI(n28210), .I0(n2637_adj_4137), 
            .I1(VCC_net), .CO(n28211));
    SB_LUT4 div_46_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4213));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n27701), .I0(displacement_23__N_205[11]), 
            .I1(n14_adj_4030), .CO(n27702));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_205[10]), 
            .I2(n15_adj_4031), .I3(n27700), .O(displacement_23__N_81[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n27700), .I0(displacement_23__N_205[10]), 
            .I1(n15_adj_4031), .CO(n27701));
    SB_LUT4 div_46_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4212));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_205[9]), 
            .I2(n16_adj_4032), .I3(n27699), .O(displacement_23__N_81[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n27699), .I0(displacement_23__N_205[9]), 
            .I1(n16_adj_4032), .CO(n27700));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_205[8]), 
            .I2(n17_adj_4033), .I3(n27698), .O(displacement_23__N_81[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n27698), .I0(displacement_23__N_205[8]), 
            .I1(n17_adj_4033), .CO(n27699));
    SB_LUT4 communication_counter_31__I_0_i1738_3_lut (.I0(n2553_adj_4159), 
            .I1(n2620_adj_4144), .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1452_14 (.CI(n28430), .I0(n2147), 
            .I1(VCC_net), .CO(n28431));
    SB_LUT4 communication_counter_31__I_0_add_1787_23_lut (.I0(GND_net), .I1(n2638_adj_4136), 
            .I2(VCC_net), .I3(n28209), .O(n2705_adj_4117)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1452_13_lut (.I0(GND_net), .I1(n2148), 
            .I2(VCC_net), .I3(n28429), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_205[7]), 
            .I2(n18_adj_4034), .I3(n27697), .O(displacement_23__N_81[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n27697), .I0(displacement_23__N_205[7]), 
            .I1(n18_adj_4034), .CO(n27698));
    SB_CARRY communication_counter_31__I_0_add_1452_13 (.CI(n28429), .I0(n2148), 
            .I1(VCC_net), .CO(n28430));
    SB_LUT4 communication_counter_31__I_0_add_1452_12_lut (.I0(GND_net), .I1(n2149), 
            .I2(VCC_net), .I3(n28428), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1452_12 (.CI(n28428), .I0(n2149), 
            .I1(VCC_net), .CO(n28429));
    SB_LUT4 communication_counter_31__I_0_add_1452_11_lut (.I0(GND_net), .I1(n2150), 
            .I2(VCC_net), .I3(n28427), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_23 (.CI(n28209), .I0(n2638_adj_4136), 
            .I1(VCC_net), .CO(n28210));
    SB_CARRY communication_counter_31__I_0_add_1452_11 (.CI(n28427), .I0(n2150), 
            .I1(VCC_net), .CO(n28428));
    SB_LUT4 communication_counter_31__I_0_add_1787_22_lut (.I0(GND_net), .I1(n2639), 
            .I2(VCC_net), .I3(n28208), .O(n2706_adj_4116)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_205[6]), 
            .I2(n19_adj_4035), .I3(n27696), .O(displacement_23__N_81[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34169_3_lut (.I0(n12_adj_4430), .I1(n87), .I2(n35_adj_4446), 
            .I3(GND_net), .O(n40491));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34169_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n27696), .I0(displacement_23__N_205[6]), 
            .I1(n19_adj_4035), .CO(n27697));
    SB_LUT4 i13693_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13950), 
            .I3(GND_net), .O(n18200));   // verilog/coms.v(126[12] 289[6])
    defparam i13693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_205[5]), 
            .I2(n20_adj_4036), .I3(n27695), .O(displacement_23__N_81[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4211));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4210));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_add_1452_10_lut (.I0(GND_net), .I1(n2151), 
            .I2(VCC_net), .I3(n28426), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_22 (.CI(n28208), .I0(n2639), 
            .I1(VCC_net), .CO(n28209));
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n27695), .I0(displacement_23__N_205[5]), 
            .I1(n20_adj_4036), .CO(n27696));
    SB_LUT4 div_46_i1531_3_lut (.I0(n2273), .I1(n6832), .I2(n2288), .I3(GND_net), 
            .O(n2366));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1531_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_205[4]), 
            .I2(n21_adj_4037), .I3(n27694), .O(displacement_23__N_81[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_21_lut (.I0(GND_net), .I1(n2640), 
            .I2(VCC_net), .I3(n28207), .O(n2707_adj_4115)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_21 (.CI(n28207), .I0(n2640), 
            .I1(VCC_net), .CO(n28208));
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n27694), .I0(displacement_23__N_205[4]), 
            .I1(n21_adj_4037), .CO(n27695));
    SB_CARRY communication_counter_31__I_0_add_1452_10 (.CI(n28426), .I0(n2151), 
            .I1(VCC_net), .CO(n28427));
    SB_LUT4 communication_counter_31__I_0_add_1787_20_lut (.I0(GND_net), .I1(n2641), 
            .I2(VCC_net), .I3(n28206), .O(n2708_adj_4114)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_205[3]), 
            .I2(n22_adj_4038), .I3(n27693), .O(displacement_23__N_81[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n27693), .I0(displacement_23__N_205[3]), 
            .I1(n22_adj_4038), .CO(n27694));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_205[2]), 
            .I2(n23_adj_4039), .I3(n27692), .O(displacement_23__N_81[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1452_9_lut (.I0(GND_net), .I1(n2152), 
            .I2(VCC_net), .I3(n28425), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_20 (.CI(n28206), .I0(n2641), 
            .I1(VCC_net), .CO(n28207));
    SB_CARRY communication_counter_31__I_0_add_1452_9 (.CI(n28425), .I0(n2152), 
            .I1(VCC_net), .CO(n28426));
    SB_LUT4 communication_counter_31__I_0_add_1787_19_lut (.I0(GND_net), .I1(n2642_adj_4134), 
            .I2(VCC_net), .I3(n28205), .O(n2709_adj_4113)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n27692), .I0(displacement_23__N_205[2]), 
            .I1(n23_adj_4039), .CO(n27693));
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_205[1]), 
            .I2(n24_adj_4040), .I3(n27691), .O(displacement_23__N_81[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n27691), .I0(displacement_23__N_205[1]), 
            .I1(n24_adj_4040), .CO(n27692));
    SB_LUT4 div_46_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4209));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_205[0]), 
            .I2(n25_adj_4041), .I3(VCC_net), .O(displacement_23__N_81[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_205[0]), 
            .I1(n25_adj_4041), .CO(n27691));
    SB_LUT4 i13694_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13950), 
            .I3(GND_net), .O(n18201));   // verilog/coms.v(126[12] 289[6])
    defparam i13694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1452_8_lut (.I0(GND_net), .I1(n2153), 
            .I2(VCC_net), .I3(n28424), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_mux_3_i10_3_lut (.I0(communication_counter[9]), 
            .I1(n24_adj_3961), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2658));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1758_3_lut_3_lut (.I0(n2642), .I1(n6913), .I2(n2622), 
            .I3(GND_net), .O(n2703_adj_4069));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4208));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4140), 
            .I2(n2570), .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1662_3_lut (.I0(n2445), .I1(n2512), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2544_adj_4168));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4207));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_31__I_0_add_1452_8 (.CI(n28424), .I0(n2153), 
            .I1(VCC_net), .CO(n28425));
    SB_CARRY communication_counter_31__I_0_add_1787_19 (.CI(n28205), .I0(n2642_adj_4134), 
            .I1(VCC_net), .CO(n28206));
    SB_LUT4 communication_counter_31__I_0_add_1787_18_lut (.I0(GND_net), .I1(n2643_adj_4120), 
            .I2(VCC_net), .I3(n28204), .O(n2710_adj_4112)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1761_3_lut_3_lut (.I0(n2642), .I1(n6916), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1661_3_lut (.I0(n2444), .I1(n2511), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2543_adj_4169));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4206));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1659_3_lut (.I0(n2442), .I1(n2509), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2541_adj_4171));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1671_3_lut (.I0(n2454_adj_4229), 
            .I1(n2521), .I2(n2471_adj_4224), .I3(GND_net), .O(n2553_adj_4159));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1663_3_lut (.I0(n2446), .I1(n2513), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2545_adj_4167));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1664_3_lut (.I0(n2447_adj_4236), 
            .I1(n2514), .I2(n2471_adj_4224), .I3(GND_net), .O(n2546_adj_4166));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1668_3_lut (.I0(n2451_adj_4232), 
            .I1(n2518), .I2(n2471_adj_4224), .I3(GND_net), .O(n2550_adj_4162));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1452_7_lut (.I0(GND_net), .I1(n2154), 
            .I2(GND_net), .I3(n28423), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_18 (.CI(n28204), .I0(n2643_adj_4120), 
            .I1(VCC_net), .CO(n28205));
    SB_CARRY communication_counter_31__I_0_add_1452_7 (.CI(n28423), .I0(n2154), 
            .I1(GND_net), .CO(n28424));
    SB_LUT4 communication_counter_31__I_0_add_1452_6_lut (.I0(GND_net), .I1(n2155), 
            .I2(GND_net), .I3(n28422), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_17_lut (.I0(GND_net), .I1(n2644), 
            .I2(VCC_net), .I3(n28203), .O(n2711_adj_4111)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1452_6 (.CI(n28422), .I0(n2155), 
            .I1(GND_net), .CO(n28423));
    SB_CARRY communication_counter_31__I_0_add_1787_17 (.CI(n28203), .I0(n2644), 
            .I1(VCC_net), .CO(n28204));
    SB_LUT4 communication_counter_31__I_0_i1670_3_lut (.I0(n2453_adj_4230), 
            .I1(n2520), .I2(n2471_adj_4224), .I3(GND_net), .O(n2552_adj_4160));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1452_5_lut (.I0(GND_net), .I1(n2156), 
            .I2(VCC_net), .I3(n28421), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_16_lut (.I0(GND_net), .I1(n2645), 
            .I2(VCC_net), .I3(n28202), .O(n2712_adj_4110)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_16 (.CI(n28202), .I0(n2645), 
            .I1(VCC_net), .CO(n28203));
    SB_CARRY communication_counter_31__I_0_add_1452_5 (.CI(n28421), .I0(n2156), 
            .I1(VCC_net), .CO(n28422));
    SB_LUT4 communication_counter_31__I_0_add_1452_4_lut (.I0(GND_net), .I1(n2157), 
            .I2(VCC_net), .I3(n28420), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_15_lut (.I0(GND_net), .I1(n2646), 
            .I2(VCC_net), .I3(n28201), .O(n2713_adj_4109)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1762_3_lut_3_lut (.I0(n2642), .I1(n6917), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_31__I_0_add_1452_4 (.CI(n28420), .I0(n2157), 
            .I1(VCC_net), .CO(n28421));
    SB_CARRY communication_counter_31__I_0_add_1787_15 (.CI(n28201), .I0(n2646), 
            .I1(VCC_net), .CO(n28202));
    SB_LUT4 div_46_i1759_3_lut_3_lut (.I0(n2642), .I1(n6914), .I2(n2623), 
            .I3(GND_net), .O(n2704_adj_4070));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_add_1452_3_lut (.I0(GND_net), .I1(n2158), 
            .I2(GND_net), .I3(n28419), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_14_lut (.I0(GND_net), .I1(n2647), 
            .I2(VCC_net), .I3(n28200), .O(n2714_adj_4108)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i1669_3_lut (.I0(n2452_adj_4231), 
            .I1(n2519), .I2(n2471_adj_4224), .I3(GND_net), .O(n2551_adj_4161));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1452_3 (.CI(n28419), .I0(n2158), 
            .I1(GND_net), .CO(n28420));
    SB_CARRY communication_counter_31__I_0_add_1787_14 (.CI(n28200), .I0(n2647), 
            .I1(VCC_net), .CO(n28201));
    SB_LUT4 communication_counter_31__I_0_i1666_3_lut (.I0(n2449_adj_4234), 
            .I1(n2516), .I2(n2471_adj_4224), .I3(GND_net), .O(n2548_adj_4164));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1452_2 (.CI(VCC_net), .I0(n2258), 
            .I1(VCC_net), .CO(n28419));
    SB_LUT4 div_46_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4200), .I3(n28418), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_31__I_0_add_1787_13_lut (.I0(GND_net), .I1(n2648), 
            .I2(VCC_net), .I3(n28199), .O(n2715_adj_4107)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4205));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4201), .I3(n28417), .O(n3_adj_4012)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_13 (.CI(n28199), .I0(n2648), 
            .I1(VCC_net), .CO(n28200));
    SB_CARRY div_46_unary_minus_2_add_3_24 (.CI(n28417), .I0(GND_net), .I1(n3_adj_4201), 
            .CO(n28418));
    SB_LUT4 communication_counter_31__I_0_add_1787_12_lut (.I0(GND_net), .I1(n2649), 
            .I2(VCC_net), .I3(n28198), .O(n2716_adj_4106)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4202), .I3(n28416), .O(n4_adj_4007)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_12 (.CI(n28198), .I0(n2649), 
            .I1(VCC_net), .CO(n28199));
    SB_LUT4 communication_counter_31__I_0_add_1787_11_lut (.I0(GND_net), .I1(n2650), 
            .I2(VCC_net), .I3(n28197), .O(n2717_adj_4105)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_23 (.CI(n28416), .I0(GND_net), .I1(n4_adj_4202), 
            .CO(n28417));
    SB_LUT4 div_46_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4203), .I3(n28415), .O(n5_adj_4006)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_11 (.CI(n28197), .I0(n2650), 
            .I1(VCC_net), .CO(n28198));
    SB_LUT4 communication_counter_31__I_0_add_1787_10_lut (.I0(GND_net), .I1(n2651), 
            .I2(VCC_net), .I3(n28196), .O(n2718_adj_4104)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_22 (.CI(n28415), .I0(GND_net), .I1(n5_adj_4203), 
            .CO(n28416));
    SB_LUT4 div_46_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4204), .I3(n28414), .O(n6_adj_4005)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_10 (.CI(n28196), .I0(n2651), 
            .I1(VCC_net), .CO(n28197));
    SB_CARRY div_46_unary_minus_2_add_3_21 (.CI(n28414), .I0(GND_net), .I1(n6_adj_4204), 
            .CO(n28415));
    SB_LUT4 communication_counter_31__I_0_add_1787_9_lut (.I0(GND_net), .I1(n2652), 
            .I2(VCC_net), .I3(n28195), .O(n2719_adj_4103)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4205), .I3(n28413), .O(n7_adj_4004)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_9 (.CI(n28195), .I0(n2652), 
            .I1(VCC_net), .CO(n28196));
    SB_LUT4 div_46_i1760_3_lut_3_lut (.I0(n2642), .I1(n6915), .I2(n2624), 
            .I3(GND_net), .O(n2705_adj_4071));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4204));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1667_3_lut (.I0(n2450_adj_4233), 
            .I1(n2517), .I2(n2471_adj_4224), .I3(GND_net), .O(n2549_adj_4163));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_20 (.CI(n28413), .I0(GND_net), .I1(n7_adj_4205), 
            .CO(n28414));
    SB_LUT4 div_46_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4203));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13695_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13950), 
            .I3(GND_net), .O(n18202));   // verilog/coms.v(126[12] 289[6])
    defparam i13695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1665_3_lut (.I0(n2448_adj_4235), 
            .I1(n2515), .I2(n2471_adj_4224), .I3(GND_net), .O(n2547_adj_4165));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1787_8_lut (.I0(GND_net), .I1(n2653), 
            .I2(VCC_net), .I3(n28194), .O(n2720_adj_4102)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_8 (.CI(n28194), .I0(n2653), 
            .I1(VCC_net), .CO(n28195));
    SB_LUT4 communication_counter_31__I_0_add_1787_7_lut (.I0(GND_net), .I1(n2654), 
            .I2(GND_net), .I3(n28193), .O(n2721)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_7 (.CI(n28193), .I0(n2654), 
            .I1(GND_net), .CO(n28194));
    SB_LUT4 i13696_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13950), 
            .I3(GND_net), .O(n18203));   // verilog/coms.v(126[12] 289[6])
    defparam i13696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4206), .I3(n28412), .O(n8_adj_4003)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13697_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13950), 
            .I3(GND_net), .O(n18204));   // verilog/coms.v(126[12] 289[6])
    defparam i13697_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_19 (.CI(n28412), .I0(GND_net), .I1(n8_adj_4206), 
            .CO(n28413));
    SB_LUT4 communication_counter_31__I_0_add_1787_6_lut (.I0(GND_net), .I1(n2655), 
            .I2(GND_net), .I3(n28192), .O(n2722)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_6 (.CI(n28192), .I0(n2655), 
            .I1(GND_net), .CO(n28193));
    SB_LUT4 div_46_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4207), .I3(n28411), .O(n9_adj_4002)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_18 (.CI(n28411), .I0(GND_net), .I1(n9_adj_4207), 
            .CO(n28412));
    SB_LUT4 communication_counter_31__I_0_mux_3_i11_3_lut (.I0(communication_counter[10]), 
            .I1(n23_adj_3962), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2558_adj_4158));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4208), .I3(n28410), .O(n10_adj_4001)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_17 (.CI(n28410), .I0(GND_net), .I1(n10_adj_4208), 
            .CO(n28411));
    SB_LUT4 communication_counter_31__I_0_add_1787_5_lut (.I0(GND_net), .I1(n2656), 
            .I2(VCC_net), .I3(n28191), .O(n2723_adj_4101)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4209), .I3(n28409), .O(n11_adj_4000)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1787_5 (.CI(n28191), .I0(n2656), 
            .I1(VCC_net), .CO(n28192));
    SB_CARRY div_46_unary_minus_2_add_3_16 (.CI(n28409), .I0(GND_net), .I1(n11_adj_4209), 
            .CO(n28410));
    SB_LUT4 div_46_LessThan_1606_i38_3_lut (.I0(n20_adj_4437), .I1(n83), 
            .I2(n43_adj_4451), .I3(GND_net), .O(n38_adj_4448));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 communication_counter_31__I_0_add_1787_4_lut (.I0(GND_net), .I1(n2657), 
            .I2(VCC_net), .I3(n28190), .O(n2724_adj_4100)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4210), .I3(n28408), .O(n12_adj_3999)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1674_3_lut (.I0(n2457_adj_4226), 
            .I1(n2524), .I2(n2471_adj_4224), .I3(GND_net), .O(n2556));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4202));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_46_unary_minus_2_add_3_15 (.CI(n28408), .I0(GND_net), .I1(n12_adj_4210), 
            .CO(n28409));
    SB_LUT4 div_46_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4211), .I3(n28407), .O(n13_adj_3998)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1675_3_lut (.I0(n2458_adj_4225), 
            .I1(n2525), .I2(n2471_adj_4224), .I3(GND_net), .O(n2557));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_14 (.CI(n28407), .I0(GND_net), .I1(n13_adj_4211), 
            .CO(n28408));
    SB_LUT4 div_46_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4212), .I3(n28406), .O(n14_adj_3997)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_13 (.CI(n28406), .I0(GND_net), .I1(n14_adj_4212), 
            .CO(n28407));
    SB_LUT4 div_46_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4201));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4213), .I3(n28405), .O(n15_adj_3996)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13698_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13950), 
            .I3(GND_net), .O(n18205));   // verilog/coms.v(126[12] 289[6])
    defparam i13698_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1787_4 (.CI(n28190), .I0(n2657), 
            .I1(VCC_net), .CO(n28191));
    SB_LUT4 div_46_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4200));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1673_3_lut (.I0(n2456_adj_4227), 
            .I1(n2523), .I2(n2471_adj_4224), .I3(GND_net), .O(n2555));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1672_3_lut (.I0(n2455_adj_4228), 
            .I1(n2522), .I2(n2471_adj_4224), .I3(GND_net), .O(n2554));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1775_3_lut_3_lut (.I0(n2642), .I1(n6930), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1592_3_lut (.I0(n2343), .I1(n2410), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_12 (.CI(n28405), .I0(GND_net), .I1(n15_adj_4213), 
            .CO(n28406));
    SB_LUT4 div_46_i1764_3_lut_3_lut (.I0(n2642), .I1(n6919), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4214), .I3(n28404), .O(n16_adj_3995)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1787_3_lut (.I0(GND_net), .I1(n2658), 
            .I2(GND_net), .I3(n28189), .O(n2725)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1787_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1597_3_lut (.I0(n2348), .I1(n2415), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2447_adj_4236));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13699_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13950), 
            .I3(GND_net), .O(n18206));   // verilog/coms.v(126[12] 289[6])
    defparam i13699_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_11 (.CI(n28404), .I0(GND_net), .I1(n16_adj_4214), 
            .CO(n28405));
    SB_LUT4 i13700_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13950), 
            .I3(GND_net), .O(n18207));   // verilog/coms.v(126[12] 289[6])
    defparam i13700_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1787_3 (.CI(n28189), .I0(n2658), 
            .I1(GND_net), .CO(n28190));
    SB_LUT4 i13701_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13950), 
            .I3(GND_net), .O(n18208));   // verilog/coms.v(126[12] 289[6])
    defparam i13701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13702_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13950), 
            .I3(GND_net), .O(n18209));   // verilog/coms.v(126[12] 289[6])
    defparam i13702_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_31__I_0_add_1787_2 (.CI(VCC_net), .I0(n2758), 
            .I1(VCC_net), .CO(n28189));
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4041));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4215), .I3(n28403), .O(n17_adj_3994)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13703_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13950), 
            .I3(GND_net), .O(n18210));   // verilog/coms.v(126[12] 289[6])
    defparam i13703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1854_25_lut (.I0(n2768), .I1(n2735_adj_4099), 
            .I2(VCC_net), .I3(n28188), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4040));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13704_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13950), 
            .I3(GND_net), .O(n18211));   // verilog/coms.v(126[12] 289[6])
    defparam i13704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4039));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_46_unary_minus_2_add_3_10 (.CI(n28403), .I0(GND_net), .I1(n17_adj_4215), 
            .CO(n28404));
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4038));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13705_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13950), 
            .I3(GND_net), .O(n18212));   // verilog/coms.v(126[12] 289[6])
    defparam i13705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_add_1854_24_lut (.I0(GND_net), .I1(n2736_adj_4098), 
            .I2(VCC_net), .I3(n28187), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4216), .I3(n28402), .O(n18_adj_3993)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_31__I_0_add_1854_24 (.CI(n28187), .I0(n2736_adj_4098), 
            .I1(VCC_net), .CO(n28188));
    SB_LUT4 communication_counter_31__I_0_add_1854_23_lut (.I0(GND_net), .I1(n2737_adj_4097), 
            .I2(VCC_net), .I3(n28186), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1596_3_lut (.I0(n2347), .I1(n2414), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i17_3_lut (.I0(communication_counter[16]), 
            .I1(n17_adj_3968), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1958));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4037));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1335_3_lut (.I0(n1958), .I1(n2025), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_9 (.CI(n28402), .I0(GND_net), .I1(n18_adj_4216), 
            .CO(n28403));
    SB_CARRY communication_counter_31__I_0_add_1854_23 (.CI(n28186), .I0(n2737_adj_4097), 
            .I1(VCC_net), .CO(n28187));
    SB_LUT4 div_46_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4217), .I3(n28401), .O(n19_adj_3992)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_add_1854_22_lut (.I0(GND_net), .I1(n2738_adj_4096), 
            .I2(VCC_net), .I3(n28185), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_31__I_0_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_31__I_0_i1402_3_lut (.I0(n2057), .I1(n2124), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1469_3_lut (.I0(n2156), .I1(n2223), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1536_3_lut (.I0(n2255), .I1(n2322), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_8 (.CI(n28401), .I0(GND_net), .I1(n19_adj_4217), 
            .CO(n28402));
    SB_CARRY communication_counter_31__I_0_add_1854_22 (.CI(n28185), .I0(n2738_adj_4096), 
            .I1(VCC_net), .CO(n28186));
    SB_LUT4 communication_counter_31__I_0_i1603_3_lut (.I0(n2354), .I1(n2421), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2453_adj_4230));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4036));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13706_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13950), 
            .I3(GND_net), .O(n18213));   // verilog/coms.v(126[12] 289[6])
    defparam i13706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1600_3_lut (.I0(n2351), .I1(n2418), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2450_adj_4233));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1594_3_lut (.I0(n2345), .I1(n2412), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1594_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_LUT4 communication_counter_31__I_0_i1593_3_lut (.I0(n2344), .I1(n2411), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1602_3_lut (.I0(n2353), .I1(n2420), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2452_adj_4231));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1601_3_lut (.I0(n2352), .I1(n2419), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2451_adj_4232));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1598_3_lut (.I0(n2349), .I1(n2416), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2448_adj_4235));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1595_3_lut (.I0(n2346_adj_4240), 
            .I1(n2413), .I2(n2372_adj_4237), .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4035));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4034));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13707_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13950), 
            .I3(GND_net), .O(n18214));   // verilog/coms.v(126[12] 289[6])
    defparam i13707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4033));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1589_3_lut (.I0(n2340), .I1(n2407), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34170_3_lut (.I0(n40491), .I1(n86), .I2(n37_adj_4447), .I3(GND_net), 
            .O(n40492));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34170_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33335_4_lut (.I0(n41_adj_4450), .I1(n39_adj_4449), .I2(n37_adj_4447), 
            .I3(n39669), .O(n39657));
    defparam i33335_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4032));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1765_3_lut_3_lut (.I0(n2642), .I1(n6920), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_58[0]));   // verilog/TinyFPGA_B.v(120[10] 133[6])
    SB_LUT4 communication_counter_31__I_0_i1599_3_lut (.I0(n2350), .I1(n2417), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2449_adj_4234));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4031));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4030));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4029));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_mux_3_i16_3_lut (.I0(communication_counter[15]), 
            .I1(n18_adj_3967), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2058));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4028));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1403_3_lut (.I0(n2058), .I1(n2125), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1470_3_lut (.I0(n2157), .I1(n2224), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1537_3_lut (.I0(n2256), .I1(n2323), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4027));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4026));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13708_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13950), 
            .I3(GND_net), .O(n18215));   // verilog/coms.v(126[12] 289[6])
    defparam i13708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i14_3_lut (.I0(communication_counter[13]), 
            .I1(n20_adj_3965), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2258));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4025));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4024));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_3934));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1539_3_lut (.I0(n2258), .I1(n2325), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2357_adj_4239));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13709_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13950), 
            .I3(GND_net), .O(n18216));   // verilog/coms.v(126[12] 289[6])
    defparam i13709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i13_3_lut (.I0(communication_counter[12]), 
            .I1(n21_adj_3964), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2358_adj_4238));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i12_3_lut (.I0(communication_counter[11]), 
            .I1(n22_adj_3963), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2458_adj_4225));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_3984));   // verilog/TinyFPGA_B.v(208[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1607_3_lut (.I0(n2358_adj_4238), 
            .I1(n2425), .I2(n2372_adj_4237), .I3(GND_net), .O(n2457_adj_4226));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1606_3_lut (.I0(n2357_adj_4239), 
            .I1(n2424), .I2(n2372_adj_4237), .I3(GND_net), .O(n2456_adj_4227));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i15_3_lut (.I0(communication_counter[14]), 
            .I1(n19_adj_3966), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n2158));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1471_3_lut (.I0(n2158), .I1(n2225), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1257_3_lut (.I0(n1848), .I1(n1915), 
            .I2(n1877), .I3(GND_net), .O(n1947));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1330_3_lut (.I0(n1953), .I1(n2020), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1324_3_lut (.I0(n1947), .I1(n2014), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1391_3_lut (.I0(n2046), .I1(n2113), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13710_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13950), 
            .I3(GND_net), .O(n18217));   // verilog/coms.v(126[12] 289[6])
    defparam i13710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1458_3_lut (.I0(n2145), .I1(n2212), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1256_3_lut (.I0(n1847), .I1(n1914), 
            .I2(n1877), .I3(GND_net), .O(n1946));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1323_3_lut (.I0(n1946), .I1(n2013), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1390_3_lut (.I0(n2045), .I1(n2112), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1254_3_lut (.I0(n1845), .I1(n1912), 
            .I2(n1877), .I3(GND_net), .O(n1944));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1321_3_lut (.I0(n1944), .I1(n2011), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13711_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13950), 
            .I3(GND_net), .O(n18218));   // verilog/coms.v(126[12] 289[6])
    defparam i13711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1388_3_lut (.I0(n2043), .I1(n2110), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1455_3_lut (.I0(n2142), .I1(n2209), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13712_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13950), 
            .I3(GND_net), .O(n18219));   // verilog/coms.v(126[12] 289[6])
    defparam i13712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1255_3_lut (.I0(n1846), .I1(n1913), 
            .I2(n1877), .I3(GND_net), .O(n1945));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1322_3_lut (.I0(n1945), .I1(n2012), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1389_3_lut (.I0(n2044), .I1(n2111), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1456_3_lut (.I0(n2143), .I1(n2210), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1457_3_lut (.I0(n2144), .I1(n2211), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1766_3_lut_3_lut (.I0(n2642), .I1(n6921), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1524_3_lut (.I0(n2243), .I1(n2310), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13713_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13950), 
            .I3(GND_net), .O(n18220));   // verilog/coms.v(126[12] 289[6])
    defparam i13713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1523_3_lut (.I0(n2242), .I1(n2309), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1522_3_lut (.I0(n2241), .I1(n2308), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13714_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13950), 
            .I3(GND_net), .O(n18221));   // verilog/coms.v(126[12] 289[6])
    defparam i13714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i1263_3_lut (.I0(n1854), .I1(n1921), 
            .I2(n1877), .I3(GND_net), .O(n1953));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34230_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_4254), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1260_3_lut (.I0(n1851), .I1(n1918), 
            .I2(n1877), .I3(GND_net), .O(n1950));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13715_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13950), .I3(GND_net), .O(n18222));   // verilog/coms.v(126[12] 289[6])
    defparam i13715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13716_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13950), .I3(GND_net), .O(n18223));   // verilog/coms.v(126[12] 289[6])
    defparam i13716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13717_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13950), .I3(GND_net), .O(n18224));   // verilog/coms.v(126[12] 289[6])
    defparam i13717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1327_3_lut (.I0(n1950), .I1(n2017), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1394_3_lut (.I0(n2049), .I1(n2116), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1461_3_lut (.I0(n2148), .I1(n2215), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i1_3_lut (.I0(communication_counter[0]), 
            .I1(n33), .I2(communication_counter[31]), .I3(GND_net), .O(n3459));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i1464_3_lut (.I0(n2151), .I1(n2218), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1529_3_lut (.I0(n2248), .I1(n2315), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1534_3_lut (.I0(n2253), .I1(n2320), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i2_3_lut (.I0(communication_counter[1]), 
            .I1(n32_adj_3954), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n3458));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i1531_3_lut (.I0(n2250), .I1(n2317), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2287_3_lut (.I0(n3358), .I1(n10710), 
            .I2(n3362), .I3(GND_net), .O(n3457));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i2286_3_lut (.I0(n3357), .I1(n10709), 
            .I2(n3362), .I3(GND_net), .O(n3456));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i1528_3_lut (.I0(n2247), .I1(n2314), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2346_adj_4240));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n36865));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(n1854), .I1(n36865), .I2(n1855), .I3(n1857), 
            .O(n34678));
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'ha080;
    SB_LUT4 i7_4_lut (.I0(n1846), .I1(n1848), .I2(n1847), .I3(n34678), 
            .O(n18_adj_4614));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1853), .I1(n1851), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4615));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13718_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13950), .I3(GND_net), .O(n18225));   // verilog/coms.v(126[12] 289[6])
    defparam i13718_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    SB_LUT4 communication_counter_31__I_0_i2285_3_lut (.I0(n3356), .I1(n10708), 
            .I2(n3362), .I3(GND_net), .O(n3455));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 communication_counter_31__I_0_i2284_3_lut (.I0(n3355), .I1(n10707), 
            .I2(n3362), .I3(GND_net), .O(n3454));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2284_3_lut.LUT_INIT = 16'h3535;
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .n18368(n18368), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .n18367(n18367), .n18366(n18366), .n18365(n18365), .GND_net(GND_net), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_in_frame[19] ({\data_in_frame[19] }), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .rx_data({rx_data}), 
         .n18372(n18372), .n18371(n18371), .n18370(n18370), .n18369(n18369), 
         .n41916(n41916), .VCC_net(VCC_net), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .n18427(n18427), .control_mode({control_mode}), .n18428(n18428), 
         .PWMLimit({PWMLimit}), .n18429(n18429), .n18430(n18430), .n18431(n18431), 
         .n18432(n18432), .n18433(n18433), .n18421(n18421), .n18422(n18422), 
         .n18423(n18423), .n18424(n18424), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n18447(n18447), .n18448(n18448), .n18449(n18449), .n18450(n18450), 
         .n18445(n18445), .n18446(n18446), .n18443(n18443), .n18444(n18444), 
         .n18441(n18441), .n18442(n18442), .n18439(n18439), .n18440(n18440), 
         .n18437(n18437), .n18438(n18438), .n18434(n18434), .n18435(n18435), 
         .n18436(n18436), .n18425(n18425), .n18426(n18426), .n18245(n18245), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n18244(n18244), 
         .n18243(n18243), .n18242(n18242), .n18241(n18241), .n18240(n18240), 
         .n18239(n18239), .n18238(n18238), .n18237(n18237), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n18236(n18236), .n18235(n18235), .n18234(n18234), .n18233(n18233), 
         .n18232(n18232), .n18231(n18231), .n18230(n18230), .n18229(n18229), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .n18228(n18228), 
         .n18227(n18227), .n18226(n18226), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\byte_transmit_counter[1] (byte_transmit_counter[1]), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .n21(n21_adj_4564), 
         .n18225(n18225), .n18224(n18224), .n18223(n18223), .n18222(n18222), 
         .n18221(n18221), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n18220(n18220), .n35752(n35752), .n18219(n18219), .n18218(n18218), 
         .n18217(n18217), .n18216(n18216), .n18215(n18215), .n18214(n18214), 
         .n18213(n18213), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n18212(n18212), .n18211(n18211), .n18210(n18210), .n18209(n18209), 
         .n18208(n18208), .n18207(n18207), .n18206(n18206), .n18205(n18205), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .n18204(n18204), 
         .n18203(n18203), .n18202(n18202), .n18201(n18201), .n18200(n18200), 
         .n18199(n18199), .n18198(n18198), .n18197(n18197), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n18196(n18196), .n18195(n18195), .n18194(n18194), .rx_data_ready(rx_data_ready), 
         .n18193(n18193), .n18192(n18192), .n18191(n18191), .n18190(n18190), 
         .n18189(n18189), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n18188(n18188), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n36216(n36216), .n18187(n18187), .n18186(n18186), .n18185(n18185), 
         .n18184(n18184), .n18183(n18183), .n18182(n18182), .n18181(n18181), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .n18180(n18180), 
         .n18179(n18179), .n18178(n18178), .n18177(n18177), .n18176(n18176), 
         .n18175(n18175), .n18174(n18174), .n18173(n18173), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n18172(n18172), .n18171(n18171), .n18170(n18170), .n18169(n18169), 
         .n18168(n18168), .n18167(n18167), .n18166(n18166), .n18165(n18165), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .n18164(n18164), 
         .n18163(n18163), .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), 
         .\data_in[3] ({\data_in[3] }), .\data_in[2] ({\data_in[2] }), .n18162(n18162), 
         .n18161(n18161), .n18160(n18160), .n18159(n18159), .n18158(n18158), 
         .n18157(n18157), .\data_out_frame[9] ({\data_out_frame[9] }), .n18156(n18156), 
         .n18155(n18155), .n18154(n18154), .n18153(n18153), .n18152(n18152), 
         .n18151(n18151), .n18150(n18150), .n18149(n18149), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .n3761(n3761), .n16420(n16420), .n18148(n18148), .n18147(n18147), 
         .n18146(n18146), .n18145(n18145), .n18144(n18144), .n18143(n18143), 
         .n18142(n18142), .n25598(n25598), .n18141(n18141), .n18140(n18140), 
         .n18139(n18139), .n18138(n18138), .n18137(n18137), .n18136(n18136), 
         .n18135(n18135), .n18134(n18134), .n18133(n18133), .n18132(n18132), 
         .n18131(n18131), .n35990(n35990), .n18130(n18130), .n18129(n18129), 
         .n18128(n18128), .n18127(n18127), .n18126(n18126), .n18125(n18125), 
         .n18124(n18124), .n18123(n18123), .n18122(n18122), .n18121(n18121), 
         .n18120(n18120), .n18119(n18119), .n18118(n18118), .n63(n63_adj_4076), 
         .n123(n123), .n16404(n16404), .n2857(n2857), .n5(n5_adj_4077), 
         .n18114(n18114), .\Kp[7] (Kp[7]), .n18113(n18113), .\Kp[6] (Kp[6]), 
         .n42588(n42588), .n18112(n18112), .\Kp[5] (Kp[5]), .n18111(n18111), 
         .\Kp[4] (Kp[4]), .n18110(n18110), .\Kp[3] (Kp[3]), .n18109(n18109), 
         .\Kp[2] (Kp[2]), .n18108(n18108), .\Kp[1] (Kp[1]), .n18107(n18107), 
         .n16405(n16405), .n37137(n37137), .n18106(n18106), .n18105(n18105), 
         .n9783(n9783), .n18104(n18104), .n18103(n18103), .n18102(n18102), 
         .n18101(n18101), .n18100(n18100), .n18099(n18099), .n18098(n18098), 
         .n18097(n18097), .n18096(n18096), .n18095(n18095), .n18094(n18094), 
         .n18093(n18093), .n18092(n18092), .n18091(n18091), .n18090(n18090), 
         .n18089(n18089), .n18088(n18088), .n18087(n18087), .n18086(n18086), 
         .n18085(n18085), .n18084(n18084), .n18083(n18083), .n18082(n18082), 
         .n18081(n18081), .n18080(n18080), .n18079(n18079), .n18078(n18078), 
         .n18077(n18077), .n18075(n18075), .gearBoxRatio({gearBoxRatio}), 
         .n18074(n18074), .n18073(n18073), .n18072(n18072), .n18071(n18071), 
         .n18070(n18070), .n18069(n18069), .n18068(n18068), .n18067(n18067), 
         .n18066(n18066), .n18065(n18065), .n18064(n18064), .n18063(n18063), 
         .n18062(n18062), .n18061(n18061), .n18060(n18060), .n18059(n18059), 
         .n18058(n18058), .n18057(n18057), .n18056(n18056), .n18055(n18055), 
         .n18054(n18054), .n18053(n18053), .n17974(n17974), .setpoint({setpoint}), 
         .n17973(n17973), .n17972(n17972), .n17971(n17971), .n17970(n17970), 
         .n17969(n17969), .n17968(n17968), .n17967(n17967), .n17966(n17966), 
         .n17965(n17965), .n17964(n17964), .n17963(n17963), .n17962(n17962), 
         .n17961(n17961), .n17960(n17960), .n17959(n17959), .n17958(n17958), 
         .n17957(n17957), .n17956(n17956), .n17955(n17955), .n17954(n17954), 
         .n17953(n17953), .n17952(n17952), .LED_c(LED_c), .n18308(n18308), 
         .n18307(n18307), .\data_out_frame[21] ({Open_0, Open_1, Open_2, 
         Open_3, Open_4, Open_5, Open_6, \data_out_frame[21] [0]}), 
         .n35420(n35420), .\data_out_frame[22] ({Open_7, Open_8, Open_9, 
         Open_10, Open_11, Open_12, Open_13, \data_out_frame[22] [0]}), 
         .n34307(n34307), .n18306(n18306), .n18305(n18305), .n18304(n18304), 
         .n18303(n18303), .\r_SM_Main_2__N_3298[0] (r_SM_Main_2__N_3298[0]), 
         .n18302(n18302), .tx_active(tx_active), .n18301(n18301), .n33144(n33144), 
         .n17896(n17896), .n17895(n17895), .n17893(n17893), .\Kp[0] (Kp[0]), 
         .n17793(n17793), .n17791(n17791), .n17892(n17892), .n11748(n11748), 
         .n34073(n34073), .n19(n19_adj_4616), .n33787(n33787), .n33923(n33923), 
         .n33775(n33775), .n33766(n33766), .n16417(n16417), .n30686(n30686), 
         .n4423(n4423), .n4446(n4446), .n13950(n13950), .n4445(n4445), 
         .n4444(n4444), .n4443(n4443), .n4442(n4442), .n4441(n4441), 
         .n4440(n4440), .n4439(n4439), .n37188(n37188), .n4438(n4438), 
         .n4437(n4437), .n4436(n4436), .n4435(n4435), .n4434(n4434), 
         .n4433(n4433), .n16809(n16809), .n4432(n4432), .n4431(n4431), 
         .n4430(n4430), .n4429(n4429), .n4428(n4428), .n4427(n4427), 
         .n4426(n4426), .n4425(n4425), .n4424(n4424), .n18509(n18509), 
         .r_SM_Main({r_SM_Main_adj_4662}), .n17827(n17827), .r_Bit_Index({r_Bit_Index_adj_4664}), 
         .n17830(n17830), .\r_SM_Main_2__N_3295[1] (r_SM_Main_2__N_3295[1]), 
         .n17625(n17625), .n17748(n17748), .n4706(n4706), .n17989(n17989), 
         .tx_o(tx_o), .tx_enable(tx_enable), .n18539(n18539), .\r_Clock_Count[0] (r_Clock_Count[0]), 
         .n17836(n17836), .r_Bit_Index_adj_10({r_Bit_Index}), .n17833(n17833), 
         .\r_SM_Main[1]_adj_6 (r_SM_Main[1]), .\r_SM_Main[2]_adj_7 (r_SM_Main[2]), 
         .n2346(n2346), .r_Rx_Data(r_Rx_Data), .PIN_13_N_106(PIN_13_N_106), 
         .\r_Clock_Count[2] (r_Clock_Count[2]), .\r_Clock_Count[1] (r_Clock_Count[1]), 
         .\r_Clock_Count[6] (r_Clock_Count[6]), .\r_Clock_Count[4] (r_Clock_Count[4]), 
         .n16429(n16429), .n4(n4_adj_4023), .n35922(n35922), .n4684(n4684), 
         .n17619(n17619), .n17746(n17746), .n17931(n17931), .n17936(n17936), 
         .n17942(n17942), .n17980(n17980), .n17992(n17992), .n18003(n18003), 
         .n33396(n33396), .n220(n220), .n222(n222), .n224(n224_adj_4014), 
         .n225(n225), .n226(n226), .n24632(n24632), .n4_adj_8(n4), .n4_adj_9(n4_adj_4022), 
         .n16424(n16424), .n17843(n17843), .n17842(n17842), .n17841(n17841), 
         .n17840(n17840), .n17839(n17839), .n17838(n17838), .n17837(n17837), 
         .n17522(n17522)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(161[8] 181[4])
    SB_LUT4 i13385_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17892));   // verilog/coms.v(126[12] 289[6])
    defparam i13385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13284_3_lut (.I0(setpoint[0]), .I1(n4423), .I2(n36216), .I3(GND_net), 
            .O(n17791));   // verilog/coms.v(126[12] 289[6])
    defparam i13284_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13285_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n37153), .I3(GND_net), .O(n17792));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13285_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2283_3_lut (.I0(n3354), .I1(n10706), 
            .I2(n3362), .I3(GND_net), .O(n3453));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i9_4_lut (.I0(n1852), .I1(n18_adj_4614), .I2(n1845), .I3(n1844), 
            .O(n20_adj_4613));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13286_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[19] [0]), 
            .I2(n35752), .I3(GND_net), .O(n17793));   // verilog/coms.v(126[12] 289[6])
    defparam i13286_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34675_2_lut (.I0(n3362), .I1(n10705), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34675_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i10_4_lut (.I0(n1849), .I1(n20_adj_4613), .I2(n16_adj_4615), 
            .I3(n1850), .O(n1877));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i18_3_lut (.I0(communication_counter[17]), 
            .I1(n16_adj_3969), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1858));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35398_1_lut (.I0(n1778_adj_4345), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n41718));
    defparam i35398_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1767_3_lut_3_lut (.I0(n2642), .I1(n6922), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1589 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n34667));
    defparam i1_3_lut_adj_1589.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1590 (.I0(n1947), .I1(n1954), .I2(n34667), .I3(n1955), 
            .O(n15_adj_4602));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i3_4_lut_adj_1590.LUT_INIT = 16'heaaa;
    SB_LUT4 i34478_4_lut (.I0(n38_adj_4448), .I1(n18_adj_4435), .I2(n43_adj_4451), 
            .I3(n39653), .O(n40800));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34478_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i7_4_lut_adj_1591 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4600));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i7_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1953), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4601));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1592 (.I0(n19_adj_4600), .I1(n15_adj_4602), .I2(n1948), 
            .I3(n1952), .O(n22_adj_4599));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i10_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1773_3_lut_3_lut (.I0(n2642), .I1(n6928), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11_4_lut_adj_1593 (.I0(n1950), .I1(n22_adj_4599), .I2(n18_adj_4601), 
            .I3(n1949), .O(n1976_adj_4266));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1267_3_lut (.I0(n1858), .I1(n1925), 
            .I2(n1877), .I3(GND_net), .O(n1957));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1594 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n34710));
    defparam i1_3_lut_adj_1594.LUT_INIT = 16'hfefe;
    SB_LUT4 communication_counter_31__I_0_i1121_3_lut (.I0(n1648_adj_4123), 
            .I1(n1715), .I2(n1679), .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34235_3_lut (.I0(n1553_adj_4130), .I1(n1620), .I2(n1580), 
            .I3(GND_net), .O(n1652_adj_4127));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34236_3_lut (.I0(n1652_adj_4127), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1595 (.I0(n2054), .I1(n2048), .I2(n34710), .I3(n2055), 
            .O(n17_adj_4558));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i4_4_lut_adj_1595.LUT_INIT = 16'heccc;
    SB_LUT4 communication_counter_31__I_0_i1129_3_lut (.I0(n1656), .I1(n1723), 
            .I2(n1679), .I3(GND_net), .O(n1755_adj_4366));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut (.I0(n2044), .I1(n2046), .I2(n2045), .I3(n2047), 
            .O(n21_adj_4556));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1127_3_lut (.I0(n1654), .I1(n1721), 
            .I2(n1679), .I3(GND_net), .O(n1753));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1128_3_lut (.I0(n1655), .I1(n1722), 
            .I2(n1679), .I3(GND_net), .O(n1754_adj_4367));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut (.I0(n2051), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_4557));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1596 (.I0(n21_adj_4556), .I1(n17_adj_4558), .I2(n2053), 
            .I3(n2050), .O(n24_adj_4555));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1597 (.I0(n2049), .I1(n24_adj_4555), .I2(n20_adj_4557), 
            .I3(n2052), .O(n2075_adj_4254));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1334_3_lut (.I0(n1957), .I1(n2024), 
            .I2(n1976_adj_4266), .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_4_lut (.I0(n131), .I1(n39062), .I2(state[0]), .I3(n21_adj_3947), 
            .O(n19_adj_4546));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 communication_counter_31__I_0_i1131_rep_52_3_lut (.I0(n1658), 
            .I1(n1725), .I2(n1679), .I3(GND_net), .O(n1757_adj_4347));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1131_rep_52_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1774_3_lut_3_lut (.I0(n2642), .I1(n6929), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1598 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n34672));
    defparam i1_3_lut_adj_1598.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1599 (.I0(n2154), .I1(n2147), .I2(n34672), .I3(n2155), 
            .O(n18_adj_4074));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i4_4_lut_adj_1599.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut_adj_1600 (.I0(n2150), .I1(n2152), .I2(n2148), .I3(n2153), 
            .O(n24_adj_4072));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i10_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1601 (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_4073));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i8_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1602 (.I0(n2145), .I1(n24_adj_4072), .I2(n18_adj_4074), 
            .I3(n2146), .O(n26_adj_4064));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1603 (.I0(n2151), .I1(n26_adj_4064), .I2(n22_adj_4073), 
            .I3(n2149), .O(n2174_adj_4245));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i13_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1130_3_lut (.I0(n1657), .I1(n1724), 
            .I2(n1679), .I3(GND_net), .O(n1756_adj_4348));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1120_3_lut (.I0(n1647_adj_4122), 
            .I1(n1714), .I2(n1679), .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1126_3_lut (.I0(n1653_adj_4128), 
            .I1(n1720), .I2(n1679), .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1123_3_lut (.I0(n1650_adj_4125), 
            .I1(n1717), .I2(n1679), .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1401_3_lut (.I0(n2056), .I1(n2123), 
            .I2(n2075_adj_4254), .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1122_3_lut (.I0(n1649_adj_4124), 
            .I1(n1716), .I2(n1679), .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1124_3_lut (.I0(n1651_adj_4126), 
            .I1(n1718), .I2(n1679), .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1604 (.I0(n1745), .I1(n1750), .I2(n1748), .I3(n1749), 
            .O(n16_adj_4618));
    defparam i6_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1605 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n34743));
    defparam i1_3_lut_adj_1605.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1606 (.I0(n1756_adj_4348), .I1(n1757_adj_4347), 
            .I2(n1758_adj_4346), .I3(GND_net), .O(n34651));
    defparam i1_3_lut_adj_1606.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1752), .I1(n16_adj_4618), .I2(n1746), .I3(GND_net), 
            .O(n18_adj_4617));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1607 (.I0(n2248), .I1(n2253), .I2(n2251), .I3(n2249), 
            .O(n26_adj_4052));
    defparam i11_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1608 (.I0(n1754_adj_4367), .I1(n1753), .I2(n34651), 
            .I3(n1755_adj_4366), .O(n13_adj_4619));
    defparam i3_4_lut_adj_1608.LUT_INIT = 16'heccc;
    SB_LUT4 i9_4_lut_adj_1609 (.I0(n13_adj_4619), .I1(n18_adj_4617), .I2(n1751), 
            .I3(n1747), .O(n1778_adj_4345));
    defparam i9_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1610 (.I0(n2246), .I1(n2254), .I2(n34743), .I3(n2255), 
            .O(n19_adj_4054));
    defparam i4_4_lut_adj_1610.LUT_INIT = 16'heaaa;
    SB_LUT4 communication_counter_31__I_0_mux_3_i19_3_lut (.I0(communication_counter[18]), 
            .I1(n15_adj_3970), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1758_adj_4346));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1611 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4056));
    defparam i1_2_lut_adj_1611.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1612 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_4053));
    defparam i9_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i13386_3_lut (.I0(Kp[0]), .I1(\data_in_frame[2] [0]), .I2(n35752), 
            .I3(GND_net), .O(n17893));   // verilog/coms.v(126[12] 289[6])
    defparam i13386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1657_3_lut (.I0(n2462), .I1(n6879), .I2(n2471), .I3(GND_net), 
            .O(n2549));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_1613 (.I0(n19_adj_4054), .I1(n26_adj_4052), .I2(n2247), 
            .I3(n2250), .O(n28_adj_4051));
    defparam i13_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i13388_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n35752), .I3(GND_net), .O(n17895));   // verilog/coms.v(126[12] 289[6])
    defparam i13388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut_adj_1614 (.I0(n2252), .I1(n28_adj_4051), .I2(n24_adj_4053), 
            .I3(n16_adj_4056), .O(n2273_adj_4242));
    defparam i14_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1468_3_lut (.I0(n2155), .I1(n2222), 
            .I2(n2174_adj_4245), .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34222_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4242), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1530_3_lut (.I0(n2249), .I1(n2316), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34368_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_4254), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1770_3_lut_3_lut (.I0(n2642), .I1(n6925), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[17] [5]), .I1(n33923), .I2(n34073), 
            .I3(GND_net), .O(n6_adj_4567));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n16520), 
            .O(n16472));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i34224_3_lut (.I0(n2251), .I1(n2318), .I2(n2273_adj_4242), 
            .I3(GND_net), .O(n2350));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1535_3_lut (.I0(n2254), .I1(n2321), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1802_3_lut (.I0(n2649), .I1(n2716_adj_4106), 
            .I2(n2669), .I3(GND_net), .O(n2748_adj_4086));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1526_3_lut (.I0(n2245), .I1(n2312), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1527_3_lut (.I0(n2246), .I1(n2313), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1525_3_lut (.I0(n2244), .I1(n2311), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1615 (.I0(n2356), .I1(n2358_adj_4238), .I2(GND_net), 
            .I3(GND_net), .O(n36797));
    defparam i1_2_lut_adj_1615.LUT_INIT = 16'heeee;
    SB_LUT4 i13719_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13950), .I3(GND_net), .O(n18226));   // verilog/coms.v(126[12] 289[6])
    defparam i13719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n2354), .I1(n36797), .I2(n2355), .I3(n2357_adj_4239), 
            .O(n34680));
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'ha080;
    SB_LUT4 i12_4_lut_adj_1617 (.I0(n2353), .I1(n2350), .I2(n2348), .I3(n2351), 
            .O(n28_adj_4119));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1618 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n34680), 
            .O(n26_adj_4133));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i10_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1619 (.I0(n2346_adj_4240), .I1(n2349), .I2(n2352), 
            .I3(n2347), .O(n27_adj_4132));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1620 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_4135));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i9_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1621 (.I0(n25_adj_4135), .I1(n27_adj_4132), .I2(n26_adj_4133), 
            .I3(n28_adj_4119), .O(n2372_adj_4237));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1771_3_lut_3_lut (.I0(n2642), .I1(n6926), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1538_3_lut (.I0(n2257), .I1(n2324), 
            .I2(n2273_adj_4242), .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1605_3_lut (.I0(n2356), .I1(n2423), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2455_adj_4228));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1604_3_lut (.I0(n2355), .I1(n2422), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2454_adj_4229));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1772_3_lut_3_lut (.I0(n2642), .I1(n6927), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1590_3_lut (.I0(n2341), .I1(n2408), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1622 (.I0(n2456_adj_4227), .I1(n2457_adj_4226), 
            .I2(n2458_adj_4225), .I3(GND_net), .O(n34749));
    defparam i1_3_lut_adj_1622.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_3_lut (.I0(n2449_adj_4234), .I1(n2439), .I2(n2438), .I3(GND_net), 
            .O(n26_adj_4606));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i9_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1623 (.I0(n2445), .I1(n2448_adj_4235), .I2(n2451_adj_4232), 
            .I3(n2452_adj_4231), .O(n29_adj_4604));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1624 (.I0(n2440), .I1(n2454_adj_4229), .I2(n34749), 
            .I3(n2455_adj_4228), .O(n20_adj_4607));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i3_4_lut_adj_1624.LUT_INIT = 16'heaaa;
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_78_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[0]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_107[0]), 
            .I2(n15), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_4598));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_1_lut (.I0(communication_counter[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4055));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1625 (.I0(n2443), .I1(n2444), .I2(n2450_adj_4233), 
            .I3(n2453_adj_4230), .O(n28_adj_4605));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i13720_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13950), .I3(GND_net), .O(n18227));   // verilog/coms.v(126[12] 289[6])
    defparam i13720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_4597));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_4596));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_4595));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13389_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[7] [0]), 
            .I2(n35752), .I3(GND_net), .O(n17896));   // verilog/coms.v(126[12] 289[6])
    defparam i13389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13390_3_lut (.I0(encoder0_position[0]), .I1(n2755), .I2(count_enable), 
            .I3(GND_net), .O(n17897));   // quad.v(35[10] 41[6])
    defparam i13390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13721_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13950), .I3(GND_net), .O(n18228));   // verilog/coms.v(126[12] 289[6])
    defparam i13721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n35990), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n36316), .I3(n11748), .O(n33144));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'hd5f5;
    SB_LUT4 i13722_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13950), .I3(GND_net), .O(n18229));   // verilog/coms.v(126[12] 289[6])
    defparam i13722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30933_3_lut_4_lut (.I0(n16404), .I1(n2857), .I2(n33787), 
            .I3(n37137), .O(n37188));
    defparam i30933_3_lut_4_lut.LUT_INIT = 16'he000;
    SB_LUT4 i13723_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13950), .I3(GND_net), .O(n18230));   // verilog/coms.v(126[12] 289[6])
    defparam i13723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_4594));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1627 (.I0(n82), .I1(n81), .I2(n80), 
            .I3(n16505), .O(n16547));
    defparam i1_2_lut_3_lut_4_lut_adj_1627.LUT_INIT = 16'hff7f;
    SB_LUT4 i15_4_lut_adj_1628 (.I0(n29_adj_4604), .I1(n2446), .I2(n26_adj_4606), 
            .I3(n2447_adj_4236), .O(n32_adj_4603));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i22752_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4_adj_3936));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22752_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i2_2_lut (.I0(n2442), .I1(n2441), .I2(GND_net), .I3(GND_net), 
            .O(n19_adj_4608));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut_adj_1629 (.I0(n19_adj_4608), .I1(n32_adj_4603), .I2(n28_adj_4605), 
            .I3(n20_adj_4607), .O(n2471_adj_4224));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i16_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i13794_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n33766), 
            .I3(GND_net), .O(n18301));   // verilog/coms.v(126[12] 289[6])
    defparam i13794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i1591_3_lut (.I0(n2342), .I1(n2409), 
            .I2(n2372_adj_4237), .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1658_3_lut (.I0(n2441), .I1(n2508), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2540_adj_4172));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1630 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n16505));
    defparam i1_2_lut_3_lut_adj_1630.LUT_INIT = 16'hf7f7;
    SB_LUT4 communication_counter_31__I_0_i1657_3_lut (.I0(n2440), .I1(n2507), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2539_adj_4173));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1656_3_lut (.I0(n2439), .I1(n2506), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2538_adj_4174));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4431));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10_4_lut_adj_1631 (.I0(n2538_adj_4174), .I1(n2539_adj_4173), 
            .I2(n2537_adj_4175), .I3(n2540_adj_4172), .O(n28_adj_4563));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i10_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i33369_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n39691));
    defparam i33369_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i1_2_lut_adj_1632 (.I0(n2556), .I1(n2558_adj_4158), .I2(GND_net), 
            .I3(GND_net), .O(n36817));
    defparam i1_2_lut_adj_1632.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4433));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_adj_1633 (.I0(n2554), .I1(n36817), .I2(n2555), .I3(n2557), 
            .O(n34684));
    defparam i1_4_lut_adj_1633.LUT_INIT = 16'ha080;
    SB_LUT4 i14_3_lut (.I0(n2547_adj_4165), .I1(n28_adj_4563), .I2(n2549_adj_4163), 
            .I3(GND_net), .O(n32_adj_4559));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i22728_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_4610));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22728_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 communication_counter_31__I_0_i1061_3_lut (.I0(n1556), .I1(n1623), 
            .I2(n1580), .I3(GND_net), .O(n1655));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1060_3_lut (.I0(n1555), .I1(n1622), 
            .I2(n1580), .I3(GND_net), .O(n1654));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1054_3_lut (.I0(n1549), .I1(n1616), 
            .I2(n1580), .I3(GND_net), .O(n1648_adj_4123));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1634 (.I0(n34684), .I1(n2546_adj_4166), .I2(n2545_adj_4167), 
            .I3(n2553_adj_4159), .O(n30_adj_4561));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1635 (.I0(n2548_adj_4164), .I1(n2551_adj_4161), 
            .I2(n2552_adj_4160), .I3(n2550_adj_4162), .O(n31_adj_4560));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i13_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1636 (.I0(n2541_adj_4171), .I1(n2543_adj_4169), 
            .I2(n2542_adj_4170), .I3(n2544_adj_4168), .O(n29_adj_4562));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1637 (.I0(n29_adj_4562), .I1(n31_adj_4560), .I2(n30_adj_4561), 
            .I3(n32_adj_4559), .O(n2570));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1056_3_lut (.I0(n1551), .I1(n1618), 
            .I2(n1580), .I3(GND_net), .O(n1650_adj_4125));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1660_3_lut (.I0(n2443), .I1(n2510), 
            .I2(n2471_adj_4224), .I3(GND_net), .O(n2542_adj_4170));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1727_3_lut (.I0(n2542_adj_4170), 
            .I1(n2609), .I2(n2570), .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1725_3_lut (.I0(n2540_adj_4172), 
            .I1(n2607), .I2(n2570), .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13724_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13950), .I3(GND_net), .O(n18231));   // verilog/coms.v(126[12] 289[6])
    defparam i13724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1724_3_lut (.I0(n2539_adj_4173), 
            .I1(n2606), .I2(n2570), .I3(GND_net), .O(n2638_adj_4136));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1638 (.I0(n2638_adj_4136), .I1(n2640), .I2(n2639), 
            .I3(n2641), .O(n30_adj_4061));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i11_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1639 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n37033));
    defparam i1_2_lut_adj_1639.LUT_INIT = 16'heeee;
    SB_LUT4 communication_counter_31__I_0_i1055_3_lut (.I0(n1550), .I1(n1617), 
            .I2(n1580), .I3(GND_net), .O(n1649_adj_4124));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n2654), .I1(n37033), .I2(n2655), .I3(n2657), 
            .O(n34761));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'ha080;
    SB_LUT4 i15_4_lut_adj_1641 (.I0(n2650), .I1(n30_adj_4061), .I2(n2637_adj_4137), 
            .I3(n2636_adj_4138), .O(n34_adj_4057));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i15_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i1057_3_lut (.I0(n1552), .I1(n1619), 
            .I2(n1580), .I3(GND_net), .O(n1651_adj_4126));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1642 (.I0(n2645), .I1(n2651), .I2(n2646), .I3(n2649), 
            .O(n32_adj_4059));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i13_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i13725_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13950), .I3(GND_net), .O(n18232));   // verilog/coms.v(126[12] 289[6])
    defparam i13725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1059_rep_53_3_lut (.I0(n1554_adj_4131), 
            .I1(n1621), .I2(n1580), .I3(GND_net), .O(n1653_adj_4128));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1059_rep_53_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut_adj_1643 (.I0(n2652), .I1(n2648), .I2(n2653), .I3(n2647), 
            .O(n33_adj_4058));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1644 (.I0(n2642_adj_4134), .I1(n34761), .I2(n2643_adj_4120), 
            .I3(n2644), .O(n31_adj_4060));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i12_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1645 (.I0(n31_adj_4060), .I1(n33_adj_4058), .I2(n32_adj_4059), 
            .I3(n34_adj_4057), .O(n2669));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i18_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1768_3_lut_3_lut (.I0(n2642), .I1(n6923), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_31__I_0_i1726_3_lut (.I0(n2541_adj_4171), 
            .I1(n2608), .I2(n2570), .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1063_3_lut (.I0(n1558), .I1(n1625), 
            .I2(n1580), .I3(GND_net), .O(n1657));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1062_rep_54_3_lut (.I0(n1557), 
            .I1(n1624), .I2(n1580), .I3(GND_net), .O(n1656));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1062_rep_54_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1793_3_lut (.I0(n2640), .I1(n2707_adj_4115), 
            .I2(n2669), .I3(GND_net), .O(n2739_adj_4095));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1053_3_lut (.I0(n1548), .I1(n1615), 
            .I2(n1580), .I3(GND_net), .O(n1647_adj_4122));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_3_lut_4_lut (.I0(n16420), .I1(n3761), .I2(n37188), .I3(n19_adj_4616), 
            .O(n36316));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'hff1f;
    SB_LUT4 i1_2_lut_adj_1646 (.I0(n1647_adj_4122), .I1(n1646_adj_4121), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3946));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i1_2_lut_adj_1646.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1647 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n34659));
    defparam i1_3_lut_adj_1647.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1648 (.I0(n1653_adj_4128), .I1(n1652_adj_4127), 
            .I2(n1651_adj_4126), .I3(n10_adj_3946), .O(n16_adj_3944));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i7_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1649 (.I0(n1648_adj_4123), .I1(n1654), .I2(n34659), 
            .I3(n1655), .O(n11_adj_3945));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i2_4_lut_adj_1649.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut_adj_1650 (.I0(n11_adj_3945), .I1(n16_adj_3944), .I2(n1649_adj_4124), 
            .I3(n1650_adj_4125), .O(n1679));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i8_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i20_3_lut (.I0(communication_counter[19]), 
            .I1(n14_adj_3971), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1658));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_4593));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_4592));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1763_3_lut_3_lut (.I0(n2642), .I1(n6918), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_3996), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13726_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13950), .I3(GND_net), .O(n18233));   // verilog/coms.v(126[12] 289[6])
    defparam i13726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1271_3_lut (.I0(n381), .I1(n6766), .I2(n1886), .I3(GND_net), 
            .O(n1980));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13727_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13950), .I3(GND_net), .O(n18234));   // verilog/coms.v(126[12] 289[6])
    defparam i13727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1340_3_lut (.I0(n1980), .I1(n6782), .I2(n1991), .I3(GND_net), 
            .O(n2082));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1407_3_lut (.I0(n2082), .I1(n6799), .I2(n2093), .I3(GND_net), 
            .O(n2181));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1472_3_lut (.I0(n2181), .I1(n6817), .I2(n2192), .I3(GND_net), 
            .O(n2277));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1472_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13728_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13950), .I3(GND_net), .O(n18235));   // verilog/coms.v(126[12] 289[6])
    defparam i13728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1535_3_lut (.I0(n2277), .I1(n6836), .I2(n2288), .I3(GND_net), 
            .O(n2370));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1535_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13729_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13950), .I3(GND_net), .O(n18236));   // verilog/coms.v(126[12] 289[6])
    defparam i13729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i367_4_lut (.I0(n34342), .I1(n4_adj_4610), .I2(n533), 
            .I3(n98), .O(n34344));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i367_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i13730_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13950), .I3(GND_net), .O(n18237));   // verilog/coms.v(126[12] 289[6])
    defparam i13730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22760_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_3936), .I3(GND_net), 
            .O(n6_adj_3935));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22760_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_i458_4_lut (.I0(n34344), .I1(n6_adj_3935), .I2(n671), 
            .I3(n97), .O(n34346));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i458_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i18900_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13950), .I3(GND_net), .O(n18238));
    defparam i18900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22800_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4611), .I3(GND_net), 
            .O(n8_adj_4609));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22800_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_i547_4_lut (.I0(n34346), .I1(n8_adj_4609), .I2(n806), 
            .I3(n96), .O(n914));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i547_4_lut.LUT_INIT = 16'h5659;
    SB_LUT4 i13732_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13950), .I3(GND_net), .O(n18239));   // verilog/coms.v(126[12] 289[6])
    defparam i13732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i634_3_lut (.I0(n914), .I1(n6661), .I2(n938), .I3(GND_net), 
            .O(n1043));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13733_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13950), .I3(GND_net), .O(n18240));   // verilog/coms.v(126[12] 289[6])
    defparam i13733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13734_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13950), .I3(GND_net), .O(n18241));   // verilog/coms.v(126[12] 289[6])
    defparam i13734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13735_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13950), .I3(GND_net), .O(n18242));   // verilog/coms.v(126[12] 289[6])
    defparam i13735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33653_3_lut (.I0(n40492), .I1(n85), .I2(n39_adj_4449), .I3(GND_net), 
            .O(n39975));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33653_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i719_3_lut (.I0(n1043), .I1(n6669), .I2(n1067), .I3(GND_net), 
            .O(n1169));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i802_3_lut (.I0(n1169), .I1(n6678), .I2(n1193), .I3(GND_net), 
            .O(n1292));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i883_3_lut (.I0(n1292), .I1(n6688), .I2(n1316), .I3(GND_net), 
            .O(n1412));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i24_3_lut (.I0(n16_adj_4433), .I1(n91), 
            .I2(n27_adj_4442), .I3(GND_net), .O(n24_adj_4440));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34508_4_lut (.I0(n24_adj_4440), .I1(n14_adj_4431), .I2(n27_adj_4442), 
            .I3(n39691), .O(n40830));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34508_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34509_3_lut (.I0(n40830), .I1(n90), .I2(n29_adj_4443), .I3(GND_net), 
            .O(n40831));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34509_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34395_3_lut (.I0(n40831), .I1(n89), .I2(n31_adj_4444), .I3(GND_net), 
            .O(n40717));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34395_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34320_4_lut (.I0(n41_adj_4450), .I1(n39_adj_4449), .I2(n37_adj_4447), 
            .I3(n39673), .O(n40642));
    defparam i34320_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34605_4_lut (.I0(n39975), .I1(n40800), .I2(n43_adj_4451), 
            .I3(n39657), .O(n40927));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34605_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33651_3_lut (.I0(n40717), .I1(n88), .I2(n33_adj_4445), .I3(GND_net), 
            .O(n39973));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33651_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i962_3_lut (.I0(n1412), .I1(n6699), .I2(n1436), .I3(GND_net), 
            .O(n1529));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1039_3_lut (.I0(n1529), .I1(n6711), .I2(n1553), .I3(GND_net), 
            .O(n1643));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1114_3_lut (.I0(n1643), .I1(n6724), .I2(n1667), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13736_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13950), .I3(GND_net), .O(n18243));   // verilog/coms.v(126[12] 289[6])
    defparam i13736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1187_3_lut (.I0(n1754), .I1(n6738), .I2(n1778), .I3(GND_net), 
            .O(n1862));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1258_3_lut (.I0(n1862), .I1(n6753), .I2(n1886), .I3(GND_net), 
            .O(n1967));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1327_3_lut (.I0(n1967), .I1(n6769), .I2(n1991), .I3(GND_net), 
            .O(n2069));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13737_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13950), .I3(GND_net), .O(n18244));   // verilog/coms.v(126[12] 289[6])
    defparam i13737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1394_3_lut (.I0(n2069), .I1(n6786), .I2(n2093), .I3(GND_net), 
            .O(n2168));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4435));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33331_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n39653));
    defparam i33331_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1459_3_lut (.I0(n2168), .I1(n6804), .I2(n2192), .I3(GND_net), 
            .O(n2264));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1459_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4000), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1651 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n16508));
    defparam i1_2_lut_adj_1651.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4437));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i1522_3_lut (.I0(n2264), .I1(n6823), .I2(n2288), .I3(GND_net), 
            .O(n2357));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1583_3_lut (.I0(n2357), .I1(n6843), .I2(n2381), .I3(GND_net), 
            .O(n2447));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1652 (.I0(n80), .I1(n16505), .I2(GND_net), .I3(GND_net), 
            .O(n16502));
    defparam i1_2_lut_adj_1652.LUT_INIT = 16'hdddd;
    SB_LUT4 i22720_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3983));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22720_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13795_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n33766), 
            .I3(GND_net), .O(n18302));   // verilog/coms.v(126[12] 289[6])
    defparam i13795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13796_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n33766), 
            .I3(GND_net), .O(n18303));   // verilog/coms.v(126[12] 289[6])
    defparam i13796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i368_4_lut (.I0(n510), .I1(n2_adj_3983), .I2(n533), 
            .I3(n99), .O(n648));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i368_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4591));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1653 (.I0(n81), .I1(n80), .I2(n16505), 
            .I3(GND_net), .O(n16498));
    defparam i1_2_lut_3_lut_adj_1653.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13797_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n33766), 
            .I3(GND_net), .O(n18304));   // verilog/coms.v(126[12] 289[6])
    defparam i13797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22792_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4612), .I3(GND_net), 
            .O(n6_adj_4611));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22792_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_i459_4_lut (.I0(n648), .I1(n4_adj_3936), .I2(n671), 
            .I3(n98), .O(n783));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i459_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i13798_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n33766), 
            .I3(GND_net), .O(n18305));   // verilog/coms.v(126[12] 289[6])
    defparam i13798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34646_4_lut (.I0(n39973), .I1(n40927), .I2(n43_adj_4451), 
            .I3(n40642), .O(n40968));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34646_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i548_4_lut (.I0(n783), .I1(n6_adj_4611), .I2(n806), 
            .I3(n97), .O(n915));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i548_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_46_i635_3_lut (.I0(n915), .I1(n6662), .I2(n938), .I3(GND_net), 
            .O(n1044));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i720_3_lut (.I0(n1044), .I1(n6670), .I2(n1067), .I3(GND_net), 
            .O(n1170));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i803_3_lut (.I0(n1170), .I1(n6679), .I2(n1193), .I3(GND_net), 
            .O(n1293));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34647_3_lut (.I0(n40968), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n40969));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i34647_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i884_3_lut (.I0(n1293), .I1(n6689), .I2(n1316), .I3(GND_net), 
            .O(n1413));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13392_3_lut (.I0(encoder1_position[0]), .I1(n2705), .I2(count_enable_adj_4011), 
            .I3(GND_net), .O(n17899));   // quad.v(35[10] 41[6])
    defparam i13392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4590));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i971_3_lut (.I0(n377), .I1(n6708), .I2(n1436), .I3(GND_net), 
            .O(n1538));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4589));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4588));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1654 (.I0(n83), .I1(n82), .I2(n16498), 
            .I3(GND_net), .O(n16495));
    defparam i1_2_lut_3_lut_adj_1654.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(n84), .I1(n83), .I2(n16547), 
            .I3(GND_net), .O(n16491));
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1656 (.I0(n85), .I1(n84), .I2(n16495), 
            .I3(GND_net), .O(n16544));
    defparam i1_2_lut_3_lut_adj_1656.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1657 (.I0(n86), .I1(n85), .I2(n16491), 
            .I3(GND_net), .O(n16485));
    defparam i1_2_lut_3_lut_adj_1657.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1658 (.I0(n87), .I1(n86), .I2(n16544), 
            .I3(GND_net), .O(n16541));
    defparam i1_2_lut_3_lut_adj_1658.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1659 (.I0(n88), .I1(n87), .I2(n16485), 
            .I3(GND_net), .O(n16538));
    defparam i1_2_lut_3_lut_adj_1659.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1660 (.I0(n89), .I1(n88), .I2(n16541), 
            .I3(GND_net), .O(n16535));
    defparam i1_2_lut_3_lut_adj_1660.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1661 (.I0(n90), .I1(n89), .I2(n16538), 
            .I3(GND_net), .O(n16475));
    defparam i1_2_lut_3_lut_adj_1661.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4409));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33414_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n39736));
    defparam i33414_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4411));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4413));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33387_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n39709));
    defparam i33387_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4415));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4391));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n40969), .I1(n16502), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'hceef;
    SB_LUT4 i32805_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n39125));
    defparam i32805_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4393));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4395));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32811_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n39131));
    defparam i32811_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4370));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32848_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n39168));
    defparam i32848_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4372));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4374));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32861_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n39181));
    defparam i32861_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4351));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32896_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n39216));
    defparam i32896_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4353));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32910_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n39230));
    defparam i32910_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4355));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4329));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32961_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n39281));
    defparam i32961_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4331));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32967_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n39287));
    defparam i32967_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4333));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4311));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33022_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n39342));
    defparam i33022_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4313));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33051_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n39372));
    defparam i33051_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4315));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4299));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33110_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n39432));
    defparam i33110_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4301));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4287));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33133_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n39455));
    defparam i33133_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4289));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4275));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33153_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n39475));
    defparam i33153_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1596_3_lut (.I0(n2370), .I1(n6856), .I2(n2381), .I3(GND_net), 
            .O(n2460));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4277));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_78_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[1]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_107[1]), 
            .I2(n15), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13799_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n33766), 
            .I3(GND_net), .O(n18306));   // verilog/coms.v(126[12] 289[6])
    defparam i13799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22784_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4612));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i22784_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_3_lut_adj_1663 (.I0(n97), .I1(n96), .I2(n16520), 
            .I3(GND_net), .O(n16514));
    defparam i1_2_lut_3_lut_adj_1663.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut (.I0(n95), .I1(n94), .I2(n93), .I3(n16529), 
            .O(n16520));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(n94), .I1(n93), .I2(n16529), 
            .I3(GND_net), .O(n16523));
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1665 (.I0(n92), .I1(n91), .I2(n90), .I3(n16535), 
            .O(n16529));
    defparam i1_2_lut_4_lut_adj_1665.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1666 (.I0(n91), .I1(n90), .I2(n16535), 
            .I3(GND_net), .O(n16532));
    defparam i1_2_lut_3_lut_adj_1666.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n16472), 
            .O(n249));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 i4_4_lut_adj_1667 (.I0(n34307), .I1(n30686), .I2(n16809), 
            .I3(n6_adj_4567), .O(n35420));
    defparam i4_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 i13738_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13950), .I3(GND_net), .O(n18245));   // verilog/coms.v(126[12] 289[6])
    defparam i13738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14002_3_lut_4_lut (.I0(r_SM_Main_adj_4662[2]), .I1(r_SM_Main_adj_4662[0]), 
            .I2(r_SM_Main_2__N_3295[1]), .I3(r_SM_Main_adj_4662[1]), .O(n18509));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14002_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 div_46_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4453));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1048_3_lut (.I0(n1538), .I1(n6720), .I2(n1553), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33308_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n39630));
    defparam i33308_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1123_3_lut (.I0(n1652), .I1(n6733), .I2(n1667), .I3(GND_net), 
            .O(n1763));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4455));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_4_lut_adj_1668 (.I0(n16417), .I1(tx_active), .I2(r_SM_Main_2__N_3298[0]), 
            .I3(n25598), .O(n19_adj_4616));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_4_lut_adj_1668.LUT_INIT = 16'h5455;
    SB_LUT4 div_46_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4457));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33237_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n39559));
    defparam i33237_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1655_3_lut (.I0(n2460), .I1(n6877), .I2(n2471), .I3(GND_net), 
            .O(n2547));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33185_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n39507));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33185_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4268));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33197_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n39519));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33197_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4260));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4256));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33205_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n39527));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33205_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4251));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1196_3_lut (.I0(n1763), .I1(n6747), .I2(n1778), .I3(GND_net), 
            .O(n1871));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4459));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33215_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n39537));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33215_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4247));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33227_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n39549));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam i33227_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1592_3_lut (.I0(n2366), .I1(n6852), .I2(n2381), .I3(GND_net), 
            .O(n2456));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1267_3_lut (.I0(n1871), .I1(n6762), .I2(n1886), .I3(GND_net), 
            .O(n1976));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n17522), .O(n33396));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 div_46_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4475));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4479));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4587));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4586));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13393_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n34976), 
            .I3(GND_net), .O(n17900));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33169_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n39491));
    defparam i33169_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 communication_counter_31__I_0_i584_3_lut_4_lut (.I0(n36607), .I1(n746), 
            .I2(n11515), .I3(n852), .O(n954));
    defparam communication_counter_31__I_0_i584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 communication_counter_31__I_0_i585_3_lut_4_lut (.I0(n36607), .I1(n746), 
            .I2(n11516), .I3(n748), .O(n955));
    defparam communication_counter_31__I_0_i585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 communication_counter_31__I_0_i587_3_lut_4_lut (.I0(n36607), .I1(n746), 
            .I2(n11518), .I3(n855), .O(n957));
    defparam communication_counter_31__I_0_i587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 communication_counter_31__I_0_i586_rep_65_3_lut_4_lut (.I0(n36607), 
            .I1(n746), .I2(n11517), .I3(n749), .O(n956));
    defparam communication_counter_31__I_0_i586_rep_65_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1669 (.I0(control_mode[0]), .I1(n16421), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_3985));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i1_2_lut_3_lut_adj_1669.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1670 (.I0(control_mode[0]), .I1(n16421), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(186[5:22])
    defparam i1_2_lut_3_lut_adj_1670.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4481));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13800_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n33766), 
            .I3(GND_net), .O(n18307));   // verilog/coms.v(126[12] 289[6])
    defparam i13800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13801_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n33766), 
            .I3(GND_net), .O(n18308));   // verilog/coms.v(126[12] 289[6])
    defparam i13801_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4477));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33201_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n39523));
    defparam i33201_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4497));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4501));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4585));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4584));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33047_2_lut_4_lut (.I0(n2705_adj_4071), .I1(n84), .I2(n2714), 
            .I3(n93), .O(n39368));
    defparam i33047_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 communication_counter_31__I_0_i990_rep_58_3_lut (.I0(n1453), .I1(n1520), 
            .I2(n1481), .I3(GND_net), .O(n1552));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i990_rep_58_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i991_3_lut (.I0(n1454), .I1(n1521), 
            .I2(n1481), .I3(GND_net), .O(n1553_adj_4130));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i993_3_lut (.I0(n1456), .I1(n1523), 
            .I2(n1481), .I3(GND_net), .O(n1555));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i989_3_lut (.I0(n1452), .I1(n1519), 
            .I2(n1481), .I3(GND_net), .O(n1551));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i992_3_lut (.I0(n1455), .I1(n1522), 
            .I2(n1481), .I3(GND_net), .O(n1554_adj_4131));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i995_3_lut (.I0(n1458), .I1(n1525), 
            .I2(n1481), .I3(GND_net), .O(n1557));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705_adj_4071), 
            .I3(GND_net), .O(n14_adj_4503));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 communication_counter_31__I_0_i994_rep_59_3_lut (.I0(n1457), .I1(n1524), 
            .I2(n1481), .I3(GND_net), .O(n1556));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i994_rep_59_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i988_3_lut (.I0(n1451), .I1(n1518), 
            .I2(n1481), .I3(GND_net), .O(n1550));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i987_3_lut (.I0(n1450), .I1(n1517), 
            .I2(n1481), .I3(GND_net), .O(n1549));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i986_3_lut (.I0(n1449), .I1(n1516), 
            .I2(n1481), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1671 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n34642));
    defparam i1_3_lut_adj_1671.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1672 (.I0(n1554_adj_4131), .I1(n1551), .I2(n34642), 
            .I3(n1555), .O(n11_adj_4043));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i3_4_lut_adj_1672.LUT_INIT = 16'heccc;
    SB_LUT4 i5_4_lut_adj_1673 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_4042));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1674 (.I0(n13_adj_4042), .I1(n11_adj_4043), .I2(n1553_adj_4130), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i7_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4583));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_mux_3_i21_3_lut (.I0(communication_counter[20]), 
            .I1(n13_adj_3972), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1558));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4582));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4581));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4580));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4579));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_78_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[2]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_107[2]), 
            .I2(n15), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_78_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[3]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_107[3]), 
            .I2(n15), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4578));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4577));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1336_3_lut (.I0(n1976), .I1(n6778), .I2(n1991), .I3(GND_net), 
            .O(n2078));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1336_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4576));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4575));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_i919_3_lut (.I0(n1350), .I1(n1417_adj_4154), 
            .I2(n1382), .I3(GND_net), .O(n1449));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i923_3_lut (.I0(n1354), .I1(n1421), 
            .I2(n1382), .I3(GND_net), .O(n1453));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i927_3_lut (.I0(n1358), .I1(n1425), 
            .I2(n1382), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i925_3_lut (.I0(n1356), .I1(n1423), 
            .I2(n1382), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i924_3_lut (.I0(n1355), .I1(n1422), 
            .I2(n1382), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i922_3_lut (.I0(n1353), .I1(n1420_adj_4157), 
            .I2(n1382), .I3(GND_net), .O(n1452));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i920_3_lut (.I0(n1351), .I1(n1418_adj_4155), 
            .I2(n1382), .I3(GND_net), .O(n1450));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i921_3_lut (.I0(n1352), .I1(n1419_adj_4156), 
            .I2(n1382), .I3(GND_net), .O(n1451));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i926_rep_60_3_lut (.I0(n1357), .I1(n1424), 
            .I2(n1382), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i926_rep_60_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1675 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n36727));
    defparam i1_2_lut_adj_1675.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n1454), .I1(n36727), .I2(n1455), .I3(n1457), 
            .O(n34645));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1677 (.I0(n34645), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_4075));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1678 (.I0(n1453), .I1(n12_adj_4075), .I2(n1449), 
            .I3(n1448), .O(n1481));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i6_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i22_3_lut (.I0(communication_counter[21]), 
            .I1(n12_adj_3973), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1458));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4499));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4574));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33114_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n39436));
    defparam i33114_2_lut_4_lut.LUT_INIT = 16'hf99f;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n2731({n2732, n2733, n2734, 
            n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
            n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
            n2751, n2752, n2753, n2754, n2755}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .n18466(n18466), .clk32MHz(clk32MHz), .n18467(n18467), 
            .n18468(n18468), .n18469(n18469), .n18470(n18470), .n18471(n18471), 
            .n18451(n18451), .n18452(n18452), .n18472(n18472), .n18473(n18473), 
            .n18462(n18462), .n18463(n18463), .n18464(n18464), .n18465(n18465), 
            .n18453(n18453), .n18454(n18454), .n18455(n18455), .n18456(n18456), 
            .n18457(n18457), .n18458(n18458), .n18459(n18459), .n18460(n18460), 
            .n18461(n18461), .data_o({quadA_debounced, quadB_debounced}), 
            .count_enable(count_enable), .n17897(n17897), .n18498(n18498), 
            .n34976(n34976), .reg_B({reg_B}), .n17900(n17900), .PIN_2_c_0(PIN_2_c_0), 
            .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(212[15] 217[4])
    SB_LUT4 mux_78_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[4]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_107[4]), 
            .I2(n15), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4573));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13858_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n33775), .I3(GND_net), .O(n18365));   // verilog/coms.v(126[12] 289[6])
    defparam i13858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4572));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(130[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1403_3_lut (.I0(n2078), .I1(n6795), .I2(n2093), .I3(GND_net), 
            .O(n2177));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4571));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13404_3_lut (.I0(quadB_debounced_adj_4010), .I1(reg_B_adj_4672[0]), 
            .I2(n34961), .I3(GND_net), .O(n17911));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13415_4_lut (.I0(n17721), .I1(state[1]), .I2(state_3__N_337[1]), 
            .I3(n17561), .O(n17922));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13415_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i13425_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1035), .I3(GND_net), .O(n17932));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i855_3_lut (.I0(n1254), .I1(n1321), 
            .I2(n1283), .I3(GND_net), .O(n1353));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i854_3_lut (.I0(n1253), .I1(n1320), 
            .I2(n1283), .I3(GND_net), .O(n1352));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13919_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18426));   // verilog/coms.v(126[12] 289[6])
    defparam i13919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i857_3_lut (.I0(n1256), .I1(n1323), 
            .I2(n1283), .I3(GND_net), .O(n1355));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i856_3_lut (.I0(n1255), .I1(n1322), 
            .I2(n1283), .I3(GND_net), .O(n1354));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i853_3_lut (.I0(n1252), .I1(n1319), 
            .I2(n1283), .I3(GND_net), .O(n1351));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i852_3_lut (.I0(n1251), .I1(n1318), 
            .I2(n1283), .I3(GND_net), .O(n1350));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i859_3_lut (.I0(n1258), .I1(n1325), 
            .I2(n1283), .I3(GND_net), .O(n1357));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i858_rep_61_3_lut (.I0(n1257), .I1(n1324), 
            .I2(n1283), .I3(GND_net), .O(n1356));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i858_rep_61_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1679 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n34612));
    defparam i1_3_lut_adj_1679.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1680 (.I0(n1351), .I1(n1354), .I2(n34612), .I3(n1355), 
            .O(n8_adj_4062));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i2_4_lut_adj_1680.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1681 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4063));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i1_2_lut_adj_1681.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1682 (.I0(n1352), .I1(n7_adj_4063), .I2(n1353), 
            .I3(n8_adj_4062), .O(n1382));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i5_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i23_3_lut (.I0(communication_counter[22]), 
            .I1(n11_adj_3974), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n1358));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4570));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4569));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    \pwm(32000000,20000,32000000,23,1)  PWM (.VCC_net(VCC_net), .PIN_19_c_0(PIN_19_c_0), 
            .CLK_c(CLK_c), .\half_duty_new[0] (half_duty_new[0]), .n18513(n18513), 
            .\half_duty[0][2] (\half_duty[0] [2]), .n18514(n18514), .\half_duty[0][3] (\half_duty[0] [3]), 
            .n18515(n18515), .\half_duty[0][4] (\half_duty[0] [4]), .n18517(n18517), 
            .\half_duty[0][6] (\half_duty[0] [6]), .n18518(n18518), .\half_duty[0][7] (\half_duty[0] [7]), 
            .n18512(n18512), .\half_duty[0][1] (\half_duty[0] [1]), .GND_net(GND_net), 
            .n1035(n1035), .n17932(n17932), .\half_duty[0][0] (\half_duty[0] [0]), 
            .\half_duty_new[1] (half_duty_new[1]), .\half_duty_new[2] (half_duty_new[2]), 
            .\half_duty_new[3] (half_duty_new[3]), .\half_duty_new[4] (half_duty_new[4]), 
            .\half_duty_new[6] (half_duty_new[6]), .\half_duty_new[7] (half_duty_new[7]), 
            .pwm_setpoint({pwm_setpoint})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(112[43] 118[3])
    SB_LUT4 mux_78_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_3943), .I3(n15_adj_3985), .O(motor_state_23__N_107[5]));   // verilog/TinyFPGA_B.v(187[5] 190[10])
    defparam mux_78_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_77_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_107[5]), 
            .I2(n15), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(186[5] 190[10])
    defparam mux_77_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13918_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18425));   // verilog/coms.v(126[12] 289[6])
    defparam i13918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13436_3_lut (.I0(color[22]), .I1(blue[6]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17943));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1683 (.I0(bit_ctr[6]), .I1(n39069), .I2(n17536), 
            .I3(GND_net), .O(n32690));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1683.LUT_INIT = 16'hcaca;
    SB_LUT4 i13438_3_lut (.I0(color[21]), .I1(blue[5]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17945));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13439_3_lut (.I0(color[20]), .I1(blue[4]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17946));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13440_3_lut (.I0(color[19]), .I1(blue[3]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17947));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13441_3_lut (.I0(color[23]), .I1(blue[7]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17948));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13442_3_lut (.I0(color[18]), .I1(blue[2]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17949));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13443_3_lut (.I0(color[17]), .I1(blue[1]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17950));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2206_3_lut (.I0(n3245), .I1(n3312), 
            .I2(n3263), .I3(GND_net), .O(n3344));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2205_3_lut (.I0(n3244), .I1(n3311), 
            .I2(n3263), .I3(GND_net), .O(n3343));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n3246), .I1(n3343), .I2(n3313), .I3(n3263), 
            .O(n36643));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'hfcee;
    SB_LUT4 communication_counter_31__I_0_i2208_3_lut (.I0(n3247), .I1(n3314), 
            .I2(n3263), .I3(GND_net), .O(n3346));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2213_3_lut (.I0(n3252), .I1(n3319), 
            .I2(n3263), .I3(GND_net), .O(n3351));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n3249), .I1(n3351), .I2(n3316), .I3(n3263), 
            .O(n36693));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n36693), .I1(n3251), .I2(n3318), .I3(n3263), 
            .O(n36695));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n3242), .I1(n36695), .I2(n3309), .I3(n3263), 
            .O(n36697));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n3240), .I1(n36697), .I2(n3307), .I3(n3263), 
            .O(n36699));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n3239), .I1(n36699), .I2(n3306), .I3(n3263), 
            .O(n36701));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_2_lut_adj_1690 (.I0(n3356), .I1(n3358), .I2(GND_net), .I3(GND_net), 
            .O(n36953));
    defparam i1_2_lut_adj_1690.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n3253), .I1(n3344), .I2(n3320), .I3(n3263), 
            .O(n36641));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n36643), .I1(n3243), .I2(n3310), .I3(n3263), 
            .O(n36645));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'hfaee;
    SB_LUT4 communication_counter_31__I_0_i2202_3_lut (.I0(n3241), .I1(n3308), 
            .I2(n3263), .I3(GND_net), .O(n3340));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n3354), .I1(n36953), .I2(n3355), .I3(n3357), 
            .O(n34730));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n34730), .I1(n3340), .I2(n36645), .I3(n36641), 
            .O(n36651));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n3237), .I1(n36651), .I2(n3304), .I3(n3263), 
            .O(n36653));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n3236), .I1(n36701), .I2(n3303), .I3(n3263), 
            .O(n36703));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n3353), .I1(n3250), .I2(n3317), .I3(n3263), 
            .O(n36757));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'hfaee;
    SB_LUT4 i13929_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[6] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18436));   // verilog/coms.v(126[12] 289[6])
    defparam i13929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1698 (.I0(n3248), .I1(n3346), .I2(n3315), .I3(n3263), 
            .O(n28));
    defparam i3_4_lut_adj_1698.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n36703), .I1(n3235), .I2(n3302), .I3(n3263), 
            .O(n46_adj_4622));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n36653), .I1(n3233), .I2(n3300), .I3(n3263), 
            .O(n47_adj_4621));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hfaee;
    SB_LUT4 communication_counter_31__I_0_i2199_3_lut (.I0(n3238), .I1(n3305), 
            .I2(n3263), .I3(GND_net), .O(n3337));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n3234), .I1(n3337), .I2(n3301), .I3(n3263), 
            .O(n36613));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'hfcee;
    SB_LUT4 communication_counter_31__I_0_i2192_3_lut (.I0(n3231), .I1(n3298), 
            .I2(n3263), .I3(GND_net), .O(n3330));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n47_adj_4621), .I1(n46_adj_4622), .I2(n28), 
            .I3(n36757), .O(n36763));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n3232), .I1(n36613), .I2(n3299), .I3(n3263), 
            .O(n36615));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n37078), .I1(n36615), .I2(n36763), 
            .I3(n3330), .O(n3362));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i3_3_lut (.I0(communication_counter[2]), 
            .I1(n31_adj_3955), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n3358));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2217_3_lut (.I0(n3256), .I1(n3323), 
            .I2(n3263), .I3(GND_net), .O(n3355));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2215_3_lut (.I0(n3254), .I1(n3321), 
            .I2(n3263), .I3(GND_net), .O(n3353));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13928_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[6] [0]), 
            .I2(n35752), .I3(GND_net), .O(n18435));   // verilog/coms.v(126[12] 289[6])
    defparam i13928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2216_3_lut (.I0(n3255), .I1(n3322), 
            .I2(n3263), .I3(GND_net), .O(n3354));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33990_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i33990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13927_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[7] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18434));   // verilog/coms.v(126[12] 289[6])
    defparam i13927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33991_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i33991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2139_3_lut (.I0(n3146), .I1(n3213), 
            .I2(n3164), .I3(GND_net), .O(n3245));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2137_3_lut (.I0(n3144), .I1(n3211), 
            .I2(n3164), .I3(GND_net), .O(n3243));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2135_3_lut (.I0(n3142), .I1(n3209), 
            .I2(n3164), .I3(GND_net), .O(n3241));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13931_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[6] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18438));   // verilog/coms.v(126[12] 289[6])
    defparam i13931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2142_3_lut (.I0(n3149), .I1(n3216), 
            .I2(n3164), .I3(GND_net), .O(n3248));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33992_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i33992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33993_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i33993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2138_3_lut (.I0(n3145), .I1(n3212), 
            .I2(n3164), .I3(GND_net), .O(n3244));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2140_3_lut (.I0(n3147), .I1(n3214), 
            .I2(n3164), .I3(GND_net), .O(n3246));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2129_3_lut (.I0(n3136), .I1(n3203), 
            .I2(n3164), .I3(GND_net), .O(n3235));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2127_3_lut (.I0(n3134), .I1(n3201), 
            .I2(n3164), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2128_3_lut (.I0(n3135), .I1(n3202), 
            .I2(n3164), .I3(GND_net), .O(n3234));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2126_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3164), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2149_3_lut (.I0(n3156), .I1(n3223), 
            .I2(n3164), .I3(GND_net), .O(n3255));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2148_3_lut (.I0(n3155), .I1(n3222), 
            .I2(n3164), .I3(GND_net), .O(n3254));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2134_3_lut (.I0(n3141), .I1(n3208), 
            .I2(n3164), .I3(GND_net), .O(n3240));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34377_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34190_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2141_3_lut (.I0(n3148), .I1(n3215), 
            .I2(n3164), .I3(GND_net), .O(n3247));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2147_3_lut (.I0(n3154), .I1(n3221), 
            .I2(n3164), .I3(GND_net), .O(n3253));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2136_3_lut (.I0(n3143), .I1(n3210), 
            .I2(n3164), .I3(GND_net), .O(n3242));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2151_3_lut (.I0(n3158), .I1(n3225), 
            .I2(n3164), .I3(GND_net), .O(n3257));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2150_3_lut (.I0(n3157), .I1(n3224), 
            .I2(n3164), .I3(GND_net), .O(n3256));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2070_3_lut (.I0(n3045), .I1(n3112), 
            .I2(n3065), .I3(GND_net), .O(n3144));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34197_3_lut (.I0(n2953), .I1(n3020), .I2(n2966), .I3(GND_net), 
            .O(n3052));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2075_3_lut (.I0(n3050), .I1(n3117), 
            .I2(n3065), .I3(GND_net), .O(n3149));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2072_3_lut (.I0(n3047), .I1(n3114), 
            .I2(n3065), .I3(GND_net), .O(n3146));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2058_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3065), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_mux_3_i5_3_lut (.I0(communication_counter[4]), 
            .I1(n29_adj_3957), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n3158));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2083_3_lut (.I0(n3058), .I1(n3125), 
            .I2(n3065), .I3(GND_net), .O(n3157));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2082_3_lut (.I0(n3057), .I1(n3124), 
            .I2(n3065), .I3(GND_net), .O(n3156));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2071_3_lut (.I0(n3046), .I1(n3113), 
            .I2(n3065), .I3(GND_net), .O(n3145));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2071_3_lut.LUT_INIT = 16'hcaca;
    motorControl control (.GND_net(GND_net), .\Kp[6] (Kp[6]), .motor_state({motor_state}), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .setpoint({setpoint}), .\Kp[2] (Kp[2]), 
            .\Kp[7] (Kp[7]), .duty({duty}), .VCC_net(VCC_net), .PWMLimit({PWMLimit}), 
            .clk32MHz(clk32MHz), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .n41708(n41708)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(192[16] 205[4])
    SB_LUT4 div_46_i1468_3_lut (.I0(n2177), .I1(n6813), .I2(n2192), .I3(GND_net), 
            .O(n2273));   // verilog/TinyFPGA_B.v(208[21:53])
    defparam div_46_i1468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2073_3_lut (.I0(n3048), .I1(n3115), 
            .I2(n3065), .I3(GND_net), .O(n3147));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2069_3_lut (.I0(n3044), .I1(n3111), 
            .I2(n3065), .I3(GND_net), .O(n3143));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2066_3_lut (.I0(n3041), .I1(n3108), 
            .I2(n3065), .I3(GND_net), .O(n3140));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2065_3_lut (.I0(n3040), .I1(n3107), 
            .I2(n3065), .I3(GND_net), .O(n3139));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2064_3_lut (.I0(n3039), .I1(n3106), 
            .I2(n3065), .I3(GND_net), .O(n3138));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2062_3_lut (.I0(n3037), .I1(n3104), 
            .I2(n3065), .I3(GND_net), .O(n3136));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2061_3_lut (.I0(n3036), .I1(n3103), 
            .I2(n3065), .I3(GND_net), .O(n3135));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2060_3_lut (.I0(n3035), .I1(n3102), 
            .I2(n3065), .I3(GND_net), .O(n3134));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2059_3_lut (.I0(n3034), .I1(n3101), 
            .I2(n3065), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2079_3_lut (.I0(n3054), .I1(n3121), 
            .I2(n3065), .I3(GND_net), .O(n3153));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2068_3_lut (.I0(n3043), .I1(n3110), 
            .I2(n3065), .I3(GND_net), .O(n3142));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2074_3_lut (.I0(n3049), .I1(n3116), 
            .I2(n3065), .I3(GND_net), .O(n3148));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2009_rep_12_3_lut (.I0(n2952), 
            .I1(n3019), .I2(n2966), .I3(GND_net), .O(n3051));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2009_rep_12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34204_3_lut (.I0(n2947), .I1(n3014), .I2(n2966), .I3(GND_net), 
            .O(n3046));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i34204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2011_rep_14_3_lut (.I0(n2954), 
            .I1(n3021), .I2(n2966), .I3(GND_net), .O(n3053));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2011_rep_14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2008_3_lut (.I0(n2951), .I1(n3018), 
            .I2(n2966), .I3(GND_net), .O(n3050));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2003_3_lut (.I0(n2946), .I1(n3013), 
            .I2(n2966), .I3(GND_net), .O(n3045));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2006_3_lut (.I0(n2949), .I1(n3016), 
            .I2(n2966), .I3(GND_net), .O(n3048));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2002_3_lut (.I0(n2945), .I1(n3012), 
            .I2(n2966), .I3(GND_net), .O(n3044));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2001_3_lut (.I0(n2944), .I1(n3011), 
            .I2(n2966), .I3(GND_net), .O(n3043));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2007_3_lut (.I0(n2950), .I1(n3017), 
            .I2(n2966), .I3(GND_net), .O(n3049));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1995_3_lut (.I0(n2938), .I1(n3005), 
            .I2(n2966), .I3(GND_net), .O(n3037));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1993_3_lut (.I0(n2936), .I1(n3003), 
            .I2(n2966), .I3(GND_net), .O(n3035));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1994_3_lut (.I0(n2937), .I1(n3004), 
            .I2(n2966), .I3(GND_net), .O(n3036));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1992_3_lut (.I0(n2935), .I1(n3002), 
            .I2(n2966), .I3(GND_net), .O(n3034));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1999_3_lut (.I0(n2942), .I1(n3009), 
            .I2(n2966), .I3(GND_net), .O(n3041));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1997_3_lut (.I0(n2940), .I1(n3007), 
            .I2(n2966), .I3(GND_net), .O(n3039));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1998_3_lut (.I0(n2941), .I1(n3008), 
            .I2(n2966), .I3(GND_net), .O(n3040));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1996_3_lut (.I0(n2939), .I1(n3006), 
            .I2(n2966), .I3(GND_net), .O(n3038));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i1991_3_lut (.I0(n2934), .I1(n3001), 
            .I2(n2966), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2005_3_lut (.I0(n2948), .I1(n3015), 
            .I2(n2966), .I3(GND_net), .O(n3047));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2013_3_lut (.I0(n2956), .I1(n3023), 
            .I2(n2966), .I3(GND_net), .O(n3055));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2000_3_lut (.I0(n2943), .I1(n3010), 
            .I2(n2966), .I3(GND_net), .O(n3042));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2012_3_lut (.I0(n2955), .I1(n3022), 
            .I2(n2966), .I3(GND_net), .O(n3054));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13930_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[6] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18437));   // verilog/coms.v(126[12] 289[6])
    defparam i13930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_mux_3_i6_3_lut (.I0(communication_counter[5]), 
            .I1(n28_adj_3958), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n3058));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2015_3_lut (.I0(n2958), .I1(n3025), 
            .I2(n2966), .I3(GND_net), .O(n3057));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1705 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n34777));
    defparam i1_3_lut_adj_1705.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1706 (.I0(n3054), .I1(n3042), .I2(n34777), .I3(n3055), 
            .O(n29));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i6_4_lut_adj_1706.LUT_INIT = 16'heccc;
    SB_LUT4 i14_4_lut_adj_1707 (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37_adj_3952));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1708 (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i13_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1709 (.I0(n37_adj_3952), .I1(n29), .I2(n3049), 
            .I3(n3043), .O(n42_adj_3948));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i19_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1710 (.I0(n3044), .I1(n3048), .I2(n3045), .I3(n3052), 
            .O(n40_adj_3950));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1711 (.I0(n3047), .I1(n36), .I2(n3033), .I3(n3032), 
            .O(n41_adj_3949));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i18_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1712 (.I0(n3050), .I1(n3053), .I2(n3046), .I3(n3051), 
            .O(n39_adj_3951));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i16_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1713 (.I0(n39_adj_3951), .I1(n41_adj_3949), .I2(n40_adj_3950), 
            .I3(n42_adj_3948), .O(n3065));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i22_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i2014_3_lut (.I0(n2957), .I1(n3024), 
            .I2(n2966), .I3(GND_net), .O(n3056));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2081_3_lut (.I0(n3056), .I1(n3123), 
            .I2(n3065), .I3(GND_net), .O(n3155));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13933_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[6] [5]), 
            .I2(n35752), .I3(GND_net), .O(n18440));   // verilog/coms.v(126[12] 289[6])
    defparam i13933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2080_3_lut (.I0(n3055), .I1(n3122), 
            .I2(n3065), .I3(GND_net), .O(n3154));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2067_3_lut (.I0(n3042), .I1(n3109), 
            .I2(n3065), .I3(GND_net), .O(n3141));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1714 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n34725));
    defparam i1_3_lut_adj_1714.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1715 (.I0(n3141), .I1(n3154), .I2(n34725), .I3(n3155), 
            .O(n30));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i6_4_lut_adj_1715.LUT_INIT = 16'heaaa;
    SB_LUT4 i16_4_lut_adj_1716 (.I0(n3150), .I1(n3148), .I2(n3142), .I3(n3153), 
            .O(n40_adj_3941));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i16_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i13932_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[6] [4]), 
            .I2(n35752), .I3(GND_net), .O(n18439));   // verilog/coms.v(126[12] 289[6])
    defparam i13932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1717 (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i2_2_lut_adj_1717.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1718 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38_adj_3942));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i14_4_lut_adj_1718.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1719 (.I0(n3139), .I1(n40_adj_3941), .I2(n30), 
            .I3(n3140), .O(n44));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i20_4_lut_adj_1719.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1720 (.I0(n3143), .I1(n3147), .I2(n3152), .I3(n3145), 
            .O(n42_adj_3940));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i18_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1721 (.I0(n3132), .I1(n38_adj_3942), .I2(n26), 
            .I3(n3131), .O(n43_adj_3939));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i19_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1722 (.I0(n3146), .I1(n3149), .I2(n3151), .I3(n3144), 
            .O(n41));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i17_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41), .I1(n43_adj_3939), .I2(n42_adj_3940), 
            .I3(n44), .O(n3164));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_i2063_3_lut (.I0(n3038), .I1(n3105), 
            .I2(n3065), .I3(GND_net), .O(n3137));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2133_3_lut (.I0(n3140), .I1(n3207), 
            .I2(n3164), .I3(GND_net), .O(n3239));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2131_3_lut (.I0(n3138), .I1(n3205), 
            .I2(n3164), .I3(GND_net), .O(n3237));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2132_3_lut (.I0(n3139), .I1(n3206), 
            .I2(n3164), .I3(GND_net), .O(n3238));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2130_3_lut (.I0(n3137), .I1(n3204), 
            .I2(n3164), .I3(GND_net), .O(n3236));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13935_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[6] [7]), 
            .I2(n35752), .I3(GND_net), .O(n18442));   // verilog/coms.v(126[12] 289[6])
    defparam i13935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_31__I_0_i2125_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3164), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2146_3_lut (.I0(n3153), .I1(n3220), 
            .I2(n3164), .I3(GND_net), .O(n3252));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1723 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n34782));
    defparam i1_3_lut_adj_1723.LUT_INIT = 16'hfefe;
    SB_LUT4 i17_4_lut_adj_1724 (.I0(n3242), .I1(n3253), .I2(n3247), .I3(n3250), 
            .O(n42));
    defparam i17_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_LUT4 i13934_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[6] [6]), 
            .I2(n35752), .I3(GND_net), .O(n18441));   // verilog/coms.v(126[12] 289[6])
    defparam i13934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13937_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[5] [1]), 
            .I2(n35752), .I3(GND_net), .O(n18444));   // verilog/coms.v(126[12] 289[6])
    defparam i13937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1725 (.I0(n3240), .I1(n3254), .I2(n34782), .I3(n3255), 
            .O(n31_adj_3938));
    defparam i6_4_lut_adj_1725.LUT_INIT = 16'heaaa;
    SB_LUT4 i13_3_lut (.I0(n3252), .I1(n3231), .I2(n3230), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13936_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[5] [0]), 
            .I2(n35752), .I3(GND_net), .O(n18443));   // verilog/coms.v(126[12] 289[6])
    defparam i13936_3_lut.LUT_INIT = 16'hacac;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n18494(n18494), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n18495(n18495), .n18475(n18475), .n18476(n18476), 
            .n18477(n18477), .n18478(n18478), .n18479(n18479), .n18480(n18480), 
            .n18496(n18496), .n18497(n18497), .n18492(n18492), .n18493(n18493), 
            .n18490(n18490), .n18491(n18491), .n18488(n18488), .n18489(n18489), 
            .n18486(n18486), .n18487(n18487), .n18484(n18484), .n18485(n18485), 
            .n18481(n18481), .n18482(n18482), .n18483(n18483), .data_o({quadA_debounced_adj_4009, 
            quadB_debounced_adj_4010}), .count_enable(count_enable_adj_4011), 
            .n17899(n17899), .n2681({n2682, n2683, n2684, n2685, n2686, 
            n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
            n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
            n2703, n2704, n2705}), .GND_net(GND_net), .n18510(n18510), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B_adj_4672}), .PIN_7_c_1(PIN_7_c_1), 
            .n34961(n34961), .n17911(n17911)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(220[15] 225[4])
    SB_LUT4 i18_4_lut_adj_1726 (.I0(n3246), .I1(n3244), .I2(n3249), .I3(n3248), 
            .O(n43));
    defparam i18_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1727 (.I0(n3236), .I1(n3238), .I2(n3237), .I3(n3239), 
            .O(n40));
    defparam i15_4_lut_adj_1727.LUT_INIT = 16'hfffe;
    SB_LUT4 i13939_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[5] [3]), 
            .I2(n35752), .I3(GND_net), .O(n18446));   // verilog/coms.v(126[12] 289[6])
    defparam i13939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13938_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[5] [2]), 
            .I2(n35752), .I3(GND_net), .O(n18445));   // verilog/coms.v(126[12] 289[6])
    defparam i13938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21_4_lut_adj_1728 (.I0(n31_adj_3938), .I1(n42), .I2(n3241), 
            .I3(n3243), .O(n46));
    defparam i21_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1729 (.I0(n3232), .I1(n3234), .I2(n3233), .I3(n3235), 
            .O(n39));
    defparam i14_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1730 (.I0(n43), .I1(n3245), .I2(n38), .I3(n3251), 
            .O(n47));
    defparam i22_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 communication_counter_31__I_0_mux_3_i4_3_lut (.I0(communication_counter[3]), 
            .I1(n30_adj_3956), .I2(communication_counter[31]), .I3(GND_net), 
            .O(n3258));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2219_3_lut (.I0(n3258), .I1(n3325), 
            .I2(n3263), .I3(GND_net), .O(n3357));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_31__I_0_i2218_3_lut (.I0(n3257), .I1(n3324), 
            .I2(n3263), .I3(GND_net), .O(n3356));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam communication_counter_31__I_0_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33276_3_lut (.I0(n10709), .I1(n10708), .I2(n10710), .I3(GND_net), 
            .O(n39045));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i33276_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1731 (.I0(n3356), .I1(n3357), .I2(GND_net), .I3(GND_net), 
            .O(n37047));
    defparam i1_2_lut_adj_1731.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut_adj_1732 (.I0(n2951), .I1(n2948), .I2(n2946), .I3(n2945), 
            .O(n38_adj_4549));   // verilog/TinyFPGA_B.v(50[6:33])
    defparam i16_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 i33254_4_lut (.I0(n39045), .I1(n10705), .I2(n10706), .I3(n10707), 
            .O(n39042));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i33254_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33279_4_lut (.I0(n3354), .I1(n3353), .I2(n3355), .I3(n3358), 
            .O(n39047));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i33279_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47_4_lut (.I0(n39047), .I1(n39042), .I2(n3362), .I3(n37047), 
            .O(n34555));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i47_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i33403_2_lut (.I0(communication_counter[0]), .I1(communication_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n39040));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i33403_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46_4_lut (.I0(n39040), .I1(n39038), .I2(communication_counter[31]), 
            .I3(n34555), .O(color_23__N_34));   // verilog/TinyFPGA_B.v(50[6:36])
    defparam i46_4_lut.LUT_INIT = 16'h3035;
    SB_LUT4 i13444_3_lut (.I0(color[16]), .I1(blue[0]), .I2(color_23__N_34), 
            .I3(GND_net), .O(n17951));   // verilog/TinyFPGA_B.v(47[8] 55[4])
    defparam i13444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13445_3_lut (.I0(setpoint[23]), .I1(n4446), .I2(n36216), 
            .I3(GND_net), .O(n17952));   // verilog/coms.v(126[12] 289[6])
    defparam i13445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13446_3_lut (.I0(setpoint[22]), .I1(n4445), .I2(n36216), 
            .I3(GND_net), .O(n17953));   // verilog/coms.v(126[12] 289[6])
    defparam i13446_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (timer, clk32MHz, n32678, VCC_net, bit_ctr, GND_net, 
            n32688, n32680, n32744, n32746, n32748, n32682, n32734, 
            n32736, n32738, n32742, n32730, n32732, n32726, n32728, 
            n32722, n32724, n32718, n32720, n32684, start, n32716, 
            n32714, n32686, n39074, n19, n39095, \state[0] , n155, 
            n39081, n39092, n39091, n39090, \state[1] , n37153, 
            n39089, n39088, n32712, n18052, \neo_pixel_transmitter.t0 , 
            n18051, n18050, n18049, n18048, n18047, n18046, n18045, 
            n18044, n18043, n18042, n18041, n18040, n18039, n18038, 
            n18037, n18036, n18035, n18034, n18033, n18032, n18031, 
            n18030, n18029, n18028, n18027, n18026, n18025, n18024, 
            n18023, n32710, n32708, n39080, n39087, n39094, n32702, 
            n32700, n32694, n32698, n32696, n18000, n32692, n39079, 
            n39086, n39093, n39085, n39070, n32690, n17922, n39084, 
            n39083, n39069, \state_3__N_337[1] , n131, n17536, n39082, 
            n21, n17792, n17561, n17721, n39078, n39077, n39072, 
            n39071, \color[16] , \color[17] , \color[18] , \color[19] , 
            \color[22] , \color[23] , \color[20] , \color[21] , n39067, 
            n39065, n39068, n39073, n39064, PIN_8_c, n39063, n39076, 
            n39075, n175, n39062) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [31:0]timer;
    input clk32MHz;
    input n32678;
    input VCC_net;
    output [31:0]bit_ctr;
    input GND_net;
    input n32688;
    input n32680;
    input n32744;
    input n32746;
    input n32748;
    input n32682;
    input n32734;
    input n32736;
    input n32738;
    input n32742;
    input n32730;
    input n32732;
    input n32726;
    input n32728;
    input n32722;
    input n32724;
    input n32718;
    input n32720;
    input n32684;
    output start;
    input n32716;
    input n32714;
    input n32686;
    output n39074;
    input n19;
    output n39095;
    output \state[0] ;
    output n155;
    output n39081;
    output n39092;
    output n39091;
    output n39090;
    output \state[1] ;
    output n37153;
    output n39089;
    output n39088;
    input n32712;
    input n18052;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n18051;
    input n18050;
    input n18049;
    input n18048;
    input n18047;
    input n18046;
    input n18045;
    input n18044;
    input n18043;
    input n18042;
    input n18041;
    input n18040;
    input n18039;
    input n18038;
    input n18037;
    input n18036;
    input n18035;
    input n18034;
    input n18033;
    input n18032;
    input n18031;
    input n18030;
    input n18029;
    input n18028;
    input n18027;
    input n18026;
    input n18025;
    input n18024;
    input n18023;
    input n32710;
    input n32708;
    output n39080;
    output n39087;
    output n39094;
    input n32702;
    input n32700;
    input n32694;
    input n32698;
    input n32696;
    input n18000;
    input n32692;
    output n39079;
    output n39086;
    output n39093;
    output n39085;
    output n39070;
    input n32690;
    input n17922;
    output n39084;
    output n39083;
    output n39069;
    output \state_3__N_337[1] ;
    output n131;
    output n17536;
    output n39082;
    output n21;
    input n17792;
    output n17561;
    output n17721;
    output n39078;
    output n39077;
    output n39072;
    output n39071;
    input \color[16] ;
    input \color[17] ;
    input \color[18] ;
    input \color[19] ;
    input \color[22] ;
    input \color[23] ;
    input \color[20] ;
    input \color[21] ;
    output n39067;
    output n39065;
    output n39068;
    output n39073;
    output n39064;
    output PIN_8_c;
    output n39063;
    output n39076;
    output n39075;
    output n175;
    output n39062;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n28649, n1501, n1532, n28650, n2890, n2791, n2819, n28880, 
        n28881, n2891, n2792, n28879, n4;
    wire [31:0]n1;
    
    wire n27636;
    wire [31:0]one_wire_N_488;
    
    wire \neo_pixel_transmitter.done_N_545 , n33752, \neo_pixel_transmitter.done , 
        n2892, n2793, n28878, n1601, n1502, n28648, n1602, n1503, 
        n28647, n1603, n1504, n28646, n2893, n2794, n28877, n27637, 
        n35812, n2894, n2795, n28876, n1604, n1505, n28645, n2895, 
        n2796, n28875, n1605, n1506, n28644, n2896, n2797, n28874, 
        n1606, n1507, n28643, n1607, n1508, n28642, n2897, n2798, 
        n28873, n1608, n1509, n41703, n28641, n2898, n2799, n28872, 
        n1609, n2899, n2800, n28871, n1499, n1400, n1433, n28640, 
        n1500, n1401, n28639, n2900, n2801, n28870, n1402, n28638, 
        n2901, n2802, n28869, n1403, n28637, n2902, n2803, n28868, 
        n1404, n28636, n2903, n2804, n28867, n1405, n28635, n1406, 
        n28634, n2904, n2805, n28866, n1407, n28633, n2905, n2806, 
        n28865, n1408, n28632, n2302, n2292, n22, n2299, n2309, 
        n30, n2294, n2306, n2297, n34, n2301, n2307, n2291, 
        n2305, n32_adj_3797, n2298, n2295, n2304, n2300, n33_adj_3798, 
        n2308, n2296, n2303, n2293, n31, n2324, n2423, n41714, 
        n2906, n2807, n28864, n1409, n41705, n28631, n2907, n2808, 
        n28863, n2908, n2809, n41704, n28862, n27458, n27450, 
        n2909, n2786, n2687, n2720, n28861, n2787, n2688, n28860, 
        n1301, n1334, n28630, n2788, n2689, n28859, n2789, n2690, 
        n28858, n1302, n28629, n1303, n28628, n2790, n2691, n28857, 
        n2692, n28856, n2693, n28855, n1304, n28627, n1305, n28626, 
        n2694, n28854, n1306, n28625, n25, n27, n29, n26, n16, 
        n2695, n28853, n1307, n28624, n1308, n28623, n21_c, n28, 
        n30_adj_3799, n23, n17, n22_adj_3800, n24, n16437, n24843, 
        n25384, n57, n136, n165, n37097, n2696, n28852, n2697, 
        n28851, n1309, n41707, n28622, n2698, n28850, n2699, n28849, 
        n2700, n28848, n1202, n1235, n28621, n1203, n28620, n2701, 
        n28847, n1204, n28619, n1205, n28618, n2702, n28846, n1206, 
        n28617, n1207, n28616, n1208, n28615, n2703, n28845, n2704, 
        n28844, n1209, n41709, n28614, n1103, n1136, n28613, n2705, 
        n28843, n1104, n28612, n2706, n28842, n27459, n2707, n28841, 
        n2708, n28840, n2709, n41706, n28839, n1105, n28611, n2588, 
        n2621, n28838, n1106, n28610, n2589, n28837, n2590, n28836, 
        n2591, n28835, n1107, n28609, n1108, n28608, n2592, n28834, 
        n1109, n41710, n28607, n4_adj_3801, n28606, n1037;
    wire [31:0]n1070;
    
    wire n1005, n28605, n2593, n28833, n2594, n28832, n1006, n28604, 
        n1007, n28603, n2595, n28831, n1008, n28602, n2596, n28830, 
        n1009, n28601, n27451, n2597, n28829, n905, n28600, n41690;
    wire [31:0]n971;
    
    wire n906, n28599, n34363, n28598, n2598, n28828, n17645, 
        n28597, n2599, n28827, n2600, n28826, n15165, n28596, 
        n2601, n28825, n2602, n28824, n27457, n2603, n28823, n2604, 
        n28822, n2605, n28821, n2606, n28820, n2607, n28819, n2608, 
        n28818, n2609, n41711, n28817, n2489, n2522, n28816, n2490, 
        n28815, n2491, n28814, n2492, n28813, n2493, n28812, n27478, 
        n2494, n28811;
    wire [31:0]n133;
    
    wire n28343, n28342, n28341, n2495, n28810, n2496, n28809, 
        n28340, n2497, n28808, n28339, n2498, n28807, n2499, n28806, 
        n28338, n28337, n28336, n28335, n2500, n28805, n2501, 
        n28804, n2502, n28803, n27477, n28334, n2503, n28802, 
        n2504, n28801, n28333, n2505, n28800, n28332, n2506, n28799, 
        n2507, n28798, n28331, n27476, n166, n168, n2508, n28797, 
        n28330, n28329, n2509, n41712, n28796, n28328, n28327, 
        n27475, n2390, n28795, n2391, n28794, n28326, n27474, 
        n2392, n28793, n28325, n28324, n2406, n2402, n22_adj_3803, 
        n2395, n2408, n2394, n2399, n32_adj_3804, n2409, n25276, 
        n2404, n2393, n36, n2407, n2398, n2401, n2405, n34_adj_3806, 
        n28792, n2397, n35, n2403, n2396, n2400, n33_adj_3807, 
        n28323, n28791, n28322, n28790, n27456, n27473, n27449, 
        n28789, n28321, n28788, n28787, n28786, n28320, n28319, 
        n28785, n28784, n28318, n28783, n28782, n28781, n28780, 
        n28317, n28316, n28779, n28315, n28778, n27455, n28314, 
        n27472, n25466, n16_adj_3809, n17_adj_3810, n28313, n28777, 
        n27448, n27471, n28776, n27454, n28775, n28774, n28773, 
        n28772, n24_adj_3811, n34_adj_3812, n22_adj_3813, n38, n36_adj_3814, 
        n37, n35_adj_3815, n30590, n36_adj_3816, n25_adj_3817, n34_adj_3818, 
        n40, n38_adj_3819, n39, n37_adj_3820, n27470, n28771, n28770, 
        n28769, n838, n807, n60, n28768, n28767, n28766, n28765, 
        n28764, n28763, n28762, n28761, n28760, n28759, n28758, 
        n41715, n28757, n2192, n2225, n28756, n2193, n28755, n2194, 
        n28754, n2195, n28753, n2196, n28752, n62, n2197, n28751, 
        n8, n34512, n7, n25502, n12, n2198, n28750, n2199, n28749, 
        n2200, n28748, n2201, n28747, n27469, n2202, n28746, n2203, 
        n28745, n2204, n28744, n14, n9, n30_adj_3821, n27453, 
        n48, n46, n47, n45, n44, n2205, n28743, n43, n54, 
        n49, n2206, n28742, n34361, n2207, n28741, n37149, n4488, 
        n40_adj_3822, n2208, n28740, n2209, n41716, n28739, n2093, 
        n2126, n28738, n2094, n28737, n2095, n28736, n2096, n28735, 
        n2097, n28734, n27468, n2098, n28733, n14_adj_3823, n12_adj_3824, 
        n16_adj_3825, n28_adj_3826, n9_adj_3827, n11, n10, n19765, 
        n38_adj_3829, n2099, n28732, n2100, n28731, n2101, n28730, 
        n25258, n2102, n28729, n2103, n28728, n36_adj_3830, n3182, 
        n3083, n3116, n28963, n2104, n28727, n3183, n3084, n28962, 
        n2105, n28726, n3184, n3085, n28961, n2106, n28725, n3185, 
        n3086, n28960, n3186, n3087, n28959, n26_adj_3831, n2107, 
        n28724;
    wire [3:0]state_3__N_337;
    
    wire n2108, n28723, n3187, n3088, n28958, n2109, n41717, n28722, 
        n3188, n3089, n28957, n1994, n2027, n28721, n1995, n28720, 
        n3189, n3090, n28956, n1996, n28719, n3190, n3091, n28955, 
        n1997, n28718, n3191, n3092, n28954, n3192, n3093, n28953, 
        n1998, n28717, n3193, n3094, n28952, n27467, n3194, n3095, 
        n28951, n1999, n28716, n3195, n3096, n28950, n2000, n28715, 
        n3196, n3097, n28949, n2001, n28714, n3197, n3098, n28948, 
        n2002, n28713, n27466, n42, n3198, n3099, n28947, n40_adj_3832, 
        n2003, n28712, n3199, n3100, n28946, n2004, n28711, n2005, 
        n28710, n3200, n3101, n28945, n2006, n28709, n3201, n3102, 
        n28944, n2007, n28708, n3202, n3103, n28943, n3203, n3104, 
        n28942, n2008, n28707, n3204, n3105, n28941, n2009, n41720, 
        n28706, n3205, n3106, n28940, n41, n3206, n3107, n28939, 
        n1895, n1928, n28705, n1896, n28704, n3207, n3108, n28938, 
        n3208, n3109, n41719, n28937, n1897, n28703, n3209, n1898, 
        n28702, n39_adj_3833, n2984, n3017, n28936, n27465, n1899, 
        n28701, n2985, n28935, n1900, n28700, n27464, n38_adj_3834, 
        n2986, n28934, n2987, n28933, n1901, n28699, n1902, n28698, 
        n2988, n28932, n1903, n28697, n2989, n28931, n1904, n28696, 
        n2990, n28930, n2991, n28929, n1905, n28695, n2992, n28928, 
        n1906, n28694, n2993, n28927, n2994, n28926, n1907, n28693, 
        n2995, n28925, n1908, n28692, n1909, n41721, n28691, n37309, 
        n2996, n28924, n37310, n37367, n2997, n28923, n37366, 
        n2998, n28922, n1796, n1829, n28690, n1797, n28689, n2999, 
        n28921, n1798, n28688, n39_adj_3840, n3000, n28920, n1799, 
        n28687, n3001, n28919, n1800, n28686, n1801, n28685, n3002, 
        n28918, n1802, n28684, n3003, n28917, n1803, n28683, n3004, 
        n28916, n27463, n1804, n28682, n3005, n28915, n1805, n28681, 
        n3006, n28914, n1806, n28680, n3007, n28913, n1807, n28679, 
        n3008, n28912, n1808, n28678, n3009, n41722, n28911, n1809, 
        n41723, n28677, n1631, n41726, n2885, n2918, n28910, n1697, 
        n1730, n28676, n2886, n28909, n1698, n28675, n1699, n28674, 
        n2887, n28908, n41724, n1700, n28673, n2888, n28907, n1701, 
        n28672, n37_adj_3851, n1702, n28671, n2889, n28906, n27452, 
        n27462, n1703, n28670, n28905, n28904, n1704, n28669, 
        n1705, n28668, n28903, n1706, n28667, n34_adj_3858, n28902, 
        n1707, n28666, n28901, n28900, n1708, n28665, n42_adj_3859, 
        n46_adj_3860, n1709, n41725, n28664, n28899, n28898, n28897, 
        n28896, n35817, n27461, n1598, n28663, n1599, n28662, 
        n17503, n28895, n1600, n28661, \neo_pixel_transmitter.done_N_551 , 
        n33686, n27666, n28894, n27665, n28660, n27664, n27663, 
        n28893, n28659, n33_adj_3862, n20_adj_3863, n27662, n13_adj_3864, 
        n28892, n18_adj_3865, n22_adj_3866, n27661, n27660, n28658, 
        n28891, n28890, n27659, n28657, n28889, n28656, n27658, 
        n27657, n28888, n28887, n27656, n28655, n27655, n28886, 
        n27654, n28654, n27653, n27652, n28885, n27651, n28884, 
        n27650, n27460, n27649, n28883, n28653, n28882, n28652, 
        n27648, n27647, n27646, n27645, n28651, n27644, n27643, 
        n27642, n27641, n27640, n27639, n27638, n18_adj_3867, n22_adj_3868, 
        n20_adj_3869, n21_adj_3870, n19_adj_3871, n34_adj_3872, n41_adj_3873, 
        n38_adj_3874, n43_adj_3875, n40_adj_3876, n46_adj_3877, n39_adj_3878, 
        n47_adj_3879, n24_adj_3880, n22_adj_3881, n23_adj_3882, n21_adj_3883, 
        n40_adj_3884, n44_adj_3885, n42_adj_3886, n43_adj_3887, n41_adj_3888, 
        n38_adj_3889, n46_adj_3890, n50, n37_adj_3891, n26_adj_3892, 
        n24_adj_3893, n25_adj_3894, n23_adj_3895, n18_adj_3896, n28_adj_3897, 
        n26_adj_3898, n27_adj_3899, n25_adj_3900, n25528, n48_adj_3901, 
        n46_adj_3902, n47_adj_3903, n45_adj_3904, n44_adj_3905, n43_adj_3906, 
        n54_adj_3907, n49_adj_3908, n25560, n41779, n5_adj_3909, n42_adj_3910, 
        n46_adj_3911, n44_adj_3912, n45_adj_3913, n43_adj_3914, n40_adj_3915, 
        n20_adj_3916, n48_adj_3917, n52, n39_adj_3918, n15_adj_3919, 
        n29806, n15157, n18_adj_3920, n25344, n30_adj_3921, n28_adj_3922, 
        n29_adj_3923, n27_adj_3924, n7534, n41776, n708, n28_adj_3925, 
        n32_adj_3926, n30_adj_3927, n31_adj_3928, n29_adj_3929;
    
    SB_CARRY mod_5_add_1071_11 (.CI(n28649), .I0(n1501), .I1(n1532), .CO(n28650));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n28880), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n28880), .I0(n2791), .I1(n2819), .CO(n28881));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n28879), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n28879), .I0(n2792), .I1(n2819), .CO(n28880));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_488[2]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n27636), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n33752), .D(\neo_pixel_transmitter.done_N_545 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n28878), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n28648), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n28878), .I0(n2793), .I1(n2819), .CO(n28879));
    SB_CARRY mod_5_add_1071_10 (.CI(n28648), .I0(n1502), .I1(n1532), .CO(n28649));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n28647), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(VCC_net), 
            .D(n32678));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1071_9 (.CI(n28647), .I0(n1503), .I1(n1532), .CO(n28648));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n28646), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n28877), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n27636), .I0(timer[1]), .I1(n1[1]), .CO(n27637));
    SB_LUT4 sub_14_add_2_2_lut (.I0(n4), .I1(timer[0]), .I2(n1[0]), .I3(VCC_net), 
            .O(n35812)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n27636));
    SB_CARRY mod_5_add_1942_18 (.CI(n28877), .I0(n2794), .I1(n2819), .CO(n28878));
    SB_CARRY mod_5_add_1071_8 (.CI(n28646), .I0(n1504), .I1(n1532), .CO(n28647));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n28876), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n28876), .I0(n2795), .I1(n2819), .CO(n28877));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n28645), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n28645), .I0(n1505), .I1(n1532), .CO(n28646));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n28875), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n28644), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n28644), .I0(n1506), .I1(n1532), .CO(n28645));
    SB_CARRY mod_5_add_1942_16 (.CI(n28875), .I0(n2796), .I1(n2819), .CO(n28876));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n28874), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n28643), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n28643), .I0(n1507), .I1(n1532), .CO(n28644));
    SB_CARRY mod_5_add_1942_15 (.CI(n28874), .I0(n2797), .I1(n2819), .CO(n28875));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n28642), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n28873), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n28642), .I0(n1508), .I1(n1532), .CO(n28643));
    SB_CARRY mod_5_add_1942_14 (.CI(n28873), .I0(n2798), .I1(n2819), .CO(n28874));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n41703), 
            .I3(n28641), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n28872), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_3 (.CI(n28641), .I0(n1509), .I1(n41703), .CO(n28642));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n41703), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_13 (.CI(n28872), .I0(n2799), .I1(n2819), .CO(n28873));
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n41703), 
            .CO(n28641));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n28871), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28640), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n28871), .I0(n2800), .I1(n2819), .CO(n28872));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28639), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n28870), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28639), .I0(n1401), .I1(n1433), .CO(n28640));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28638), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n28870), .I0(n2801), .I1(n2819), .CO(n28871));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n28869), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n28638), .I0(n1402), .I1(n1433), .CO(n28639));
    SB_CARRY mod_5_add_1942_10 (.CI(n28869), .I0(n2802), .I1(n2819), .CO(n28870));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28637), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n28637), .I0(n1403), .I1(n1433), .CO(n28638));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n28868), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28636), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n28868), .I0(n2803), .I1(n2819), .CO(n28869));
    SB_CARRY mod_5_add_1004_8 (.CI(n28636), .I0(n1404), .I1(n1433), .CO(n28637));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n28867), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28635), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n28867), .I0(n2804), .I1(n2819), .CO(n28868));
    SB_CARRY mod_5_add_1004_7 (.CI(n28635), .I0(n1405), .I1(n1433), .CO(n28636));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28634), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n28866), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28634), .I0(n1406), .I1(n1433), .CO(n28635));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28633), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n28866), .I0(n2805), .I1(n2819), .CO(n28867));
    SB_CARRY mod_5_add_1004_5 (.CI(n28633), .I0(n1407), .I1(n1433), .CO(n28634));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n28865), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28632), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut (.I0(bit_ctr[12]), .I1(n22), .I2(n2299), .I3(n2309), 
            .O(n30));
    defparam i11_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut (.I0(n2294), .I1(n30), .I2(n2306), .I3(n2297), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_3797));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_3798));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33_adj_3798), .I2(n32_adj_3797), 
            .I3(n34), .O(n2324));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFE bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(VCC_net), 
            .D(n32688));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(VCC_net), 
            .D(n32680));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i35394_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41714));
    defparam i35394_1_lut.LUT_INIT = 16'h5555;
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n32744));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n32746));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n32748));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(VCC_net), 
            .D(n32682));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n32734));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n32736));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n32738));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n32742));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n32730));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n32732));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n32726));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n32728));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n32722));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n32724));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n32718));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n32720));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n32684));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n32716));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n32714));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(VCC_net), 
            .D(n32686));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_6 (.CI(n28865), .I0(n2806), .I1(n2819), .CO(n28866));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n28864), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28632), .I0(n1408), .I1(n1433), .CO(n28633));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n41705), 
            .I3(n28631), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n28631), .I0(n1409), .I1(n41705), .CO(n28632));
    SB_CARRY mod_5_add_1942_5 (.CI(n28864), .I0(n2807), .I1(n2819), .CO(n28865));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n28863), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n28863), .I0(n2808), .I1(n2819), .CO(n28864));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n41704), 
            .I3(n28862), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_13_lut (.I0(n19), .I1(bit_ctr[11]), .I2(GND_net), .I3(n27458), 
            .O(n39074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n27450), 
            .O(n39095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_3 (.CI(n28862), .I0(n2809), .I1(n41704), .CO(n28863));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n41704), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n41704), 
            .CO(n28862));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n28861), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n41705), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n28860), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n41705), 
            .CO(n28631));
    SB_CARRY mod_5_add_1875_24 (.CI(n28860), .I0(n2688), .I1(n2720), .CO(n28861));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28630), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n28859), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n28859), .I0(n2689), .I1(n2720), .CO(n28860));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n28858), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28629), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n28858), .I0(n2690), .I1(n2720), .CO(n28859));
    SB_CARRY mod_5_add_937_10 (.CI(n28629), .I0(n1302), .I1(n1334), .CO(n28630));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28628), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n28857), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28628), .I0(n1303), .I1(n1334), .CO(n28629));
    SB_CARRY mod_5_add_1875_21 (.CI(n28857), .I0(n2691), .I1(n2720), .CO(n28858));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n28856), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n28856), .I0(n2692), .I1(n2720), .CO(n28857));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n28855), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n28855), .I0(n2693), .I1(n2720), .CO(n28856));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28627), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n28627), .I0(n1304), .I1(n1334), .CO(n28628));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28626), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n28854), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n28626), .I0(n1305), .I1(n1334), .CO(n28627));
    SB_CARRY mod_5_add_1875_18 (.CI(n28854), .I0(n2694), .I1(n2720), .CO(n28855));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28625), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut (.I0(n25), .I1(n27), .I2(n29), .I3(n26), .O(n16));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n28853), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n28853), .I0(n2695), .I1(n2720), .CO(n28854));
    SB_CARRY mod_5_add_937_6 (.CI(n28625), .I0(n1306), .I1(n1334), .CO(n28626));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28624), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28624), .I0(n1307), .I1(n1334), .CO(n28625));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28623), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut (.I0(n21_c), .I1(n28), .I2(n30_adj_3799), .I3(n23), 
            .O(n17));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n22_adj_3800), .I2(n16), .I3(n24), 
            .O(n16437));   // verilog/neopixel.v(104[14:39])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20897_3_lut (.I0(n16437), .I1(one_wire_N_488[11]), .I2(n24843), 
            .I3(GND_net), .O(n25384));
    defparam i20897_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(n57), .I2(GND_net), .I3(GND_net), 
            .O(n155));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15267_3_lut (.I0(n136), .I1(n165), .I2(\state[0] ), .I3(GND_net), 
            .O(n37097));   // verilog/neopixel.v(16[20:25])
    defparam i15267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n28852), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n28852), .I0(n2696), .I1(n2720), .CO(n28853));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n28851), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n28623), .I0(n1308), .I1(n1334), .CO(n28624));
    SB_CARRY mod_5_add_1875_15 (.CI(n28851), .I0(n2697), .I1(n2720), .CO(n28852));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n41707), 
            .I3(n28622), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n28622), .I0(n1309), .I1(n41707), .CO(n28623));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n28850), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n41707), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_14 (.CI(n28850), .I0(n2698), .I1(n2720), .CO(n28851));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n28849), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n41707), 
            .CO(n28622));
    SB_CARRY mod_5_add_1875_13 (.CI(n28849), .I0(n2699), .I1(n2720), .CO(n28850));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n28848), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28621), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28620), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n28848), .I0(n2700), .I1(n2720), .CO(n28849));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n28847), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28620), .I0(n1203), .I1(n1235), .CO(n28621));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28619), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28619), .I0(n1204), .I1(n1235), .CO(n28620));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28618), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n28847), .I0(n2701), .I1(n2720), .CO(n28848));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n28846), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28618), .I0(n1205), .I1(n1235), .CO(n28619));
    SB_CARRY mod_5_add_1875_10 (.CI(n28846), .I0(n2702), .I1(n2720), .CO(n28847));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28617), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28617), .I0(n1206), .I1(n1235), .CO(n28618));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28616), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n28616), .I0(n1207), .I1(n1235), .CO(n28617));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28615), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n28845), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n28615), .I0(n1208), .I1(n1235), .CO(n28616));
    SB_CARRY mod_5_add_1875_9 (.CI(n28845), .I0(n2703), .I1(n2720), .CO(n28846));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n28844), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n41709), 
            .I3(n28614), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n28614), .I0(n1209), .I1(n41709), .CO(n28615));
    SB_CARRY mod_5_add_1875_8 (.CI(n28844), .I0(n2704), .I1(n2720), .CO(n28845));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n41709), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n41709), 
            .CO(n28614));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28613), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n28843), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28612), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n28843), .I0(n2705), .I1(n2720), .CO(n28844));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n28842), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n27458), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27459));
    SB_CARRY mod_5_add_803_8 (.CI(n28612), .I0(n1104), .I1(n1136), .CO(n28613));
    SB_CARRY mod_5_add_1875_6 (.CI(n28842), .I0(n2706), .I1(n2720), .CO(n28843));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n28841), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n28841), .I0(n2707), .I1(n2720), .CO(n28842));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n28840), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n28840), .I0(n2708), .I1(n2720), .CO(n28841));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n41706), 
            .I3(n28839), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n28839), .I0(n2709), .I1(n41706), .CO(n28840));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28611), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n41706), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n41706), 
            .CO(n28839));
    SB_CARRY mod_5_add_803_7 (.CI(n28611), .I0(n1105), .I1(n1136), .CO(n28612));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n28838), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28610), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n28837), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n28837), .I0(n2589), .I1(n2621), .CO(n28838));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n28836), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28610), .I0(n1106), .I1(n1136), .CO(n28611));
    SB_CARRY mod_5_add_1808_22 (.CI(n28836), .I0(n2590), .I1(n2621), .CO(n28837));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n28835), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28609), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28609), .I0(n1107), .I1(n1136), .CO(n28610));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28608), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28608), .I0(n1108), .I1(n1136), .CO(n28609));
    SB_CARRY mod_5_add_1808_21 (.CI(n28835), .I0(n2591), .I1(n2621), .CO(n28836));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n28834), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n41710), 
            .I3(n28607), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n28607), .I0(n1109), .I1(n41710), .CO(n28608));
    SB_CARRY mod_5_add_1808_20 (.CI(n28834), .I0(n2592), .I1(n2621), .CO(n28835));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n41710), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n41710), 
            .CO(n28607));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n1037), .I1(n4_adj_3801), .I2(VCC_net), 
            .I3(n28606), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_736_7_lut (.I0(GND_net), .I1(n1005), .I2(VCC_net), 
            .I3(n28605), .O(n1070[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n28833), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28605), .I0(n1005), .I1(VCC_net), .CO(n28606));
    SB_CARRY mod_5_add_1808_19 (.CI(n28833), .I0(n2593), .I1(n2621), .CO(n28834));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n28832), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_6_lut (.I0(GND_net), .I1(n1006), .I2(VCC_net), 
            .I3(n28604), .O(n1070[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_6 (.CI(n28604), .I0(n1006), .I1(VCC_net), .CO(n28605));
    SB_CARRY mod_5_add_1808_18 (.CI(n28832), .I0(n2594), .I1(n2621), .CO(n28833));
    SB_LUT4 mod_5_add_736_5_lut (.I0(GND_net), .I1(n1007), .I2(VCC_net), 
            .I3(n28603), .O(n1070[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n28831), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28603), .I0(n1007), .I1(VCC_net), .CO(n28604));
    SB_LUT4 mod_5_add_736_4_lut (.I0(GND_net), .I1(n1008), .I2(VCC_net), 
            .I3(n28602), .O(n1070[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n28831), .I0(n2595), .I1(n2621), .CO(n28832));
    SB_CARRY mod_5_add_736_4 (.CI(n28602), .I0(n1008), .I1(VCC_net), .CO(n28603));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n28830), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_3_lut (.I0(GND_net), .I1(n1009), .I2(GND_net), 
            .I3(n28601), .O(n1070[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_5 (.CI(n27450), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27451));
    SB_CARRY mod_5_add_736_3 (.CI(n28601), .I0(n1009), .I1(GND_net), .CO(n28602));
    SB_CARRY mod_5_add_1808_16 (.CI(n28830), .I0(n2596), .I1(n2621), .CO(n28831));
    SB_LUT4 mod_5_add_736_2_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(VCC_net), .O(n1070[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(GND_net), 
            .CO(n28601));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n28829), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_7_lut (.I0(n41690), .I1(n905), .I2(VCC_net), 
            .I3(n28600), .O(n4_adj_3801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_15 (.CI(n28829), .I0(n2597), .I1(n2621), .CO(n28830));
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28599), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n28599), .I0(n906), .I1(VCC_net), .CO(n28600));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n34363), .I2(VCC_net), 
            .I3(n28598), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n28828), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n28828), .I0(n2598), .I1(n2621), .CO(n28829));
    SB_CARRY mod_5_add_669_5 (.CI(n28598), .I0(n34363), .I1(VCC_net), 
            .CO(n28599));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17645), .I2(VCC_net), 
            .I3(n28597), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n28597), .I0(n17645), .I1(VCC_net), 
            .CO(n28598));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n28827), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n28827), .I0(n2599), .I1(n2621), .CO(n28828));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n28826), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n15165), .I2(GND_net), 
            .I3(n28596), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n28596), .I0(n15165), .I1(GND_net), 
            .CO(n28597));
    SB_CARRY mod_5_add_1808_12 (.CI(n28826), .I0(n2600), .I1(n2621), .CO(n28827));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28596));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n28825), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n28825), .I0(n2601), .I1(n2621), .CO(n28826));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n28824), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_12_lut (.I0(n19), .I1(bit_ctr[10]), .I2(GND_net), .I3(n27457), 
            .O(n39081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_10 (.CI(n28824), .I0(n2602), .I1(n2621), .CO(n28825));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n28823), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n28823), .I0(n2603), .I1(n2621), .CO(n28824));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n28822), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n28822), .I0(n2604), .I1(n2621), .CO(n28823));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n28821), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n28821), .I0(n2605), .I1(n2621), .CO(n28822));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n28820), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n28820), .I0(n2606), .I1(n2621), .CO(n28821));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n28819), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n28819), .I0(n2607), .I1(n2621), .CO(n28820));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n28818), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n28818), .I0(n2608), .I1(n2621), .CO(n28819));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n41711), 
            .I3(n28817), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n28817), .I0(n2609), .I1(n41711), .CO(n28818));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n41711), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n41711), 
            .CO(n28817));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n28816), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n28815), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n28815), .I0(n2490), .I1(n2522), .CO(n28816));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n28814), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n28814), .I0(n2491), .I1(n2522), .CO(n28815));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n28813), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n28813), .I0(n2492), .I1(n2522), .CO(n28814));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n28812), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n27478), 
            .O(n39092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_19 (.CI(n28812), .I0(n2493), .I1(n2522), .CO(n28813));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n28811), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n28811), .I0(n2494), .I1(n2522), .CO(n28812));
    SB_LUT4 timer_1138_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28343), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1138_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28342), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_32 (.CI(n28342), .I0(GND_net), .I1(timer[30]), 
            .CO(n28343));
    SB_LUT4 timer_1138_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28341), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n28810), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_31 (.CI(n28341), .I0(GND_net), .I1(timer[29]), 
            .CO(n28342));
    SB_CARRY mod_5_add_1741_17 (.CI(n28810), .I0(n2495), .I1(n2522), .CO(n28811));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n28809), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28340), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n28809), .I0(n2496), .I1(n2522), .CO(n28810));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n28808), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_30 (.CI(n28340), .I0(GND_net), .I1(timer[28]), 
            .CO(n28341));
    SB_CARRY mod_5_add_1741_15 (.CI(n28808), .I0(n2497), .I1(n2522), .CO(n28809));
    SB_LUT4 timer_1138_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28339), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_29 (.CI(n28339), .I0(GND_net), .I1(timer[27]), 
            .CO(n28340));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n28807), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n28807), .I0(n2498), .I1(n2522), .CO(n28808));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n28806), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28338), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_28 (.CI(n28338), .I0(GND_net), .I1(timer[26]), 
            .CO(n28339));
    SB_LUT4 timer_1138_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28337), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_13 (.CI(n28806), .I0(n2499), .I1(n2522), .CO(n28807));
    SB_CARRY timer_1138_add_4_27 (.CI(n28337), .I0(GND_net), .I1(timer[25]), 
            .CO(n28338));
    SB_LUT4 timer_1138_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28336), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_26 (.CI(n28336), .I0(GND_net), .I1(timer[24]), 
            .CO(n28337));
    SB_LUT4 timer_1138_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28335), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n28805), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n28805), .I0(n2500), .I1(n2522), .CO(n28806));
    SB_CARRY timer_1138_add_4_25 (.CI(n28335), .I0(GND_net), .I1(timer[23]), 
            .CO(n28336));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n28804), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n28804), .I0(n2501), .I1(n2522), .CO(n28805));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n28803), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n27477), 
            .O(n39091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_10 (.CI(n28803), .I0(n2502), .I1(n2522), .CO(n28804));
    SB_LUT4 timer_1138_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28334), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n28802), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n28802), .I0(n2503), .I1(n2522), .CO(n28803));
    SB_CARRY timer_1138_add_4_24 (.CI(n28334), .I0(GND_net), .I1(timer[22]), 
            .CO(n28335));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n28801), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28333), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n28801), .I0(n2504), .I1(n2522), .CO(n28802));
    SB_CARRY timer_1138_add_4_23 (.CI(n28333), .I0(GND_net), .I1(timer[21]), 
            .CO(n28334));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n28800), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28332), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n28800), .I0(n2505), .I1(n2522), .CO(n28801));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n28799), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n28799), .I0(n2506), .I1(n2522), .CO(n28800));
    SB_CARRY timer_1138_add_4_22 (.CI(n28332), .I0(GND_net), .I1(timer[20]), 
            .CO(n28333));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n28798), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28331), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_21 (.CI(n28331), .I0(GND_net), .I1(timer[19]), 
            .CO(n28332));
    SB_CARRY add_21_32 (.CI(n27477), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27478));
    SB_LUT4 add_21_31_lut (.I0(n19), .I1(bit_ctr[29]), .I2(GND_net), .I3(n27476), 
            .O(n39090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i140_4_lut (.I0(n165), .I1(n136), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n166));   // verilog/neopixel.v(16[20:25])
    defparam i140_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i30899_4_lut (.I0(\state[1] ), .I1(start), .I2(n166), .I3(n168), 
            .O(n37153));   // verilog/neopixel.v(16[20:25])
    defparam i30899_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mod_5_add_1741_5 (.CI(n28798), .I0(n2507), .I1(n2522), .CO(n28799));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n28797), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28330), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_20 (.CI(n28330), .I0(GND_net), .I1(timer[18]), 
            .CO(n28331));
    SB_LUT4 timer_1138_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28329), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n27476), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27477));
    SB_CARRY mod_5_add_1741_4 (.CI(n28797), .I0(n2508), .I1(n2522), .CO(n28798));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n41712), 
            .I3(n28796), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1138_add_4_19 (.CI(n28329), .I0(GND_net), .I1(timer[17]), 
            .CO(n28330));
    SB_LUT4 timer_1138_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28328), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n28796), .I0(n2509), .I1(n41712), .CO(n28797));
    SB_CARRY timer_1138_add_4_18 (.CI(n28328), .I0(GND_net), .I1(timer[16]), 
            .CO(n28329));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n41712), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1138_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28327), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_30_lut (.I0(n19), .I1(bit_ctr[28]), .I2(GND_net), .I3(n27475), 
            .O(n39089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n41712), 
            .CO(n28796));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n28795), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_17 (.CI(n28327), .I0(GND_net), .I1(timer[15]), 
            .CO(n28328));
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n28794), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28326), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n28794), .I0(n2391), .I1(n2423), .CO(n28795));
    SB_CARRY add_21_30 (.CI(n27475), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27476));
    SB_LUT4 add_21_29_lut (.I0(n19), .I1(bit_ctr[27]), .I2(GND_net), .I3(n27474), 
            .O(n39088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n32712));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n28793), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_16 (.CI(n28326), .I0(GND_net), .I1(timer[14]), 
            .CO(n28327));
    SB_LUT4 timer_1138_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28325), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_15 (.CI(n28325), .I0(GND_net), .I1(timer[13]), 
            .CO(n28326));
    SB_CARRY mod_5_add_1674_20 (.CI(n28793), .I0(n2392), .I1(n2423), .CO(n28794));
    SB_LUT4 timer_1138_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28324), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(n2406), .I1(n2402), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_3803));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1387 (.I0(n2395), .I1(n2408), .I2(n2394), .I3(n2399), 
            .O(n32_adj_3804));
    defparam i12_4_lut_adj_1387.LUT_INIT = 16'hfffe;
    SB_LUT4 i20790_2_lut (.I0(bit_ctr[11]), .I1(n2409), .I2(GND_net), 
            .I3(GND_net), .O(n25276));
    defparam i20790_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16_4_lut (.I0(n2404), .I1(n32_adj_3804), .I2(n22_adj_3803), 
            .I3(n2393), .O(n36));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n18052));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n18051));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n18050));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n18049));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n18048));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n18047));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n18046));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n18045));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n18044));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n18043));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1138__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n18042));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n18041));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_12 (.CI(n27457), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27458));
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n18040));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i14_4_lut_adj_1388 (.I0(n2407), .I1(n2398), .I2(n2401), .I3(n2405), 
            .O(n34_adj_3806));
    defparam i14_4_lut_adj_1388.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n18039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n18038));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n18037));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n18036));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n28792), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n18035));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_29 (.CI(n27474), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27475));
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n18034));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n18033));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i15_4_lut_adj_1389 (.I0(n2397), .I1(n2392), .I2(n25276), .I3(n2391), 
            .O(n35));
    defparam i15_4_lut_adj_1389.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n18032));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n18031));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n18030));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i13_4_lut_adj_1390 (.I0(n2390), .I1(n2403), .I2(n2396), .I3(n2400), 
            .O(n33_adj_3807));
    defparam i13_4_lut_adj_1390.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n33_adj_3807), .I1(n35), .I2(n34_adj_3806), 
            .I3(n36), .O(n2423));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1138_add_4_14 (.CI(n28324), .I0(GND_net), .I1(timer[12]), 
            .CO(n28325));
    SB_CARRY mod_5_add_1674_19 (.CI(n28792), .I0(n2393), .I1(n2423), .CO(n28793));
    SB_LUT4 timer_1138_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28323), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n18029));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n18028));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n18027));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n18026));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n18025));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n18024));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n18023));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1138_add_4_13 (.CI(n28323), .I0(GND_net), .I1(timer[11]), 
            .CO(n28324));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n28791), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n32710));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n32708));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i35392_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41712));
    defparam i35392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1138_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28322), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_18 (.CI(n28791), .I0(n2394), .I1(n2423), .CO(n28792));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n28790), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(n19), .I1(bit_ctr[9]), .I2(GND_net), .I3(n27456), 
            .O(n39080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_28_lut (.I0(n19), .I1(bit_ctr[26]), .I2(GND_net), .I3(n27473), 
            .O(n39087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_17 (.CI(n28790), .I0(n2395), .I1(n2423), .CO(n28791));
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n27449), 
            .O(n39094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n28789), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_12 (.CI(n28322), .I0(GND_net), .I1(timer[10]), 
            .CO(n28323));
    SB_CARRY mod_5_add_1674_16 (.CI(n28789), .I0(n2396), .I1(n2423), .CO(n28790));
    SB_LUT4 timer_1138_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28321), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n32702));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n32700));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n28788), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n28788), .I0(n2397), .I1(n2423), .CO(n28789));
    SB_CARRY timer_1138_add_4_11 (.CI(n28321), .I0(GND_net), .I1(timer[9]), 
            .CO(n28322));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n28787), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n28787), .I0(n2398), .I1(n2423), .CO(n28788));
    SB_CARRY add_21_11 (.CI(n27456), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27457));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n28786), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(VCC_net), 
            .D(n32694));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_1138_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28320), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n28786), .I0(n2399), .I1(n2423), .CO(n28787));
    SB_CARRY timer_1138_add_4_10 (.CI(n28320), .I0(GND_net), .I1(timer[8]), 
            .CO(n28321));
    SB_LUT4 timer_1138_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28319), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n28785), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n28785), .I0(n2400), .I1(n2423), .CO(n28786));
    SB_CARRY timer_1138_add_4_9 (.CI(n28319), .I0(GND_net), .I1(timer[7]), 
            .CO(n28320));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n28784), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28318), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n28784), .I0(n2401), .I1(n2423), .CO(n28785));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n28783), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_28 (.CI(n27473), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27474));
    SB_CARRY mod_5_add_1674_10 (.CI(n28783), .I0(n2402), .I1(n2423), .CO(n28784));
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n32698));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n28782), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n28782), .I0(n2403), .I1(n2423), .CO(n28783));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n28781), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n28781), .I0(n2404), .I1(n2423), .CO(n28782));
    SB_CARRY timer_1138_add_4_8 (.CI(n28318), .I0(GND_net), .I1(timer[6]), 
            .CO(n28319));
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n32696));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n28780), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1138_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28317), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n27449), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27450));
    SB_CARRY timer_1138_add_4_7 (.CI(n28317), .I0(GND_net), .I1(timer[5]), 
            .CO(n28318));
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n18000));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n32692));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_7 (.CI(n28780), .I0(n2405), .I1(n2423), .CO(n28781));
    SB_LUT4 timer_1138_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28316), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1138_add_4_6 (.CI(n28316), .I0(GND_net), .I1(timer[4]), 
            .CO(n28317));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n28779), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n28779), .I0(n2406), .I1(n2423), .CO(n28780));
    SB_LUT4 timer_1138_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28315), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n28778), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1138_add_4_5 (.CI(n28315), .I0(GND_net), .I1(timer[3]), 
            .CO(n28316));
    SB_LUT4 add_21_10_lut (.I0(n19), .I1(bit_ctr[8]), .I2(GND_net), .I3(n27455), 
            .O(n39079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 timer_1138_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28314), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_27_lut (.I0(n19), .I1(bit_ctr[25]), .I2(GND_net), .I3(n27472), 
            .O(n39086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_5 (.CI(n28778), .I0(n2407), .I1(n2423), .CO(n28779));
    SB_LUT4 i20978_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n25466));
    defparam i20978_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1391 (.I0(n1405), .I1(n25466), .I2(n1403), .I3(n1406), 
            .O(n16_adj_3809));
    defparam i6_4_lut_adj_1391.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1392 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_3810));
    defparam i7_4_lut_adj_1392.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1393 (.I0(n17_adj_3810), .I1(n1408), .I2(n16_adj_3809), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1393.LUT_INIT = 16'hfffe;
    SB_LUT4 i35383_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41703));
    defparam i35383_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1138_add_4_4 (.CI(n28314), .I0(GND_net), .I1(timer[2]), 
            .CO(n28315));
    SB_LUT4 timer_1138_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28313), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n28777), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_3_lut (.I0(n19), .I1(bit_ctr[1]), .I2(GND_net), .I3(n27448), 
            .O(n39093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_10 (.CI(n27455), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27456));
    SB_CARRY timer_1138_add_4_3 (.CI(n28313), .I0(GND_net), .I1(timer[1]), 
            .CO(n28314));
    SB_CARRY add_21_27 (.CI(n27472), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27473));
    SB_LUT4 timer_1138_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1138_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_26_lut (.I0(n19), .I1(bit_ctr[24]), .I2(GND_net), .I3(n27471), 
            .O(n39085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_4 (.CI(n28777), .I0(n2408), .I1(n2423), .CO(n28778));
    SB_CARRY add_21_26 (.CI(n27471), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27472));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n41714), 
            .I3(n28776), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n28776), .I0(n2409), .I1(n41714), .CO(n28777));
    SB_CARRY timer_1138_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28313));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n41714), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n27454), 
            .O(n39070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n41714), 
            .CO(n28776));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n28775), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n28774), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n32690));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1607_20 (.CI(n28774), .I0(n2292), .I1(n2324), .CO(n28775));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17922));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n28773), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n28773), .I0(n2293), .I1(n2324), .CO(n28774));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n28772), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut_adj_1394 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_3811));
    defparam i3_2_lut_adj_1394.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1395 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_3812));
    defparam i13_4_lut_adj_1395.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), .I3(GND_net), 
            .O(n22_adj_3813));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut (.I0(n2490), .I1(n34_adj_3812), .I2(n24_adj_3811), 
            .I3(n2494), .O(n38));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1396 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_3814));
    defparam i15_4_lut_adj_1396.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1397 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_3813), 
            .O(n37));
    defparam i16_4_lut_adj_1397.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1398 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_3815));
    defparam i14_4_lut_adj_1398.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35_adj_3815), .I1(n37), .I2(n36_adj_3814), 
            .I3(n38), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35391_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41711));
    defparam i35391_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35368_1_lut (.I0(n30590), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41690));   // verilog/neopixel.v(22[26:36])
    defparam i35368_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35390_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41710));
    defparam i35390_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1399 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_3816));
    defparam i14_4_lut_adj_1399.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_3817));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1400 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_3818));
    defparam i12_4_lut_adj_1400.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1401 (.I0(n25_adj_3817), .I1(n36_adj_3816), .I2(n2594), 
            .I3(n2589), .O(n40));
    defparam i18_4_lut_adj_1401.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1402 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_3819));
    defparam i16_4_lut_adj_1402.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_3818), .I2(n2603), .I3(GND_net), 
            .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1403 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_3820));
    defparam i15_4_lut_adj_1403.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37_adj_3820), .I1(n39), .I2(n38_adj_3819), 
            .I3(n40), .O(n2621));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35386_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41706));
    defparam i35386_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_25_lut (.I0(n19), .I1(bit_ctr[23]), .I2(GND_net), .I3(n27470), 
            .O(n39084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1607_18 (.CI(n28772), .I0(n2294), .I1(n2324), .CO(n28773));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n28771), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i742_3_lut (.I0(n1008), .I1(n1070[27]), .I2(n1037), 
            .I3(GND_net), .O(n1107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35373_2_lut (.I0(n30590), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i35373_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i35375_2_lut (.I0(n30590), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i35375_2_lut.LUT_INIT = 16'h4444;
    SB_CARRY mod_5_add_1607_17 (.CI(n28771), .I0(n2295), .I1(n2324), .CO(n28772));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n28770), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n28770), .I0(n2296), .I1(n2324), .CO(n28771));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n28769), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n28769), .I0(n2297), .I1(n2324), .CO(n28770));
    SB_LUT4 mod_5_i675_3_lut (.I0(n15165), .I1(n971[27]), .I2(n30590), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n15165));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n28768), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n28768), .I0(n2298), .I1(n2324), .CO(n28769));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n28767), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n28767), .I0(n2299), .I1(n2324), .CO(n28768));
    SB_CARRY add_21_9 (.CI(n27454), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27455));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n28766), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n28766), .I0(n2300), .I1(n2324), .CO(n28767));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n28765), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n28765), .I0(n2301), .I1(n2324), .CO(n28766));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n28764), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n28764), .I0(n2302), .I1(n2324), .CO(n28765));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n28763), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n28763), .I0(n2303), .I1(n2324), .CO(n28764));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n28762), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n28762), .I0(n2304), .I1(n2324), .CO(n28763));
    SB_CARRY add_21_25 (.CI(n27470), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27471));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n28761), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n28761), .I0(n2305), .I1(n2324), .CO(n28762));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n28760), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n28760), .I0(n2306), .I1(n2324), .CO(n28761));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n28759), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n28759), .I0(n2307), .I1(n2324), .CO(n28760));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n28758), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n28758), .I0(n2308), .I1(n2324), .CO(n28759));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n41715), 
            .I3(n28757), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n28757), .I0(n2309), .I1(n41715), .CO(n28758));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n41715), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n41715), 
            .CO(n28757));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n28756), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n28755), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n28755), .I0(n2193), .I1(n2225), .CO(n28756));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n28754), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n28754), .I0(n2194), .I1(n2225), .CO(n28755));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n28753), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n28753), .I0(n2195), .I1(n2225), .CO(n28754));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n28752), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i33333_3_lut_4_lut (.I0(n62), .I1(bit_ctr[28]), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17645));
    defparam i33333_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_CARRY mod_5_add_1540_16 (.CI(n28752), .I0(n2196), .I1(n2225), .CO(n28753));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n28751), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY mod_5_add_1540_15 (.CI(n28751), .I0(n2197), .I1(n2225), .CO(n28752));
    SB_LUT4 i3_3_lut_adj_1405 (.I0(n34363), .I1(n906), .I2(n17645), .I3(GND_net), 
            .O(n8));   // verilog/neopixel.v(22[26:36])
    defparam i3_3_lut_adj_1405.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut (.I0(n905), .I1(n8), .I2(bit_ctr[26]), .I3(n15165), 
            .O(n30590));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h0444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n30590), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28269_3_lut (.I0(n30590), .I1(n971[28]), .I2(n971[29]), .I3(GND_net), 
            .O(n34512));
    defparam i28269_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 i2_3_lut (.I0(n1005), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n7));   // verilog/neopixel.v(22[26:36])
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i4_4_lut_adj_1406 (.I0(n7), .I1(n34512), .I2(n4_adj_3801), 
            .I3(n1008), .O(n1037));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut_adj_1406.LUT_INIT = 16'hfffb;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n30590), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i743_3_lut (.I0(n1009), .I1(n1070[26]), .I2(n1037), 
            .I3(GND_net), .O(n1108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i741_3_lut (.I0(n1007), .I1(n1070[28]), .I2(n1037), 
            .I3(GND_net), .O(n1106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i739_3_lut (.I0(n1005), .I1(n1070[30]), .I2(n1037), 
            .I3(GND_net), .O(n1104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i740_3_lut (.I0(n1006), .I1(n1070[29]), .I2(n1037), 
            .I3(GND_net), .O(n1105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i744_3_lut (.I0(bit_ctr[25]), .I1(n1070[25]), .I2(n1037), 
            .I3(GND_net), .O(n1109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21013_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n25502));
    defparam i21013_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1104), .I2(n1106), .I3(n1108), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1407 (.I0(n1107), .I1(n12), .I2(n1103), .I3(n25502), 
            .O(n1136));
    defparam i6_4_lut_adj_1407.LUT_INIT = 16'hfffe;
    SB_LUT4 i35389_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41709));
    defparam i35389_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n28750), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n28750), .I0(n2198), .I1(n2225), .CO(n28751));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n28749), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n28749), .I0(n2199), .I1(n2225), .CO(n28750));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n28748), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n28748), .I0(n2200), .I1(n2225), .CO(n28749));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n28747), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n27469), 
            .O(n39083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1540_11 (.CI(n28747), .I0(n2201), .I1(n2225), .CO(n28748));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n28746), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n27448), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27449));
    SB_CARRY mod_5_add_1540_10 (.CI(n28746), .I0(n2202), .I1(n2225), .CO(n28747));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n28745), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n28745), .I0(n2203), .I1(n2225), .CO(n28746));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n28744), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1408 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1208), 
            .O(n14));
    defparam i6_4_lut_adj_1408.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1409 (.I0(bit_ctr[23]), .I1(n1202), .I2(n1209), 
            .I3(GND_net), .O(n9));
    defparam i1_3_lut_adj_1409.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1410 (.I0(n9), .I1(n14), .I2(n1203), .I3(n1207), 
            .O(n1235));
    defparam i7_4_lut_adj_1410.LUT_INIT = 16'hfffe;
    SB_LUT4 i35387_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41707));
    defparam i35387_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1411 (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_3821));
    defparam i2_2_lut_adj_1411.LUT_INIT = 16'heeee;
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n27453), 
            .O(n39069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1540_8 (.CI(n28744), .I0(n2204), .I1(n2225), .CO(n28745));
    SB_LUT4 i20_4_lut_adj_1412 (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut_adj_1412.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1413 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut_adj_1413.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1414 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut_adj_1414.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1415 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut_adj_1415.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1416 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut_adj_1416.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n28743), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1417 (.I0(bit_ctr[3]), .I1(n30_adj_3821), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut_adj_1417.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_7 (.CI(n28743), .I0(n2205), .I1(n2225), .CO(n28744));
    SB_LUT4 i21_4_lut_adj_1418 (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut_adj_1418.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n28742), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4021_2_lut_3_lut_4_lut (.I0(n62), .I1(bit_ctr[28]), .I2(bit_ctr[27]), 
            .I3(n34361), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i4021_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_CARRY add_21_24 (.CI(n27469), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27470));
    SB_CARRY mod_5_add_1540_6 (.CI(n28742), .I0(n2206), .I1(n2225), .CO(n28743));
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_337[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n28741), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n28741), .I0(n2207), .I1(n2225), .CO(n28742));
    SB_LUT4 i2026_4_lut (.I0(n37149), .I1(\state_3__N_337[1] ), .I2(\state[1] ), 
            .I3(start), .O(n4488));
    defparam i2026_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i12_4_lut_adj_1419 (.I0(\state[1] ), .I1(n4488), .I2(\state[0] ), 
            .I3(n131), .O(n17536));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_4_lut_adj_1419.LUT_INIT = 16'h3530;
    SB_LUT4 i16_4_lut_adj_1420 (.I0(n2786), .I1(n2792), .I2(n2791), .I3(n2794), 
            .O(n40_adj_3822));
    defparam i16_4_lut_adj_1420.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n28740), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n28740), .I0(n2208), .I1(n2225), .CO(n28741));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n41716), 
            .I3(n28739), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n28739), .I0(n2209), .I1(n41716), .CO(n28740));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n41716), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n41716), 
            .CO(n28739));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n28738), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n28737), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n28737), .I0(n2094), .I1(n2126), .CO(n28738));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n28736), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n28736), .I0(n2095), .I1(n2126), .CO(n28737));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n28735), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n28735), .I0(n2096), .I1(n2126), .CO(n28736));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n28734), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n28734), .I0(n2097), .I1(n2126), .CO(n28735));
    SB_LUT4 add_21_23_lut (.I0(n19), .I1(bit_ctr[21]), .I2(GND_net), .I3(n27468), 
            .O(n39082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n28733), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n28733), .I0(n2098), .I1(n2126), .CO(n28734));
    SB_LUT4 i5_3_lut (.I0(n1308), .I1(n1304), .I2(n1305), .I3(GND_net), 
            .O(n14_adj_3823));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut_adj_1421 (.I0(n1301), .I1(n1302), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_3824));
    defparam i3_2_lut_adj_1421.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1422 (.I0(n1306), .I1(n14_adj_3823), .I2(bit_ctr[22]), 
            .I3(n1309), .O(n16_adj_3825));
    defparam i7_4_lut_adj_1422.LUT_INIT = 16'hfeee;
    SB_LUT4 i8_4_lut (.I0(n1307), .I1(n16_adj_3825), .I2(n12_adj_3824), 
            .I3(n1303), .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_3826));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1423 (.I0(one_wire_N_488[2]), .I1(one_wire_N_488[4]), 
            .I2(one_wire_N_488[3]), .I3(GND_net), .O(n136));   // verilog/neopixel.v(53[15:25])
    defparam i2_3_lut_adj_1423.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_adj_1424 (.I0(one_wire_N_488[4]), .I1(n35812), .I2(one_wire_N_488[3]), 
            .I3(GND_net), .O(n165));   // verilog/neopixel.v(6[16:24])
    defparam i1_3_lut_adj_1424.LUT_INIT = 16'heaea;
    SB_LUT4 i7_4_lut_adj_1425 (.I0(n9_adj_3827), .I1(n11), .I2(n10), .I3(n24843), 
            .O(n168));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1425.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1426 (.I0(n168), .I1(n165), .I2(GND_net), .I3(GND_net), 
            .O(n21));   // verilog/neopixel.v(6[16:24])
    defparam i2_2_lut_adj_1426.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(n136), .I1(n168), .I2(GND_net), .I3(GND_net), 
            .O(n19765));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1428 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_3829));
    defparam i15_4_lut_adj_1428.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n28732), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n28732), .I0(n2099), .I1(n2126), .CO(n28733));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n28731), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n28731), .I0(n2100), .I1(n2126), .CO(n28732));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n28730), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n28730), .I0(n2101), .I1(n2126), .CO(n28731));
    SB_LUT4 i20772_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n25258));
    defparam i20772_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n28729), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n28729), .I0(n2102), .I1(n2126), .CO(n28730));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n28728), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n28728), .I0(n2103), .I1(n2126), .CO(n28729));
    SB_LUT4 i13_4_lut_adj_1429 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n25258), 
            .O(n36_adj_3830));
    defparam i13_4_lut_adj_1429.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n28963), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n28727), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n28962), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n28962), .I0(n3084), .I1(n3116), .CO(n28963));
    SB_CARRY mod_5_add_1473_8 (.CI(n28727), .I0(n2104), .I1(n2126), .CO(n28728));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n28726), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n28961), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n28726), .I0(n2105), .I1(n2126), .CO(n28727));
    SB_CARRY mod_5_add_2143_27 (.CI(n28961), .I0(n3085), .I1(n3116), .CO(n28962));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n28725), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n28960), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n28725), .I0(n2106), .I1(n2126), .CO(n28726));
    SB_CARRY mod_5_add_2143_26 (.CI(n28960), .I0(n3086), .I1(n3116), .CO(n28961));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n28959), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut (.I0(n19765), .I1(n21), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n26_adj_3831));
    defparam i1_4_lut.LUT_INIT = 16'h3553;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n28724), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1138__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1138__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17792));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17561), .D(state_3__N_337[0]), 
            .S(n17721));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_5 (.CI(n28724), .I0(n2107), .I1(n2126), .CO(n28725));
    SB_CARRY mod_5_add_2143_25 (.CI(n28959), .I0(n3087), .I1(n3116), .CO(n28960));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n28723), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n28958), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n28723), .I0(n2108), .I1(n2126), .CO(n28724));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n41717), 
            .I3(n28722), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n28722), .I0(n2109), .I1(n41717), .CO(n28723));
    SB_CARRY mod_5_add_2143_24 (.CI(n28958), .I0(n3088), .I1(n3116), .CO(n28959));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n28957), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n41717), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n41717), 
            .CO(n28722));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n28721), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n28957), .I0(n3089), .I1(n3116), .CO(n28958));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n28720), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n28956), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n28720), .I0(n1995), .I1(n2027), .CO(n28721));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n28719), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n28956), .I0(n3090), .I1(n3116), .CO(n28957));
    SB_CARRY mod_5_add_1406_16 (.CI(n28719), .I0(n1996), .I1(n2027), .CO(n28720));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n28955), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n28718), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n28955), .I0(n3091), .I1(n3116), .CO(n28956));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n28954), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n28718), .I0(n1997), .I1(n2027), .CO(n28719));
    SB_LUT4 i15316_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_545 ));   // verilog/neopixel.v(16[20:25])
    defparam i15316_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY mod_5_add_2143_20 (.CI(n28954), .I0(n3092), .I1(n3116), .CO(n28955));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n28953), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n28717), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_23 (.CI(n27468), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27469));
    SB_CARRY mod_5_add_2143_19 (.CI(n28953), .I0(n3093), .I1(n3116), .CO(n28954));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n28952), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_22_lut (.I0(n19), .I1(bit_ctr[20]), .I2(GND_net), .I3(n27467), 
            .O(n39078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2143_18 (.CI(n28952), .I0(n3094), .I1(n3116), .CO(n28953));
    SB_CARRY mod_5_add_1406_14 (.CI(n28717), .I0(n1998), .I1(n2027), .CO(n28718));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n28951), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n28716), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n28951), .I0(n3095), .I1(n3116), .CO(n28952));
    SB_CARRY mod_5_add_1406_13 (.CI(n28716), .I0(n1999), .I1(n2027), .CO(n28717));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n28950), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n28950), .I0(n3096), .I1(n3116), .CO(n28951));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n28715), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n28715), .I0(n2000), .I1(n2027), .CO(n28716));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n28949), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n28714), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n28949), .I0(n3097), .I1(n3116), .CO(n28950));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n28948), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n28714), .I0(n2001), .I1(n2027), .CO(n28715));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n28713), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n28948), .I0(n3098), .I1(n3116), .CO(n28949));
    SB_CARRY add_21_22 (.CI(n27467), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27468));
    SB_CARRY mod_5_add_1406_10 (.CI(n28713), .I0(n2002), .I1(n2027), .CO(n28714));
    SB_LUT4 add_21_21_lut (.I0(n19), .I1(bit_ctr[19]), .I2(GND_net), .I3(n27466), 
            .O(n39077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i19_4_lut_adj_1430 (.I0(n2700), .I1(n38_adj_3829), .I2(n28_adj_3826), 
            .I3(n2705), .O(n42));
    defparam i19_4_lut_adj_1430.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n28947), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_4_lut_adj_1431 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_3832));
    defparam i17_4_lut_adj_1431.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n28712), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n28712), .I0(n2003), .I1(n2027), .CO(n28713));
    SB_CARRY mod_5_add_2143_13 (.CI(n28947), .I0(n3099), .I1(n3116), .CO(n28948));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n28946), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n28711), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n28711), .I0(n2004), .I1(n2027), .CO(n28712));
    SB_CARRY add_21_21 (.CI(n27466), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27467));
    SB_CARRY mod_5_add_2143_12 (.CI(n28946), .I0(n3100), .I1(n3116), .CO(n28947));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n28710), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n28710), .I0(n2005), .I1(n2027), .CO(n28711));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n28945), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n28709), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n28945), .I0(n3101), .I1(n3116), .CO(n28946));
    SB_CARRY mod_5_add_1406_6 (.CI(n28709), .I0(n2006), .I1(n2027), .CO(n28710));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n28944), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n28708), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n28944), .I0(n3102), .I1(n3116), .CO(n28945));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n28943), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n28943), .I0(n3103), .I1(n3116), .CO(n28944));
    SB_CARRY mod_5_add_1406_5 (.CI(n28708), .I0(n2007), .I1(n2027), .CO(n28709));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n28942), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n28707), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n28942), .I0(n3104), .I1(n3116), .CO(n28943));
    SB_CARRY mod_5_add_1406_4 (.CI(n28707), .I0(n2008), .I1(n2027), .CO(n28708));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n28941), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n41720), 
            .I3(n28706), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_7 (.CI(n28941), .I0(n3105), .I1(n3116), .CO(n28942));
    SB_CARRY mod_5_add_1406_3 (.CI(n28706), .I0(n2009), .I1(n41720), .CO(n28707));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n28940), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n41720), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_6 (.CI(n28940), .I0(n3106), .I1(n3116), .CO(n28941));
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n41720), 
            .CO(n28706));
    SB_LUT4 i18_4_lut_adj_1432 (.I0(n2687), .I1(n36_adj_3830), .I2(n2703), 
            .I3(n2695), .O(n41));
    defparam i18_4_lut_adj_1432.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n28939), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n28705), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n28939), .I0(n3107), .I1(n3116), .CO(n28940));
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n28704), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n28938), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n28704), .I0(n1896), .I1(n1928), .CO(n28705));
    SB_CARRY mod_5_add_2143_4 (.CI(n28938), .I0(n3108), .I1(n3116), .CO(n28939));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n41719), 
            .I3(n28937), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n28703), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_3 (.CI(n28937), .I0(n3109), .I1(n41719), .CO(n28938));
    SB_CARRY mod_5_add_1339_15 (.CI(n28703), .I0(n1897), .I1(n1928), .CO(n28704));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n41719), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n28702), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n41719), 
            .CO(n28937));
    SB_CARRY mod_5_add_1339_14 (.CI(n28702), .I0(n1898), .I1(n1928), .CO(n28703));
    SB_LUT4 i16_4_lut_adj_1433 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_3833));
    defparam i16_4_lut_adj_1433.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n28936), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n27465), 
            .O(n39072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n28701), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n27465), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27466));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n28935), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n28701), .I0(n1899), .I1(n1928), .CO(n28702));
    SB_CARRY mod_5_add_2076_27 (.CI(n28935), .I0(n2985), .I1(n3017), .CO(n28936));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n28700), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_19_lut (.I0(n19), .I1(bit_ctr[17]), .I2(GND_net), .I3(n27464), 
            .O(n39071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14_4_lut_adj_1434 (.I0(n2790), .I1(n2807), .I2(n2788), .I3(n2796), 
            .O(n38_adj_3834));
    defparam i14_4_lut_adj_1434.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n28934), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n28700), .I0(n1900), .I1(n1928), .CO(n28701));
    SB_CARRY mod_5_add_2076_26 (.CI(n28934), .I0(n2986), .I1(n3017), .CO(n28935));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n28933), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n28699), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n28933), .I0(n2987), .I1(n3017), .CO(n28934));
    SB_CARRY mod_5_add_1339_11 (.CI(n28699), .I0(n1901), .I1(n1928), .CO(n28700));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n28698), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n28932), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n28698), .I0(n1902), .I1(n1928), .CO(n28699));
    SB_CARRY mod_5_add_2076_24 (.CI(n28932), .I0(n2988), .I1(n3017), .CO(n28933));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n28697), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n28931), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n28697), .I0(n1903), .I1(n1928), .CO(n28698));
    SB_CARRY mod_5_add_2076_23 (.CI(n28931), .I0(n2989), .I1(n3017), .CO(n28932));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n28696), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n28930), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n28696), .I0(n1904), .I1(n1928), .CO(n28697));
    SB_CARRY mod_5_add_2076_22 (.CI(n28930), .I0(n2990), .I1(n3017), .CO(n28931));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n28929), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n28929), .I0(n2991), .I1(n3017), .CO(n28930));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n28695), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n28695), .I0(n1905), .I1(n1928), .CO(n28696));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n28928), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n28928), .I0(n2992), .I1(n3017), .CO(n28929));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n28694), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n28927), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n28694), .I0(n1906), .I1(n1928), .CO(n28695));
    SB_CARRY mod_5_add_2076_19 (.CI(n28927), .I0(n2993), .I1(n3017), .CO(n28928));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n28926), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n28693), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n28926), .I0(n2994), .I1(n3017), .CO(n28927));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n28925), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n28693), .I0(n1907), .I1(n1928), .CO(n28694));
    SB_CARRY mod_5_add_2076_17 (.CI(n28925), .I0(n2995), .I1(n3017), .CO(n28926));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n28692), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n28692), .I0(n1908), .I1(n1928), .CO(n28693));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n41721), 
            .I3(n28691), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i30989_3_lut (.I0(\color[16] ), .I1(\color[17] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n37309));
    defparam i30989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_4_lut (.I0(n39_adj_3833), .I1(n41), .I2(n40_adj_3832), 
            .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n28924), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n28924), .I0(n2996), .I1(n3017), .CO(n28925));
    SB_LUT4 i30990_3_lut (.I0(\color[18] ), .I1(\color[19] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n37310));
    defparam i30990_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1339_3 (.CI(n28691), .I0(n1909), .I1(n41721), .CO(n28692));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n41721), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i31047_3_lut (.I0(\color[22] ), .I1(\color[23] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n37367));
    defparam i31047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n28923), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n41721), 
            .CO(n28691));
    SB_CARRY mod_5_add_2076_15 (.CI(n28923), .I0(n2997), .I1(n3017), .CO(n28924));
    SB_LUT4 i31046_3_lut (.I0(\color[20] ), .I1(\color[21] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n37366));
    defparam i31046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n28922), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n28690), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n28922), .I0(n2998), .I1(n3017), .CO(n28923));
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n28689), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n28921), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n28689), .I0(n1797), .I1(n1829), .CO(n28690));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_13 (.CI(n28921), .I0(n2999), .I1(n3017), .CO(n28922));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n28688), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1435 (.I0(n2797), .I1(n2799), .I2(n2793), .I3(n2803), 
            .O(n39_adj_3840));
    defparam i15_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n28920), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n28688), .I0(n1798), .I1(n1829), .CO(n28689));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_12 (.CI(n28920), .I0(n3000), .I1(n3017), .CO(n28921));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n28687), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n28687), .I0(n1799), .I1(n1829), .CO(n28688));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n28919), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n28686), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1272_12 (.CI(n28686), .I0(n1800), .I1(n1829), .CO(n28687));
    SB_CARRY mod_5_add_2076_11 (.CI(n28919), .I0(n3001), .I1(n3017), .CO(n28920));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n28685), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n28685), .I0(n1801), .I1(n1829), .CO(n28686));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n28918), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n28684), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n28918), .I0(n3002), .I1(n3017), .CO(n28919));
    SB_CARRY mod_5_add_1272_10 (.CI(n28684), .I0(n1802), .I1(n1829), .CO(n28685));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n28917), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n28683), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n28917), .I0(n3003), .I1(n3017), .CO(n28918));
    SB_CARRY mod_5_add_1272_9 (.CI(n28683), .I0(n1803), .I1(n1829), .CO(n28684));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n28916), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n27453), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27454));
    SB_CARRY add_21_19 (.CI(n27464), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27465));
    SB_LUT4 add_21_18_lut (.I0(n19), .I1(bit_ctr[16]), .I2(GND_net), .I3(n27463), 
            .O(n39067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_8 (.CI(n28916), .I0(n3004), .I1(n3017), .CO(n28917));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n28682), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n28915), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n28682), .I0(n1804), .I1(n1829), .CO(n28683));
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n28681), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n28915), .I0(n3005), .I1(n3017), .CO(n28916));
    SB_CARRY mod_5_add_1272_7 (.CI(n28681), .I0(n1805), .I1(n1829), .CO(n28682));
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n28914), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n28680), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n28914), .I0(n3006), .I1(n3017), .CO(n28915));
    SB_CARRY mod_5_add_1272_6 (.CI(n28680), .I0(n1806), .I1(n1829), .CO(n28681));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n28913), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n28913), .I0(n3007), .I1(n3017), .CO(n28914));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n28679), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n28679), .I0(n1807), .I1(n1829), .CO(n28680));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n28912), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n28678), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n28912), .I0(n3008), .I1(n3017), .CO(n28913));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n41722), 
            .I3(n28911), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_4 (.CI(n28678), .I0(n1808), .I1(n1829), .CO(n28679));
    SB_CARRY mod_5_add_2076_3 (.CI(n28911), .I0(n3009), .I1(n41722), .CO(n28912));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n41723), 
            .I3(n28677), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i35406_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41726));
    defparam i35406_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n41722), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n28677), .I0(n1809), .I1(n41723), .CO(n28678));
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n41723), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n41722), 
            .CO(n28911));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n41723), 
            .CO(n28677));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n28910), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n28676), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n28909), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_26 (.CI(n28909), .I0(n2886), .I1(n2918), .CO(n28910));
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n28675), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_14 (.CI(n28675), .I0(n1698), .I1(n1730), .CO(n28676));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n28674), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_18 (.CI(n27463), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27464));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n28908), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_13 (.CI(n28674), .I0(n1699), .I1(n1730), .CO(n28675));
    SB_LUT4 i35404_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41724));
    defparam i35404_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n28673), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_25 (.CI(n28908), .I0(n2887), .I1(n2918), .CO(n28909));
    SB_CARRY mod_5_add_1205_12 (.CI(n28673), .I0(n1700), .I1(n1730), .CO(n28674));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n28907), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n28672), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n28907), .I0(n2888), .I1(n2918), .CO(n28908));
    SB_LUT4 i13_4_lut_adj_1436 (.I0(n2801), .I1(n2787), .I2(n2806), .I3(n2798), 
            .O(n37_adj_3851));
    defparam i13_4_lut_adj_1436.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1205_11 (.CI(n28672), .I0(n1701), .I1(n1730), .CO(n28673));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n28671), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n28906), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n28671), .I0(n1702), .I1(n1730), .CO(n28672));
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n27452), 
            .O(n39065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_17_lut (.I0(n19), .I1(bit_ctr[15]), .I2(GND_net), .I3(n27462), 
            .O(n39068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_23 (.CI(n28906), .I0(n2889), .I1(n2918), .CO(n28907));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n28670), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n28670), .I0(n1703), .I1(n1730), .CO(n28671));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n28905), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n28905), .I0(n2890), .I1(n2918), .CO(n28906));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n28904), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n28669), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n28669), .I0(n1704), .I1(n1730), .CO(n28670));
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_21 (.CI(n28904), .I0(n2891), .I1(n2918), .CO(n28905));
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n28668), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n39073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1205_7 (.CI(n28668), .I0(n1705), .I1(n1730), .CO(n28669));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n28903), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n28903), .I0(n2892), .I1(n2918), .CO(n28904));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n28667), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_2_lut (.I0(n2789), .I1(n2802), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_3858));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n28902), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n28902), .I0(n2893), .I1(n2918), .CO(n28903));
    SB_CARRY mod_5_add_1205_6 (.CI(n28667), .I0(n1706), .I1(n1730), .CO(n28668));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n28666), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n28901), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n28901), .I0(n2894), .I1(n2918), .CO(n28902));
    SB_CARRY mod_5_add_1205_5 (.CI(n28666), .I0(n1707), .I1(n1730), .CO(n28667));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n28900), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n28665), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_17 (.CI(n27462), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27463));
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1437 (.I0(n2804), .I1(n2795), .I2(n2800), .I3(n2808), 
            .O(n42_adj_3859));
    defparam i18_4_lut_adj_1437.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1205_4 (.CI(n28665), .I0(n1708), .I1(n1730), .CO(n28666));
    SB_LUT4 i22_4_lut_adj_1438 (.I0(n37_adj_3851), .I1(n39_adj_3840), .I2(n38_adj_3834), 
            .I3(n40_adj_3822), .O(n46_adj_3860));
    defparam i22_4_lut_adj_1438.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n41725), 
            .I3(n28664), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_7 (.CI(n27452), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27453));
    SB_CARRY mod_5_add_2009_17 (.CI(n28900), .I0(n2895), .I1(n2918), .CO(n28901));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n28899), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_3 (.CI(n28664), .I0(n1709), .I1(n41725), .CO(n28665));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27448));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n41725), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_16 (.CI(n28899), .I0(n2896), .I1(n2918), .CO(n28900));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n28898), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n28898), .I0(n2897), .I1(n2918), .CO(n28899));
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n28897), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n28897), .I0(n2898), .I1(n2918), .CO(n28898));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n28896), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n41725), 
            .CO(n28664));
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_adj_1439 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(n25384), .I3(GND_net), .O(n35817));
    defparam i2_3_lut_adj_1439.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_2009_13 (.CI(n28896), .I0(n2899), .I1(n2918), .CO(n28897));
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n27461), 
            .O(n39064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n28663), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n28662), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i43_4_lut (.I0(start), .I1(n35817), .I2(\state[1] ), .I3(n26_adj_3831), 
            .O(n17503));
    defparam i43_4_lut.LUT_INIT = 16'h3530;
    SB_CARRY mod_5_add_1138_13 (.CI(n28662), .I0(n1599), .I1(n1631), .CO(n28663));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n28895), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n28895), .I0(n2900), .I1(n2918), .CO(n28896));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n28661), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n17503), .D(\neo_pixel_transmitter.done_N_551 ), 
            .R(n33686));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_488[22]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n27666), .O(n22_adj_3800)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n28894), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_488[25]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n27665), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_11 (.CI(n28894), .I0(n2901), .I1(n2918), .CO(n28895));
    SB_CARRY sub_14_add_2_32 (.CI(n27665), .I0(timer[30]), .I1(n1[30]), 
            .CO(n27666));
    SB_CARRY mod_5_add_1138_12 (.CI(n28661), .I0(n1600), .I1(n1631), .CO(n28662));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n28660), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_488[28]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n27664), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n27451), 
            .O(n39063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_31 (.CI(n27664), .I0(timer[29]), .I1(n1[29]), 
            .CO(n27665));
    SB_LUT4 sub_14_add_2_30_lut (.I0(GND_net), .I1(timer[28]), .I2(n1[28]), 
            .I3(n27663), .O(one_wire_N_488[28])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_30 (.CI(n27663), .I0(timer[28]), .I1(n1[28]), 
            .CO(n27664));
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_551 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n28893), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n28660), .I0(n1601), .I1(n1631), .CO(n28661));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n28659), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2805), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_3862));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1440 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_3863));
    defparam i8_4_lut_adj_1440.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_488[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n27662), .O(n21_c)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n27662), .I0(timer[27]), .I1(n1[27]), 
            .CO(n27663));
    SB_CARRY mod_5_add_2009_10 (.CI(n28893), .I0(n2902), .I1(n2918), .CO(n28894));
    SB_LUT4 i1_3_lut_adj_1441 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_3864));
    defparam i1_3_lut_adj_1441.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n28892), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3865));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n13_adj_3864), .I1(n20_adj_3863), .I2(n1605), 
            .I3(n1599), .O(n22_adj_3866));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1442 (.I0(n1601), .I1(n22_adj_3866), .I2(n18_adj_3865), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1442.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_28_lut (.I0(one_wire_N_488[19]), .I1(timer[26]), 
            .I2(n1[26]), .I3(n27661), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1138_10 (.CI(n28659), .I0(n1602), .I1(n1631), .CO(n28660));
    SB_CARRY sub_14_add_2_28 (.CI(n27661), .I0(timer[26]), .I1(n1[26]), 
            .CO(n27662));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n27660), .O(one_wire_N_488[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_27 (.CI(n27660), .I0(timer[25]), .I1(n1[25]), 
            .CO(n27661));
    SB_CARRY mod_5_add_2009_9 (.CI(n28892), .I0(n2903), .I1(n2918), .CO(n28893));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n28658), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n28891), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n28658), .I0(n1603), .I1(n1631), .CO(n28659));
    SB_CARRY mod_5_add_2009_8 (.CI(n28891), .I0(n2904), .I1(n2918), .CO(n28892));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n28890), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n28890), .I0(n2905), .I1(n2918), .CO(n28891));
    SB_LUT4 sub_14_add_2_26_lut (.I0(one_wire_N_488[12]), .I1(timer[24]), 
            .I2(n1[24]), .I3(n27659), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n28657), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n28889), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n28657), .I0(n1604), .I1(n1631), .CO(n28658));
    SB_CARRY sub_14_add_2_26 (.CI(n27659), .I0(timer[24]), .I1(n1[24]), 
            .CO(n27660));
    SB_CARRY mod_5_add_2009_6 (.CI(n28889), .I0(n2906), .I1(n2918), .CO(n28890));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n28656), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_488[21]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n27658), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n27658), .I0(timer[23]), .I1(n1[23]), 
            .CO(n27659));
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n27657), .O(one_wire_N_488[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n28888), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n28656), .I0(n1605), .I1(n1631), .CO(n28657));
    SB_CARRY mod_5_add_2009_5 (.CI(n28888), .I0(n2907), .I1(n2918), .CO(n28889));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n28887), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_24 (.CI(n27657), .I0(timer[22]), .I1(n1[22]), 
            .CO(n27658));
    SB_LUT4 sub_14_add_2_23_lut (.I0(GND_net), .I1(timer[21]), .I2(n1[21]), 
            .I3(n27656), .O(one_wire_N_488[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n27451), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27452));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n28655), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_23 (.CI(n27656), .I0(timer[21]), .I1(n1[21]), 
            .CO(n27657));
    SB_CARRY mod_5_add_2009_4 (.CI(n28887), .I0(n2908), .I1(n2918), .CO(n28888));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_488[16]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n27655), .O(n30_adj_3799)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n27655), .I0(timer[20]), .I1(n1[20]), 
            .CO(n27656));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n41724), 
            .I3(n28886), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n27654), .O(one_wire_N_488[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n28886), .I0(n2909), .I1(n41724), .CO(n28887));
    SB_CARRY mod_5_add_1138_6 (.CI(n28655), .I0(n1606), .I1(n1631), .CO(n28656));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n28654), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n41724), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_5 (.CI(n28654), .I0(n1607), .I1(n1631), .CO(n28655));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n41724), 
            .CO(n28886));
    SB_CARRY sub_14_add_2_21 (.CI(n27654), .I0(timer[19]), .I1(n1[19]), 
            .CO(n27655));
    SB_CARRY add_21_16 (.CI(n27461), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27462));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n27653), .O(one_wire_N_488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n27653), .I0(timer[18]), .I1(n1[18]), 
            .CO(n27654));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_488[13]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n27652), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n27652), .I0(timer[17]), .I1(n1[17]), 
            .CO(n27653));
    SB_LUT4 i35405_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41725));
    defparam i35405_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n28885), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n27651), .O(one_wire_N_488[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n28884), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_18 (.CI(n27651), .I0(timer[16]), .I1(n1[16]), 
            .CO(n27652));
    SB_LUT4 sub_14_add_2_17_lut (.I0(one_wire_N_488[14]), .I1(timer[15]), 
            .I2(n1[15]), .I3(n27650), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_25 (.CI(n28884), .I0(n2787), .I1(n2819), .CO(n28885));
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n27460), 
            .O(n39076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_17 (.CI(n27650), .I0(timer[15]), .I1(n1[15]), 
            .CO(n27651));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n27649), .O(one_wire_N_488[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n28883), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n28653), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n28883), .I0(n2788), .I1(n2819), .CO(n28884));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n28882), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n28653), .I0(n1608), .I1(n1631), .CO(n28654));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n41726), 
            .I3(n28652), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_16 (.CI(n27649), .I0(timer[14]), .I1(n1[14]), 
            .CO(n27650));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n27648), .O(one_wire_N_488[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_3 (.CI(n28652), .I0(n1609), .I1(n41726), .CO(n28653));
    SB_CARRY sub_14_add_2_15 (.CI(n27648), .I0(timer[13]), .I1(n1[13]), 
            .CO(n27649));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n27647), .O(one_wire_N_488[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n27647), .I0(timer[12]), .I1(n1[12]), 
            .CO(n27648));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n27646), .O(one_wire_N_488[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n27646), .I0(timer[11]), .I1(n1[11]), 
            .CO(n27647));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n41726), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n41726), 
            .CO(n28652));
    SB_LUT4 sub_14_add_2_12_lut (.I0(one_wire_N_488[9]), .I1(timer[10]), 
            .I2(n1[10]), .I3(n27645), .O(n24843)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_23 (.CI(n28882), .I0(n2789), .I1(n2819), .CO(n28883));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n28651), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_12 (.CI(n27645), .I0(timer[10]), .I1(n1[10]), 
            .CO(n27646));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n27644), .O(one_wire_N_488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n28881), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n28650), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_11 (.CI(n27644), .I0(timer[9]), .I1(n1[9]), 
            .CO(n27645));
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_488[11]), .I1(timer[8]), 
            .I2(n1[8]), .I3(n27643), .O(n9_adj_3827)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_10 (.CI(n27643), .I0(timer[8]), .I1(n1[8]), 
            .CO(n27644));
    SB_LUT4 sub_14_add_2_9_lut (.I0(n16437), .I1(timer[7]), .I2(n1[7]), 
            .I3(n27642), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_15 (.CI(n27460), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27461));
    SB_CARRY sub_14_add_2_9 (.CI(n27642), .I0(timer[7]), .I1(n1[7]), .CO(n27643));
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_488[5]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n27641), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1071_12 (.CI(n28650), .I0(n1500), .I1(n1532), .CO(n28651));
    SB_CARRY sub_14_add_2_8 (.CI(n27641), .I0(timer[6]), .I1(n1[6]), .CO(n27642));
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n27459), 
            .O(n39075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n27640), .O(one_wire_N_488[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n27640), .I0(timer[5]), .I1(n1[5]), .CO(n27641));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n27639), .O(one_wire_N_488[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n27639), .I0(timer[4]), .I1(n1[4]), .CO(n27640));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n27638), .O(one_wire_N_488[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n27638), .I0(timer[3]), .I1(n1[3]), .CO(n27639));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n27637), .O(one_wire_N_488[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_22 (.CI(n28881), .I0(n2790), .I1(n2819), .CO(n28882));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n28649), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_4 (.CI(n27637), .I0(timer[2]), .I1(n1[2]), .CO(n27638));
    SB_LUT4 i23_4_lut (.I0(n33_adj_3862), .I1(n46_adj_3860), .I2(n42_adj_3859), 
            .I3(n34_adj_3858), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1443 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_3867));
    defparam i7_4_lut_adj_1443.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_14 (.CI(n27459), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27460));
    SB_LUT4 i9_4_lut_adj_1444 (.I0(n1705), .I1(n1703), .I2(n1700), .I3(n1699), 
            .O(n22_adj_3868));
    defparam i9_4_lut_adj_1444.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_3869));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_4_lut_adj_1445 (.I0(n1698), .I1(n1702), .I2(n1707), .I3(n1697), 
            .O(n21_adj_3870));
    defparam i8_4_lut_adj_1445.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut (.I0(n1706), .I1(bit_ctr[18]), .I2(n1709), .I3(GND_net), 
            .O(n19_adj_3871));
    defparam i6_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1446 (.I0(n19_adj_3871), .I1(n21_adj_3870), .I2(n20_adj_3869), 
            .I3(n22_adj_3868), .O(n1730));
    defparam i12_4_lut_adj_1446.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut_adj_1447 (.I0(bit_ctr[6]), .I1(n2888), .I2(n2909), 
            .I3(GND_net), .O(n34_adj_3872));
    defparam i9_3_lut_adj_1447.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1448 (.I0(n2897), .I1(n2891), .I2(n2893), .I3(n2892), 
            .O(n41_adj_3873));
    defparam i16_4_lut_adj_1448.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2901), .I1(n2889), .I2(n2903), .I3(GND_net), 
            .O(n38_adj_3874));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1449 (.I0(n2886), .I1(n2885), .I2(n2898), .I3(n2894), 
            .O(n43_adj_3875));
    defparam i18_4_lut_adj_1449.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1450 (.I0(n2902), .I1(n2887), .I2(n2896), .I3(n2895), 
            .O(n40_adj_3876));
    defparam i15_4_lut_adj_1450.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1451 (.I0(n41_adj_3873), .I1(n2890), .I2(n34_adj_3872), 
            .I3(n2905), .O(n46_adj_3877));
    defparam i21_4_lut_adj_1451.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1452 (.I0(n2904), .I1(n2906), .I2(n2908), .I3(n2900), 
            .O(n39_adj_3878));
    defparam i14_4_lut_adj_1452.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1453 (.I0(n43_adj_3875), .I1(n2907), .I2(n38_adj_3874), 
            .I3(n2899), .O(n47_adj_3879));
    defparam i22_4_lut_adj_1453.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_3879), .I1(n39_adj_3878), .I2(n46_adj_3877), 
            .I3(n40_adj_3876), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35403_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41723));
    defparam i35403_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35402_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41722));
    defparam i35402_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1454 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_3880));
    defparam i10_4_lut_adj_1454.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1455 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_3881));
    defparam i8_4_lut_adj_1455.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1456 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_3882));
    defparam i9_4_lut_adj_1456.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1457 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_3883));
    defparam i7_3_lut_adj_1457.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1458 (.I0(n21_adj_3883), .I1(n23_adj_3882), .I2(n22_adj_3881), 
            .I3(n24_adj_3880), .O(n1829));
    defparam i13_4_lut_adj_1458.LUT_INIT = 16'hfffe;
    SB_LUT4 i35401_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41721));
    defparam i35401_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1459 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_3884));
    defparam i14_4_lut_adj_1459.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1460 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_3885));
    defparam i18_4_lut_adj_1460.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1461 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_3886));
    defparam i16_4_lut_adj_1461.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1462 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_3887));
    defparam i17_4_lut_adj_1462.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1463 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_3888));
    defparam i15_4_lut_adj_1463.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_3889));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_3884), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_3890));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1464 (.I0(n41_adj_3888), .I1(n43_adj_3887), .I2(n42_adj_3886), 
            .I3(n44_adj_3885), .O(n50));
    defparam i24_4_lut_adj_1464.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_3891));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_3891), .I1(n50), .I2(n46_adj_3890), 
            .I3(n38_adj_3889), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35399_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41719));
    defparam i35399_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1465 (.I0(n1906), .I1(n1900), .I2(n1905), .I3(n1895), 
            .O(n26_adj_3892));
    defparam i11_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1466 (.I0(n1902), .I1(n1897), .I2(n1908), .I3(n1901), 
            .O(n24_adj_3893));
    defparam i9_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1467 (.I0(n1899), .I1(n1904), .I2(n1896), .I3(n1903), 
            .O(n25_adj_3894));
    defparam i10_4_lut_adj_1467.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1468 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1898), 
            .I3(n1909), .O(n23_adj_3895));
    defparam i8_4_lut_adj_1468.LUT_INIT = 16'hfefa;
    SB_LUT4 i14_4_lut_adj_1469 (.I0(n23_adj_3895), .I1(n25_adj_3894), .I2(n24_adj_3893), 
            .I3(n26_adj_3892), .O(n1928));
    defparam i14_4_lut_adj_1469.LUT_INIT = 16'hfffe;
    SB_LUT4 i35400_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41720));
    defparam i35400_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1470 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3896));
    defparam i2_2_lut_adj_1470.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1471 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_3897));
    defparam i12_4_lut_adj_1471.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1472 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_3898));
    defparam i10_4_lut_adj_1472.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1473 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_3899));
    defparam i11_4_lut_adj_1473.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1474 (.I0(bit_ctr[15]), .I1(n18_adj_3896), .I2(n2006), 
            .I3(n2009), .O(n25_adj_3900));
    defparam i9_4_lut_adj_1474.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1475 (.I0(n25_adj_3900), .I1(n27_adj_3899), .I2(n26_adj_3898), 
            .I3(n28_adj_3897), .O(n2027));
    defparam i15_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i35397_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41717));
    defparam i35397_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21038_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n25528));
    defparam i21038_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1476 (.I0(n3196), .I1(n3208), .I2(n3199), .I3(n3188), 
            .O(n48_adj_3901));
    defparam i20_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1477 (.I0(n3195), .I1(n3202), .I2(n3187), .I3(n3194), 
            .O(n46_adj_3902));
    defparam i18_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1478 (.I0(n3200), .I1(n3185), .I2(n3182), .I3(n3192), 
            .O(n47_adj_3903));
    defparam i19_4_lut_adj_1478.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1479 (.I0(n3201), .I1(n3197), .I2(n3190), .I3(n3183), 
            .O(n45_adj_3904));
    defparam i17_4_lut_adj_1479.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1480 (.I0(n3184), .I1(n3205), .I2(n3206), .I3(n3186), 
            .O(n44_adj_3905));
    defparam i16_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1481 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n25528), 
            .O(n43_adj_3906));
    defparam i15_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1482 (.I0(n45_adj_3904), .I1(n47_adj_3903), .I2(n46_adj_3902), 
            .I3(n48_adj_3901), .O(n54_adj_3907));
    defparam i26_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1483 (.I0(n3191), .I1(n3207), .I2(n3204), .I3(n3203), 
            .O(n49_adj_3908));
    defparam i21_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1484 (.I0(n49_adj_3908), .I1(n54_adj_3907), .I2(n43_adj_3906), 
            .I3(n44_adj_3905), .O(n25560));
    defparam i27_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\state_3__N_337[1] ), .I1(n41779), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3909));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut (.I0(n5_adj_3909), .I1(n3209), .I2(bit_ctr[3]), .I3(n25560), 
            .O(state_3__N_337[0]));
    defparam i3_4_lut.LUT_INIT = 16'h2008;
    SB_LUT4 i12_3_lut_4_lut (.I0(n175), .I1(\state[0] ), .I2(n57), .I3(\state[1] ), 
            .O(n17721));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h03aa;
    SB_LUT4 i15_4_lut_adj_1486 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_3910));
    defparam i15_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1487 (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_3911));
    defparam i19_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1488 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44_adj_3912));
    defparam i17_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1489 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45_adj_3913));
    defparam i18_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1490 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43_adj_3914));
    defparam i16_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1491 (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), 
            .I3(GND_net), .O(n40_adj_3915));
    defparam i13_3_lut_adj_1491.LUT_INIT = 16'hecec;
    SB_LUT4 i9_4_lut_adj_1492 (.I0(n1504), .I1(n18_adj_3867), .I2(n1502), 
            .I3(n1499), .O(n20_adj_3916));
    defparam i9_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1493 (.I0(n3107), .I1(n42_adj_3910), .I2(n3087), 
            .I3(n3086), .O(n48_adj_3917));
    defparam i21_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1494 (.I0(n43_adj_3914), .I1(n45_adj_3913), .I2(n44_adj_3912), 
            .I3(n46_adj_3911), .O(n52));
    defparam i25_4_lut_adj_1494.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1495 (.I0(n3095), .I1(n3084), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3918));
    defparam i12_2_lut_adj_1495.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut_adj_1496 (.I0(n39_adj_3918), .I1(n52), .I2(n48_adj_3917), 
            .I3(n40_adj_3915), .O(n3116));
    defparam i26_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), .I3(GND_net), 
            .O(n15_adj_3919));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n29806));   // verilog/neopixel.v(22[26:36])
    defparam i1_3_lut_4_lut_3_lut.LUT_INIT = 16'h9494;
    SB_LUT4 i35384_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41704));
    defparam i35384_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n136), .I3(n168), .O(n131));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h2220;
    SB_LUT4 i35385_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41705));
    defparam i35385_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(n34361), .I1(n15157), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1_2_lut_adj_1497 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_3920));
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'heeee;
    SB_LUT4 i20857_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n25344));
    defparam i20857_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1498 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_3920), 
            .O(n30_adj_3921));
    defparam i13_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1499 (.I0(n2098), .I1(n25344), .I2(n2094), .I3(n2099), 
            .O(n28_adj_3922));
    defparam i11_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1500 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_3923));
    defparam i12_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1501 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_3924));
    defparam i10_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1502 (.I0(n27_adj_3924), .I1(n29_adj_3923), .I2(n28_adj_3922), 
            .I3(n30_adj_3921), .O(n2126));
    defparam i16_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i35396_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41716));
    defparam i35396_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\neo_pixel_transmitter.done ), 
            .I3(n25384), .O(n33686));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i30897_2_lut_3_lut (.I0(n168), .I1(n165), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n37149));
    defparam i30897_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i3736_2_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[28]), .O(n7534));   // verilog/neopixel.v(22[26:36])
    defparam i3736_2_lut_4_lut.LUT_INIT = 16'h9400;
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n37366), .I2(n37367), 
            .I3(bit_ctr[2]), .O(n41776));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n41776_bdd_4_lut (.I0(n41776), .I1(n37310), .I2(n37309), .I3(bit_ctr[2]), 
            .O(n41779));
    defparam n41776_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i33142_2_lut_3_lut (.I0(start), .I1(\state[1] ), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n39062));
    defparam i33142_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i35365_2_lut_3_lut (.I0(start), .I1(\state[1] ), .I2(n26_adj_3831), 
            .I3(GND_net), .O(n33752));
    defparam i35365_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n37097), .I3(n168), .O(n175));   // verilog/neopixel.v(16[20:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h2220;
    SB_LUT4 i12_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam i12_3_lut_4_lut_3_lut.LUT_INIT = 16'h4242;
    SB_LUT4 i3746_2_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(bit_ctr[29]), .I3(bit_ctr[28]), .O(n62));   // verilog/neopixel.v(22[26:36])
    defparam i3746_2_lut_4_lut_4_lut.LUT_INIT = 16'hd642;
    SB_LUT4 i33334_3_lut_4_lut (.I0(n62), .I1(bit_ctr[28]), .I2(n29806), 
            .I3(GND_net), .O(n34361));   // verilog/neopixel.v(22[26:36])
    defparam i33334_3_lut_4_lut.LUT_INIT = 16'h7878;
    SB_LUT4 mod_5_i538_3_lut_4_lut (.I0(n62), .I1(n7534), .I2(n708), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut_4_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i1_2_lut_3_lut (.I0(n62), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(GND_net), .O(n15157));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n15157), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n34361), .O(n34363));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i1_2_lut_4_lut_adj_1503 (.I0(\neo_pixel_transmitter.done ), .I1(n16437), 
            .I2(one_wire_N_488[11]), .I3(n24843), .O(n57));
    defparam i1_2_lut_4_lut_adj_1503.LUT_INIT = 16'habbb;
    SB_LUT4 i10_4_lut_adj_1504 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_3925));
    defparam i10_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1505 (.I0(n2203), .I1(n28_adj_3925), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_3926));
    defparam i14_4_lut_adj_1505.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1506 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_3927));
    defparam i12_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1507 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_3928));
    defparam i13_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1508 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_3929));
    defparam i11_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1509 (.I0(n29_adj_3929), .I1(n31_adj_3928), .I2(n30_adj_3927), 
            .I3(n32_adj_3926), .O(n2225));
    defparam i17_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i35395_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41715));
    defparam i35395_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1510 (.I0(\state[0] ), .I1(n175), .I2(n57), .I3(\state[1] ), 
            .O(n17561));
    defparam i1_4_lut_adj_1510.LUT_INIT = 16'hafcc;
    SB_LUT4 i10_4_lut_adj_1511 (.I0(n15_adj_3919), .I1(n20_adj_3916), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, n18368, \data_in_frame[15] , n18367, n18366, 
            n18365, GND_net, \data_in_frame[2] , \data_in_frame[6] , 
            \data_in_frame[1] , \data_in_frame[5] , \data_in_frame[19] , 
            \data_in_frame[18] , \data_in_frame[17] , rx_data, n18372, 
            n18371, n18370, n18369, n41916, VCC_net, \byte_transmit_counter[0] , 
            n18427, control_mode, n18428, PWMLimit, n18429, n18430, 
            n18431, n18432, n18433, n18421, n18422, n18423, n18424, 
            \data_in_frame[7] , n18447, n18448, n18449, n18450, n18445, 
            n18446, n18443, n18444, n18441, n18442, n18439, n18440, 
            n18437, n18438, n18434, n18435, n18436, n18425, n18426, 
            n18245, \data_out_frame[20] , n18244, n18243, n18242, 
            n18241, n18240, n18239, n18238, n18237, \data_out_frame[19] , 
            n18236, n18235, n18234, n18233, n18232, n18231, n18230, 
            n18229, \data_out_frame[18] , n18228, n18227, n18226, 
            \data_out_frame[5] , \byte_transmit_counter[1] , \data_out_frame[6] , 
            \data_out_frame[7] , n21, n18225, n18224, n18223, n18222, 
            n18221, \data_out_frame[17] , n18220, n35752, n18219, 
            n18218, n18217, n18216, n18215, n18214, n18213, \data_out_frame[16] , 
            n18212, n18211, n18210, n18209, n18208, n18207, n18206, 
            n18205, \data_out_frame[15] , n18204, n18203, n18202, 
            n18201, n18200, n18199, n18198, n18197, \data_out_frame[14] , 
            n18196, n18195, n18194, rx_data_ready, n18193, n18192, 
            n18191, n18190, n18189, \data_out_frame[13] , n18188, 
            \FRAME_MATCHER.state[0] , n36216, n18187, n18186, n18185, 
            n18184, n18183, n18182, n18181, \data_out_frame[12] , 
            n18180, n18179, n18178, n18177, n18176, n18175, n18174, 
            n18173, \data_out_frame[11] , n18172, n18171, n18170, 
            n18169, n18168, n18167, n18166, n18165, \data_out_frame[10] , 
            n18164, n18163, \data_in[1] , \data_in[0] , \data_in[3] , 
            \data_in[2] , n18162, n18161, n18160, n18159, n18158, 
            n18157, \data_out_frame[9] , n18156, n18155, n18154, n18153, 
            n18152, n18151, n18150, n18149, \data_out_frame[8] , n3761, 
            n16420, n18148, n18147, n18146, n18145, n18144, n18143, 
            n18142, n25598, n18141, n18140, n18139, n18138, n18137, 
            n18136, n18135, n18134, n18133, n18132, n18131, n35990, 
            n18130, n18129, n18128, n18127, n18126, n18125, n18124, 
            n18123, n18122, n18121, n18120, n18119, n18118, n63, 
            n123, n16404, n2857, n5, n18114, \Kp[7] , n18113, 
            \Kp[6] , n42588, n18112, \Kp[5] , n18111, \Kp[4] , n18110, 
            \Kp[3] , n18109, \Kp[2] , n18108, \Kp[1] , n18107, n16405, 
            n37137, n18106, n18105, n9783, n18104, n18103, n18102, 
            n18101, n18100, n18099, n18098, n18097, n18096, n18095, 
            n18094, n18093, n18092, n18091, n18090, n18089, n18088, 
            n18087, n18086, n18085, n18084, n18083, n18082, n18081, 
            n18080, n18079, n18078, n18077, n18075, gearBoxRatio, 
            n18074, n18073, n18072, n18071, n18070, n18069, n18068, 
            n18067, n18066, n18065, n18064, n18063, n18062, n18061, 
            n18060, n18059, n18058, n18057, n18056, n18055, n18054, 
            n18053, n17974, setpoint, n17973, n17972, n17971, n17970, 
            n17969, n17968, n17967, n17966, n17965, n17964, n17963, 
            n17962, n17961, n17960, n17959, n17958, n17957, n17956, 
            n17955, n17954, n17953, n17952, LED_c, n18308, n18307, 
            \data_out_frame[21] , n35420, \data_out_frame[22] , n34307, 
            n18306, n18305, n18304, n18303, \r_SM_Main_2__N_3298[0] , 
            n18302, tx_active, n18301, n33144, n17896, n17895, n17893, 
            \Kp[0] , n17793, n17791, n17892, n11748, n34073, n19, 
            n33787, n33923, n33775, n33766, n16417, n30686, n4423, 
            n4446, n13950, n4445, n4444, n4443, n4442, n4441, 
            n4440, n4439, n37188, n4438, n4437, n4436, n4435, 
            n4434, n4433, n16809, n4432, n4431, n4430, n4429, 
            n4428, n4427, n4426, n4425, n4424, n18509, r_SM_Main, 
            n17827, r_Bit_Index, n17830, \r_SM_Main_2__N_3295[1] , n17625, 
            n17748, n4706, n17989, tx_o, tx_enable, n18539, \r_Clock_Count[0] , 
            n17836, r_Bit_Index_adj_10, n17833, \r_SM_Main[1]_adj_6 , 
            \r_SM_Main[2]_adj_7 , n2346, r_Rx_Data, PIN_13_N_106, \r_Clock_Count[2] , 
            \r_Clock_Count[1] , \r_Clock_Count[6] , \r_Clock_Count[4] , 
            n16429, n4, n35922, n4684, n17619, n17746, n17931, 
            n17936, n17942, n17980, n17992, n18003, n33396, n220, 
            n222, n224, n225, n226, n24632, n4_adj_8, n4_adj_9, 
            n16424, n17843, n17842, n17841, n17840, n17839, n17838, 
            n17837, n17522) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n18368;
    output [7:0]\data_in_frame[15] ;
    input n18367;
    input n18366;
    input n18365;
    input GND_net;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[17] ;
    output [7:0]rx_data;
    input n18372;
    input n18371;
    input n18370;
    input n18369;
    input n41916;
    input VCC_net;
    output \byte_transmit_counter[0] ;
    input n18427;
    output [7:0]control_mode;
    input n18428;
    output [23:0]PWMLimit;
    input n18429;
    input n18430;
    input n18431;
    input n18432;
    input n18433;
    input n18421;
    input n18422;
    input n18423;
    input n18424;
    output [7:0]\data_in_frame[7] ;
    input n18447;
    input n18448;
    input n18449;
    input n18450;
    input n18445;
    input n18446;
    input n18443;
    input n18444;
    input n18441;
    input n18442;
    input n18439;
    input n18440;
    input n18437;
    input n18438;
    input n18434;
    input n18435;
    input n18436;
    input n18425;
    input n18426;
    input n18245;
    output [7:0]\data_out_frame[20] ;
    input n18244;
    input n18243;
    input n18242;
    input n18241;
    input n18240;
    input n18239;
    input n18238;
    input n18237;
    output [7:0]\data_out_frame[19] ;
    input n18236;
    input n18235;
    input n18234;
    input n18233;
    input n18232;
    input n18231;
    input n18230;
    input n18229;
    output [7:0]\data_out_frame[18] ;
    input n18228;
    input n18227;
    input n18226;
    output [7:0]\data_out_frame[5] ;
    output \byte_transmit_counter[1] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    input n21;
    input n18225;
    input n18224;
    input n18223;
    input n18222;
    input n18221;
    output [7:0]\data_out_frame[17] ;
    input n18220;
    output n35752;
    input n18219;
    input n18218;
    input n18217;
    input n18216;
    input n18215;
    input n18214;
    input n18213;
    output [7:0]\data_out_frame[16] ;
    input n18212;
    input n18211;
    input n18210;
    input n18209;
    input n18208;
    input n18207;
    input n18206;
    input n18205;
    output [7:0]\data_out_frame[15] ;
    input n18204;
    input n18203;
    input n18202;
    input n18201;
    input n18200;
    input n18199;
    input n18198;
    input n18197;
    output [7:0]\data_out_frame[14] ;
    input n18196;
    input n18195;
    input n18194;
    output rx_data_ready;
    input n18193;
    input n18192;
    input n18191;
    input n18190;
    input n18189;
    output [7:0]\data_out_frame[13] ;
    input n18188;
    output \FRAME_MATCHER.state[0] ;
    output n36216;
    input n18187;
    input n18186;
    input n18185;
    input n18184;
    input n18183;
    input n18182;
    input n18181;
    output [7:0]\data_out_frame[12] ;
    input n18180;
    input n18179;
    input n18178;
    input n18177;
    input n18176;
    input n18175;
    input n18174;
    input n18173;
    output [7:0]\data_out_frame[11] ;
    input n18172;
    input n18171;
    input n18170;
    input n18169;
    input n18168;
    input n18167;
    input n18166;
    input n18165;
    output [7:0]\data_out_frame[10] ;
    input n18164;
    input n18163;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[2] ;
    input n18162;
    input n18161;
    input n18160;
    input n18159;
    input n18158;
    input n18157;
    output [7:0]\data_out_frame[9] ;
    input n18156;
    input n18155;
    input n18154;
    input n18153;
    input n18152;
    input n18151;
    input n18150;
    input n18149;
    output [7:0]\data_out_frame[8] ;
    output n3761;
    output n16420;
    input n18148;
    input n18147;
    input n18146;
    input n18145;
    input n18144;
    input n18143;
    input n18142;
    output n25598;
    input n18141;
    input n18140;
    input n18139;
    input n18138;
    input n18137;
    input n18136;
    input n18135;
    input n18134;
    input n18133;
    input n18132;
    input n18131;
    output n35990;
    input n18130;
    input n18129;
    input n18128;
    input n18127;
    input n18126;
    input n18125;
    input n18124;
    input n18123;
    input n18122;
    input n18121;
    input n18120;
    input n18119;
    input n18118;
    output n63;
    output n123;
    output n16404;
    output n2857;
    output n5;
    input n18114;
    output \Kp[7] ;
    input n18113;
    output \Kp[6] ;
    output n42588;
    input n18112;
    output \Kp[5] ;
    input n18111;
    output \Kp[4] ;
    input n18110;
    output \Kp[3] ;
    input n18109;
    output \Kp[2] ;
    input n18108;
    output \Kp[1] ;
    input n18107;
    output n16405;
    output n37137;
    input n18106;
    input n18105;
    output n9783;
    input n18104;
    input n18103;
    input n18102;
    input n18101;
    input n18100;
    input n18099;
    input n18098;
    input n18097;
    input n18096;
    input n18095;
    input n18094;
    input n18093;
    input n18092;
    input n18091;
    input n18090;
    input n18089;
    input n18088;
    input n18087;
    input n18086;
    input n18085;
    input n18084;
    input n18083;
    input n18082;
    input n18081;
    input n18080;
    input n18079;
    input n18078;
    input n18077;
    input n18075;
    output [23:0]gearBoxRatio;
    input n18074;
    input n18073;
    input n18072;
    input n18071;
    input n18070;
    input n18069;
    input n18068;
    input n18067;
    input n18066;
    input n18065;
    input n18064;
    input n18063;
    input n18062;
    input n18061;
    input n18060;
    input n18059;
    input n18058;
    input n18057;
    input n18056;
    input n18055;
    input n18054;
    input n18053;
    input n17974;
    output [23:0]setpoint;
    input n17973;
    input n17972;
    input n17971;
    input n17970;
    input n17969;
    input n17968;
    input n17967;
    input n17966;
    input n17965;
    input n17964;
    input n17963;
    input n17962;
    input n17961;
    input n17960;
    input n17959;
    input n17958;
    input n17957;
    input n17956;
    input n17955;
    input n17954;
    input n17953;
    input n17952;
    output LED_c;
    input n18308;
    input n18307;
    output [7:0]\data_out_frame[21] ;
    input n35420;
    output [7:0]\data_out_frame[22] ;
    output n34307;
    input n18306;
    input n18305;
    input n18304;
    input n18303;
    output \r_SM_Main_2__N_3298[0] ;
    input n18302;
    output tx_active;
    input n18301;
    input n33144;
    input n17896;
    input n17895;
    input n17893;
    output \Kp[0] ;
    input n17793;
    input n17791;
    input n17892;
    output n11748;
    output n34073;
    input n19;
    output n33787;
    output n33923;
    output n33775;
    output n33766;
    output n16417;
    output n30686;
    output n4423;
    output n4446;
    output n13950;
    output n4445;
    output n4444;
    output n4443;
    output n4442;
    output n4441;
    output n4440;
    output n4439;
    input n37188;
    output n4438;
    output n4437;
    output n4436;
    output n4435;
    output n4434;
    output n4433;
    output n16809;
    output n4432;
    output n4431;
    output n4430;
    output n4429;
    output n4428;
    output n4427;
    output n4426;
    output n4425;
    output n4424;
    input n18509;
    output [2:0]r_SM_Main;
    input n17827;
    output [2:0]r_Bit_Index;
    input n17830;
    output \r_SM_Main_2__N_3295[1] ;
    output n17625;
    output n17748;
    output n4706;
    input n17989;
    output tx_o;
    output tx_enable;
    input n18539;
    output \r_Clock_Count[0] ;
    input n17836;
    output [2:0]r_Bit_Index_adj_10;
    input n17833;
    output \r_SM_Main[1]_adj_6 ;
    output \r_SM_Main[2]_adj_7 ;
    output n2346;
    output r_Rx_Data;
    input PIN_13_N_106;
    output \r_Clock_Count[2] ;
    output \r_Clock_Count[1] ;
    output \r_Clock_Count[6] ;
    output \r_Clock_Count[4] ;
    output n16429;
    output n4;
    output n35922;
    output n4684;
    output n17619;
    output n17746;
    input n17931;
    input n17936;
    input n17942;
    input n17980;
    input n17992;
    input n18003;
    input n33396;
    output n220;
    output n222;
    output n224;
    output n225;
    output n226;
    output n24632;
    output n4_adj_8;
    output n4_adj_9;
    output n16424;
    input n17843;
    input n17842;
    input n17841;
    input n17840;
    input n17839;
    input n17838;
    input n17837;
    output n17522;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n18330;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    
    wire n18329, n18364;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n18363, n18362, n27520;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n27521, n18361, n18360, n18359, n18358, n18328, n18339;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    
    wire n18278;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    
    wire n33380, n27495, n6, n18277, n18276;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    
    wire n18275, n18338, n18337, n33352, n3, n34254, n30655, n6_adj_3566, 
        n30633, n27496, n18274, n18273, n18272, n18271, n18270, 
        n18269, n18268, n18336, n18267, n9, n16624, n2, n27519, 
        n18266, n33378, n27494, n18265, n18264, n18263, n18262, 
        n18261, n18260, n18290, n18289, n18288, n18287, n17338, 
        n4_c, n18400, n18259, n18399, n18258, n18257, n18398, 
        n18256, n18255, n18254, n18397, n18286, n18253, n18285, 
        n18252;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n18284, n18396, n18395, n18394, n18393, n18392, n18391, 
        n18390, n18389, n18388, n18387, n18386, n18385, n18384;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    
    wire n33952, n8, n33776, n18383, n18382, n18381;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    
    wire n16617, n34224;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    
    wire n33903, n18380;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n18379, n18378, n18377, n18376, n16715, n33986, n18375, 
        n34221, n16796, n18374, n18373, n18335, n18540;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n18541, n18542, n18543, n18544;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n18521, n17170, n16789, n34308, n18419;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n18420, n18408;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n18409, n18327, n18326, n18325, Kp_23__N_868, n34129, n18251, 
        n18324, n18323, n18322, n18321, n18250, n33856, n18249, 
        n18410, n18411, n18412, n18413, n18414, n18415, n18416, 
        n18417, n18418, n18248, n34260, n18247, n18246, n18406, 
        n18407, n18404, n18405, n2_adj_3567, n27518, n17114, n18283, 
        n12, n33376, n27493, n17187, n6_adj_3568, n18334, n16833, 
        n18320, n18282, n17037, n18281, Kp_23__N_1537, n34906, n30661, 
        n34239, n18280, n29784, n29824, n34039, n30670, n10, n29900, 
        n33968, n16937, n10_adj_3569, n35103, n30201, n39361, n5_c, 
        n14, n41767, n22, n38883, n37285, n16824, n30393, n34136, 
        n37287, n32806, n27517, n16, n12_adj_3570, n29915, n34329, 
        n34090, n33843, n6_adj_3571, n34227;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n16964, n33990, n17145, n12_adj_3572, n16093, n33374, n27492, 
        n33895, Kp_23__N_1058, n33852, n6_adj_3573, n34153, n10_adj_3574, 
        n7, n29840, n16741, n6_adj_3575, n18319, n18318, n18317, 
        n16952, n8_adj_3576, n33767, n24585, n16280, n29826, n35995, 
        Kp_23__N_1319, n30610, n30677, n14_adj_3577, n18316, n15, 
        n32808, n27516, n6_adj_3578, n6_adj_3579, n18, n34218, n20, 
        n29870, n34015, n4_adj_3580, n34203, n33849, n19_c, n6_adj_3581, 
        n34070, n30333, n5_adj_3582, n42567, n33811, n12_adj_3583, 
        n14_adj_3584, n34263, n17357, n33823, n15_adj_3585, \FRAME_MATCHER.rx_data_ready_prev , 
        n29818, n34093, n10_adj_3586, n29890, n35078, n34033, n35005, 
        n18333, n29928, n6_adj_3587, n35975, n18332, n35214, n27491, 
        n33801, n30720, n36127, n36135, n22_adj_3588, n34944, n34105, 
        n15_adj_3589, n10_adj_3590, n34027, n14_adj_3591, n34076, 
        n36136, n24, n36064, n37172, n31, n7_adj_3592, n24558, 
        n47, n18401, n33790, n33678, n211, n6_adj_3593, n25604, 
        n34012, n8_adj_3594, n34048, n16778, n6_adj_3595, n32810, 
        n27515, n4_adj_3596, n3_adj_3597, n17155, n4_adj_3598, n34099, 
        n29852, n6_adj_3599, Kp_23__N_833, n33943, n33792, n164, 
        n16_adj_3600, n17, n16397, n16295, n16_adj_3601, n17_adj_3602, 
        n33804, n63_c, n16394, n18_adj_3603, n20_adj_3604, n15_adj_3605, 
        n63_adj_3606, n10_adj_3607, n16466, n16406, n33898, n34290, 
        n6_adj_3608, n33929, n18_adj_3609, n30, n33807, n28, n29, 
        n34123, n27, n4_adj_3610, n14_adj_3611, n14_adj_3612, n13, 
        n13_adj_3613, n15_adj_3614, Kp_23__N_871, n16_adj_3615, n30692, 
        n28_adj_3616, n26, n17141, n27_adj_3617, n25, n31_adj_3618, 
        n24560, n5_adj_3619, n13888, n4_adj_3620, n19473, n25566, 
        n32816, n27514, n32824, n27513, n38993, n32832, n27512, 
        n4_adj_3621, n39102, n32898, n19484, n18020, n42, n40, 
        n41, n39, n38, n32846, n27511, n37, n48, n43, n16403, 
        n18403, n10_adj_3622, n16469, n37145, n15_adj_3623, n10_adj_3624, 
        n14_adj_3625, n20_adj_3626, n18117;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    
    wire n18116, n18115, n19_adj_3627, n37178, n32860, n27510, n16256, 
        n32874, n27509, n38991, n9818, n32892, n27508, n32938, 
        n27507, n38992, n32956, n27506, n34492, n13746;
    wire [31:0]\FRAME_MATCHER.state_31__N_2467 ;
    
    wire n6_adj_3630, n32978, n27505, n6_adj_3631, n38994, n33372, 
        n3_adj_3632, n18292, n18315, n18314, n18313, n18312, n18311, 
        n18310, n18309, n3_adj_3633, n34018, n34140, n3_adj_3634, 
        n3_adj_3635, n3_adj_3636, n33242, n3_adj_3637, n33192, n3_adj_3638, 
        n33110, n3_adj_3639, n33090, n3_adj_3640, n33076, n3_adj_3641, 
        n33054, n3_adj_3642, n33036, n3_adj_3643, n33018, n3_adj_3644, 
        n33004, n3_adj_3645, n3_adj_3646, n3_adj_3647, n3_adj_3648, 
        n3_adj_3649, n3_adj_3650, n3_adj_3651, n3_adj_3652, n3_adj_3653, 
        n3_adj_3654, n3_adj_3655, n3_adj_3656, n3_adj_3657, n3_adj_3658, 
        n3_adj_3659, n3_adj_3660, n2_adj_3661, n3_adj_3662, n2_adj_3663, 
        n3_adj_3664, n34115, n17572, n36123;
    wire [7:0]\data_out_frame[21]_c ;   // verilog/coms.v(95[12:26])
    
    wire n35111, n34814, n34884, n35096, n34928, n35199;
    wire [7:0]\data_out_frame[22]_c ;   // verilog/coms.v(95[12:26])
    
    wire n35129, n34031, n33912, n34046, n34084, n34249, n33126, 
        n42066, n33140, n33382, n33296, n33142, n33300, n33190, 
        n33304, n33188, n33292, n33198, n33308, n33186, n33312, 
        n33184, n33316, n33182, n33320, n33180, n33284, n33218, 
        n64, n33134, n24574, n25301, n7_adj_3665, n8_adj_3666, n33324, 
        n33174, n7_adj_3667, n8_adj_3668, n7_adj_3669, n8_adj_3670, 
        n33328, n33172, n33332, n33170, n33336, n33168, n33340, 
        n33166, n7_adj_3671, n8_adj_3672, n33288, n33200, n33344, 
        n33164, n33348, n33162, n7_adj_3673, n8_adj_3674, n33258, 
        n33228, n33262, n33160, n33274, n33158, n7_adj_3675, n8_adj_3676, 
        n10_adj_3677, n16410, n18357, n2540, n39174, n34543, n27504, 
        tx_transmit_N_3190, n10_adj_3678, n18356, n18355, n18354, 
        n18353, n18352, n18300, n18299, n18298, n18331, n16_adj_3679, 
        n22_adj_3680, n20_adj_3681, n24_adj_3682, n33788, n33971, 
        Kp_23__N_1444, n12_adj_3683, n13_adj_3684, n18291, n30710, 
        n34206, n33983, Kp_23__N_1328, n6_adj_3685, n16285, n34021, 
        n33940, n12_adj_3686, n14_adj_3687, n15_adj_3688, n18297, 
        n33886, n33859, n60, n70, n84, n17894, n18296, n18295, 
        n18294, n18293, n35093, n51, n73, n34209, n34170, n80, 
        n34156, n78, n29838, n79, n34323, n34251, n77, n29571, 
        n34293, n33917, n76, n34186, n75, n92, n34147, n85, 
        n33836, n82, n90, n94, n18279, n27503, n34133, n34108, 
        n33974, n81, n27502;
    wire [31:0]n93;
    
    wire n27501, n27528, n34510, n8_adj_3689;
    wire [7:0]n2236;
    
    wire n27527, n16648, n10_adj_3690, n16748, n6_adj_3691, n27526, 
        n27500, n17362, n37336, n39058, n5_adj_3692, n41878, n37337, 
        n37268, n37267, n34060, n29866, n30663, n33965, n16876, 
        n6_adj_3693, n18402, n18351, n17252, n33948, n16983, n1515, 
        n7_adj_3694, n27499, n16631, n10_adj_3695, n34054, n17307, 
        n34024, n16923, n10_adj_3696, n17040, n34302, n34320, n34173, 
        n1716, n16815, n6_adj_3697, n27525, n27524, n18350, n18349, 
        n18348, n18347, n17392, n27498, n14_adj_3698, n27523, n27497, 
        n34212, n17354, n10_adj_3699, n27522, n29832, n16086, n34087, 
        n34009, n12_adj_3700, n34275, n16668, n17256, n33932, n34257, 
        n18346, n17425, n35783, n35798, n18345, n18344, n18343, 
        n18342, n18341, n33911, n10_adj_3701, n18340, n34159, n10_adj_3702, 
        n33817, n12_adj_3703, n9_adj_3705, n224_c, n12_adj_3706, n34272, 
        n6_adj_3707, n10_adj_3708, n6_adj_3709, n12_adj_3710, n41872, 
        n6_adj_3711, n6_adj_3712, n35254, n6_adj_3713, n17259, n33758, 
        n16989, n34177, n34180, n34, n33908, n34278, n33880, n29836, 
        n15_adj_3714, n14163, n33961, n17128, n10_adj_3715, n33945, 
        n34266, n33993, n34057, n26_adj_3716, n6_adj_3717, n16066, 
        n16906, n34215, n16929, n6_adj_3718, n29810, n33795, n34326, 
        n34003, n16585, n34120, n14_adj_3719, n16_adj_3720, n34242, 
        n34006, n34111, n34245, n39105, n25608, n19_adj_3721, n39413, 
        n5_adj_3722, n37334, n41821, n37335, n37303, n37305, n41839, 
        n41833, n37304, n19_adj_3723, n39406, n5_adj_3724, n37331, 
        n41815, n37332, n37300, n37302, n41851, n41845, n37301, 
        n19_adj_3725, n41875, n8_adj_3726, n39401, n5_adj_3727, n37328, 
        n41809, n37329, n37297, n41866, n37299, n41869, n41860, 
        n41863, n41854, n41857, n41848, n41842, n37298, n4025, 
        n41836, n41830, n41824, n41827, n41818, n41812, n19_adj_3728, 
        n37325, n41743, n40612, n41803, n37326, n41881, n40616, 
        n41806;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n39029, n19_adj_3729, n6_adj_3730, n5_adj_3731, n37322, n41797, 
        n37323, n37294, n37296, n37295, n16102, n39026, n19_adj_3732, 
        n6_adj_3733, n5_adj_3734, n37319, n41791, n37320, n37291, 
        n37293, n41749, n41737, n37292, n19_adj_3735, n34043, n39382, 
        n17279, n6_adj_3736, n5_adj_3737, n37316, n41785, n37317, 
        n37288, n37290, n41761, n41755, n37289, n17265, n34199, 
        n13914, n4_adj_3738, n25610, n34236, n7_adj_3739, n41800, 
        n37194, n8_adj_3740, n41794, n38_adj_3741, n39_adj_3742, n220_c, 
        n24905, n37_adj_3743, n37190, n46, n37192, n37135, n35805, 
        n41788, n33747, n34572, n4_adj_3744, n14_adj_3745, n34455, 
        n5_adj_3746;
    wire [31:0]\FRAME_MATCHER.state_31__N_2435 ;
    
    wire n6_adj_3747, n41782, n34248, n34082, n34030, n34281, n8_adj_3748, 
        n17568, n10_adj_3749, n34305, n34051, n34114, n14_adj_3750, 
        n30703, n34284, n12_adj_3751, n16677, n6_adj_3752, n12_adj_3753, 
        n29879, n30316, n18_adj_3754, n20_adj_3755, n34233, n34036, 
        n34230, n16565, n15_adj_3756, n33875, n29828, n33883, n30665, 
        n34102, n33977, n17051, n6_adj_3757, n33833, n12_adj_3758, 
        n17085, n34079, n10_adj_3759, n29910, n34299, n33914, n29830, 
        n29848, n10_adj_3760, n1509, n33814, n17002, n34126, n10_adj_3761, 
        n34042, n17465, n34317, n16594, n33889, n33820, n41764, 
        n34066, n1664, n12_adj_3762, n54, n34162, n52, n34311, 
        n53, n51_adj_3763, n58, n56, n33999, n57, n33862, n55, 
        n64_adj_3764, n63_adj_3765, n35671, n12_adj_3766, n11, n30_adj_3767, 
        n28_adj_3768, n33935, n29_adj_3769, n17091, n17110, n27_adj_3770, 
        n17174, n12_adj_3771, n34183, n16661, n12_adj_3772, n14_adj_3773, 
        n33830, n34143, n15_adj_3774, n12_adj_3775, n34166, n6_adj_3776, 
        n41758, n16803, n1695, n14_adj_3777, n22_adj_3778, n24_adj_3779, 
        n23, n10_adj_3780, n12_adj_3781, n12_adj_3782, n34287, n6_adj_3783, 
        n8_adj_3784, n7_adj_3785, n41752, n16812, n41746, n41740, 
        n41734, n41728, n41731;
    
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18330));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18329));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18368));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18367));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18366));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18365));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n18364));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18363));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18362));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_32 (.CI(n27520), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27521));
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18361));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n18360));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n18359));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n18358));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18328));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18339));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n18278));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_7_lut (.I0(n6), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27495), .O(n33380)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n18277));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n18276));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n18275));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18338));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18337));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n33352), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut (.I0(n34254), .I1(\data_in_frame[14] [1]), .I2(n30655), 
            .I3(n6_adj_3566), .O(n30633));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_CARRY add_44_7 (.CI(n27495), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27496));
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n18274));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n18273));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n18272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n18271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n18270));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n18269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n18268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n18336));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n18267));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[6] [2]), .I1(n9), .I2(GND_net), 
            .I3(GND_net), .O(n16624));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_31_lut (.I0(n6), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27519), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n18266));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_6_lut (.I0(n6), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27494), .O(n33378)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n18265));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n18264));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n18263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n18262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n18261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n18260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n18290));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n18289));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n18288));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n18287));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_865 (.I0(n17338), .I1(\data_in_frame[6] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_865.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18400));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n18259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18399));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n18258));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n18257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18398));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n18256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n18255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n18254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18397));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n18286));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n18253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n18285));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n18252));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n18284));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18396));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18395));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18394));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18393));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18392));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18391));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18390));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18389));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18388));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18387));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18386));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18385));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18384));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_866 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33952));
    defparam i1_2_lut_adj_866.LUT_INIT = 16'h6666;
    SB_LUT4 i13882_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n18389));
    defparam i13882_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18383));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18382));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13883_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n18390));
    defparam i13883_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18381));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut (.I0(n33952), .I1(\data_in_frame[8] [7]), .I2(n16617), 
            .I3(n4_c), .O(n34224));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[13] [2]), .O(n33903));   // verilog/coms.v(70[16:41])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18380));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18379));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18378));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18377));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18376));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_867 (.I0(n16715), .I1(\data_in_frame[8] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n33986));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18375));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13884_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n18391));
    defparam i13884_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut (.I0(n33986), .I1(n34221), .I2(\data_in_frame[6] [3]), 
            .I3(GND_net), .O(n16796));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18374));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18373));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18372));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18371));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18370));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18369));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18335));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n18540));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n18541));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n18542));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n18543));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n18544));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n41916));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), .C(clk32MHz), 
            .E(VCC_net), .D(n18521));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n18427));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_868 (.I0(\data_in_frame[13] [3]), .I1(n17170), 
            .I2(n16789), .I3(GND_net), .O(n34308));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_868.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18428));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18429));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18430));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18431));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18432));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18433));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18419));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18420));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n18421));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n18422));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n18423));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n18424));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18408));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18409));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18327));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18326));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18325));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_869 (.I0(Kp_23__N_868), .I1(\data_in_frame[11] [2]), 
            .I2(\data_in_frame[6] [7]), .I3(\data_in_frame[7] [0]), .O(n34129));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18447));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18448));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18449));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18450));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n18251));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18324));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18323));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18445));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18446));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18322));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18443));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18444));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18321));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18441));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18442));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n18250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18439));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18440));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18437));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18438));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18434));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_870 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33856));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_870.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18435));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18436));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n18425));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n18426));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n18249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18410));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18411));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18412));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18413));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18414));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18415));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18416));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18417));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18418));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n18248));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_871 (.I0(\data_in_frame[4] [6]), .I1(n34129), .I2(GND_net), 
            .I3(GND_net), .O(n34260));   // verilog/coms.v(76[16:50])
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n18247));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n18246));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n18245));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18406));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18407));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18404));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18405));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n18244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n18243));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_31 (.CI(n27519), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27520));
    SB_CARRY add_44_6 (.CI(n27494), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27495));
    SB_LUT4 add_44_30_lut (.I0(n6), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27518), .O(n2_adj_3567)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_872 (.I0(n17114), .I1(\data_in_frame[6] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n34221));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_872.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n18283));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut (.I0(n34221), .I1(n34260), .I2(\data_in_frame[11] [1]), 
            .I3(n33856), .O(n12));   // verilog/coms.v(73[16:43])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n18242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n18241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n18240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n18239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n18238));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_5_lut (.I0(n6), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27493), .O(n33376)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n18237));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut (.I0(\data_in_frame[8] [6]), .I1(n12), .I2(n34308), 
            .I3(n16617), .O(n17187));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_873 (.I0(n33903), .I1(n34224), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3568));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n18236));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n18235));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18334));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_874 (.I0(n16624), .I1(\data_in_frame[8] [4]), .I2(n33986), 
            .I3(n6_adj_3568), .O(n16833));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n18234));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13885_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n18392));
    defparam i13885_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n18233));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18320));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n18232));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n18231));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n18282));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n18230));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n18229));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n18228));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_875 (.I0(n16833), .I1(n17187), .I2(\data_in_frame[15] [4]), 
            .I3(GND_net), .O(n17037));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_875.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n18227));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n18281));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_876 (.I0(Kp_23__N_1537), .I1(n34906), .I2(n30633), 
            .I3(n30661), .O(n34239));
    defparam i3_4_lut_adj_876.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n18280));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_877 (.I0(\data_in_frame[5] [0]), .I1(n29784), .I2(GND_net), 
            .I3(GND_net), .O(n29824));
    defparam i1_2_lut_adj_877.LUT_INIT = 16'h6666;
    SB_CARRY add_44_30 (.CI(n27518), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27519));
    SB_CARRY add_44_5 (.CI(n27493), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27494));
    SB_LUT4 i4_4_lut_adj_878 (.I0(\data_in_frame[11] [6]), .I1(n34039), 
            .I2(\data_in_frame[7] [2]), .I3(n30670), .O(n10));
    defparam i4_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[4] [6]), .I1(n10), .I2(n29900), 
            .I3(GND_net), .O(n33968));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_879 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[9] [4]), 
            .I2(n33968), .I3(n16937), .O(n10_adj_3569));
    defparam i4_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_880 (.I0(n35103), .I1(n10_adj_3569), .I2(\data_in_frame[9] [5]), 
            .I3(GND_net), .O(n30201));
    defparam i5_3_lut_adj_880.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n18226));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_3_lut (.I0(\data_out_frame[5] [0]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39361));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_881 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[11] [5]), 
            .I2(\data_in_frame[7] [3]), .I3(GND_net), .O(n14));   // verilog/coms.v(77[16:35])
    defparam i5_3_lut_adj_881.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i22_3_lut (.I0(n41767), .I1(n21), 
            .I2(byte_transmit_counter[2]), .I3(GND_net), .O(n22));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13886_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n18393));
    defparam i13886_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30965_4_lut (.I0(n5_c), .I1(\byte_transmit_counter[0] ), .I2(n38883), 
            .I3(n39361), .O(n37285));
    defparam i30965_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1_2_lut_3_lut (.I0(n16824), .I1(n30393), .I2(\data_in_frame[17] [6]), 
            .I3(GND_net), .O(n34136));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i30967_4_lut (.I0(n37285), .I1(n22), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37287));
    defparam i30967_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_44_29_lut (.I0(n6), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27517), .O(n32806)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut (.I0(n16617), .I1(n14), .I2(\data_in_frame[9] [4]), 
            .I3(\data_in_frame[6] [7]), .O(n16));   // verilog/coms.v(77[16:35])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n29824), .I1(n16), .I2(n12_adj_3570), .I3(\data_in_frame[9] [3]), 
            .O(n29915));   // verilog/coms.v(77[16:35])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_882 (.I0(n29915), .I1(n34329), .I2(\data_in_frame[13] [7]), 
            .I3(\data_in_frame[14] [0]), .O(n34090));
    defparam i3_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_883 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3] [2]), 
            .I2(n33843), .I3(n6_adj_3571), .O(n16937));   // verilog/coms.v(69[16:69])
    defparam i4_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_in_frame[7] [5]), .I1(n16937), .I2(GND_net), 
            .I3(GND_net), .O(n34227));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16964));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_886 (.I0(\data_in_frame[9] [7]), .I1(n33990), .I2(n17145), 
            .I3(\data_in_frame[6] [0]), .O(n12_adj_3572));
    defparam i5_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_887 (.I0(\data_in_frame[8] [1]), .I1(n12_adj_3572), 
            .I2(n34227), .I3(\data_in_frame[10] [2]), .O(n16093));
    defparam i6_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_4_lut (.I0(n6), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27492), .O(n33374)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13887_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18394));
    defparam i13887_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_888 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n34039));
    defparam i1_2_lut_adj_888.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_889 (.I0(n35103), .I1(\data_in_frame[9] [5]), .I2(\data_in_frame[11] [7]), 
            .I3(GND_net), .O(n33895));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_889.LUT_INIT = 16'h6969;
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1058));   // verilog/coms.v(83[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_890 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33852));
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_LUT4 i13888_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18395));
    defparam i13888_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13889_3_lut_4_lut (.I0(n8), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18396));
    defparam i13889_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [0]), 
            .I2(n6_adj_3573), .I3(\data_in_frame[1] [0]), .O(n29784));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_891 (.I0(n33990), .I1(\data_in_frame[8] [0]), .I2(n29784), 
            .I3(n34153), .O(n10_adj_3574));
    defparam i4_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_892 (.I0(n7), .I1(n10_adj_3574), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n29840));
    defparam i5_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_893 (.I0(n33852), .I1(\data_in_frame[12] [1]), 
            .I2(n16741), .I3(n33895), .O(n6_adj_3575));   // verilog/coms.v(83[17:70])
    defparam i1_4_lut_adj_893.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n18225));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18319));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n18224));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n18223));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n18222));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18318));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18317));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n18221));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n18220));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_894 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[9] [7]), .I3(n6_adj_3575), .O(n16952));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 i13810_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n18317));
    defparam i13810_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_895 (.I0(n24585), .I1(n16280), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n35752));   // verilog/coms.v(253[5:27])
    defparam i3_4_lut_adj_895.LUT_INIT = 16'hfeff;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n18219));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_29 (.CI(n27517), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27518));
    SB_CARRY add_44_4 (.CI(n27492), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27493));
    SB_LUT4 i1_4_lut_adj_896 (.I0(\data_in_frame[14] [4]), .I1(n16093), 
            .I2(n29840), .I3(n16964), .O(n29826));
    defparam i1_4_lut_adj_896.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n18218));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n18217));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_897 (.I0(\data_in_frame[14] [3]), .I1(n16952), 
            .I2(n29840), .I3(\data_in_frame[12] [2]), .O(n35995));
    defparam i3_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n18216));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n18215));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_898 (.I0(n35995), .I1(n29826), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1319));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n18214));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n18213));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n18212));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n18211));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n18210));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n18209));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n18208));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n18207));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13874_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n18381));
    defparam i13874_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n18206));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n18205));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n18204));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_899 (.I0(\data_in_frame[13] [5]), .I1(n34090), 
            .I2(n30610), .I3(GND_net), .O(n30677));
    defparam i2_3_lut_adj_899.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n18203));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n18202));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_900 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [2]), 
            .I2(n34090), .I3(GND_net), .O(n14_adj_3577));
    defparam i5_3_lut_adj_900.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n18201));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n18200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18316));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_901 (.I0(n34239), .I1(n17037), .I2(Kp_23__N_1319), 
            .I3(n34136), .O(n15));
    defparam i6_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i13875_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n18382));
    defparam i13875_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_28_lut (.I0(n6), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27516), .O(n32808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_28 (.CI(n27516), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27517));
    SB_LUT4 i1_4_lut_adj_902 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [3]), 
            .I2(n6_adj_3578), .I3(n34239), .O(n6_adj_3579));
    defparam i1_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_903 (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[14] [6]), 
            .I2(n33986), .I3(\data_in_frame[21] [6]), .O(n18));   // verilog/coms.v(71[16:42])
    defparam i7_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(\data_in_frame[19] [4]), .I1(n18), .I2(\data_in_frame[13] [0]), 
            .I3(n34218), .O(n20));   // verilog/coms.v(71[16:42])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[19] [3]), .I1(n29870), .I2(n34015), 
            .I3(GND_net), .O(n4_adj_3580));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_904 (.I0(n34203), .I1(\data_in_frame[10] [7]), 
            .I2(n33849), .I3(\data_in_frame[17] [2]), .O(n19_c));   // verilog/coms.v(71[16:42])
    defparam i8_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_905 (.I0(\data_in_frame[21] [4]), .I1(n19_c), .I2(n4_adj_3580), 
            .I3(n20), .O(n6_adj_3581));
    defparam i2_4_lut_adj_905.LUT_INIT = 16'hde7b;
    SB_LUT4 i1_4_lut_adj_906 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[21] [1]), 
            .I2(n34070), .I3(n30333), .O(n5_adj_3582));
    defparam i1_4_lut_adj_906.LUT_INIT = 16'hed7b;
    SB_LUT4 i1_rep_364_2_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42567));
    defparam i1_rep_364_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_907 (.I0(n33811), .I1(\data_in_frame[20] [4]), 
            .I2(n42567), .I3(n30633), .O(n12_adj_3583));
    defparam i5_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_908 (.I0(\data_in_frame[20] [0]), .I1(\data_in_frame[19] [7]), 
            .I2(n16833), .I3(GND_net), .O(n14_adj_3584));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_908.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n18199));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_909 (.I0(n34263), .I1(n17357), .I2(\data_in_frame[13] [4]), 
            .I3(n33823), .O(n15_adj_3585));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n18198));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n18197));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n18196));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n18195));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n18194));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_910 (.I0(n29818), .I1(\data_in_frame[18] [5]), 
            .I2(n30333), .I3(n34093), .O(n10_adj_3586));
    defparam i4_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n18193));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_911 (.I0(n29890), .I1(n34015), .I2(\data_in_frame[21] [3]), 
            .I3(GND_net), .O(n35078));
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_912 (.I0(n15), .I1(n34033), .I2(n14_adj_3577), 
            .I3(\data_in_frame[18] [0]), .O(n35005));
    defparam i8_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n18192));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18333));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_913 (.I0(\data_in_frame[18] [4]), .I1(n29928), 
            .I2(\data_in_frame[18] [3]), .I3(n6_adj_3587), .O(n35975));
    defparam i4_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18332));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_4_lut_adj_914 (.I0(n15_adj_3585), .I1(\data_in_frame[17] [4]), 
            .I2(n14_adj_3584), .I3(\data_in_frame[19] [6]), .O(n35214));   // verilog/coms.v(76[16:27])
    defparam i8_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_CARRY add_44_3 (.CI(n27491), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27492));
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n18191));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n18190));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_915 (.I0(n30633), .I1(n33801), .I2(n30720), .I3(\data_in_frame[20] [6]), 
            .O(n36127));
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_916 (.I0(\data_in_frame[18] [2]), .I1(n30655), 
            .I2(n33811), .I3(n6_adj_3579), .O(n36135));
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n18189));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n18188));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_917 (.I0(n35214), .I1(n35975), .I2(n35005), .I3(n35078), 
            .O(n22_adj_3588));
    defparam i9_4_lut_adj_917.LUT_INIT = 16'hffbf;
    SB_LUT4 i13876_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n18383));
    defparam i13876_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_918 (.I0(\data_in_frame[21] [5]), .I1(n34944), 
            .I2(n34105), .I3(\data_in_frame[19] [3]), .O(n15_adj_3589));
    defparam i2_4_lut_adj_918.LUT_INIT = 16'hb77b;
    SB_LUT4 i4_4_lut_adj_919 (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[19] [7]), 
            .I2(n34906), .I3(\data_in_frame[17] [7]), .O(n10_adj_3590));
    defparam i4_4_lut_adj_919.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_920 (.I0(n5_adj_3582), .I1(\data_in_frame[21] [7]), 
            .I2(n6_adj_3581), .I3(n34027), .O(n14_adj_3591));
    defparam i1_4_lut_adj_920.LUT_INIT = 16'hfefb;
    SB_LUT4 i6_4_lut_adj_921 (.I0(n30655), .I1(n12_adj_3583), .I2(\data_in_frame[16] [2]), 
            .I3(n34076), .O(n36136));
    defparam i6_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i13877_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n18384));
    defparam i13877_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut (.I0(n15_adj_3589), .I1(n22_adj_3588), .I2(n36135), 
            .I3(n36127), .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i13878_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n18385));
    defparam i13878_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30918_4_lut (.I0(n29890), .I1(n36064), .I2(n34070), .I3(\data_in_frame[21] [2]), 
            .O(n37172));
    defparam i30918_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i12_4_lut (.I0(n37172), .I1(n24), .I2(n36136), .I3(n14_adj_3591), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_4_lut_adj_922 (.I0(n7_adj_3592), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n24558), .I3(n47), .O(n36216));
    defparam i4_4_lut_adj_922.LUT_INIT = 16'hfeff;
    SB_LUT4 i13879_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n18386));
    defparam i13879_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n18187));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13880_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n18387));
    defparam i13880_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n18186));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n18185));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n18184));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18401));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20100_2_lut (.I0(n31), .I1(n24558), .I2(GND_net), .I3(GND_net), 
            .O(n24585));
    defparam i20100_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n18183));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13881_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n18388));
    defparam i13881_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_923 (.I0(n33790), .I1(n33678), .I2(n211), .I3(n6_adj_3593), 
            .O(n25604));
    defparam i4_4_lut_adj_923.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_924 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(n34012), .I3(\data_in_frame[3] [6]), .O(n17145));   // verilog/coms.v(83[17:28])
    defparam i1_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i13866_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18373));
    defparam i13866_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_925 (.I0(\data_in_frame[4] [1]), .I1(n34048), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[1] [5]), .O(n16715));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_926 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[5] [6]), .I3(n16778), .O(n7));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n18182));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n18181));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n18180));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3595));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_27_lut (.I0(n6), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27515), .O(n32810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n18179));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13867_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18374));
    defparam i13867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n18178));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_928 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[0] [0]), .I3(n6_adj_3595), .O(n16789));   // verilog/coms.v(68[16:27])
    defparam i4_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_929 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n4_adj_3596));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_929.LUT_INIT = 16'h9696;
    SB_LUT4 i13868_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18375));
    defparam i13868_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13869_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18376));
    defparam i13869_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_930 (.I0(\data_in_frame[4] [4]), .I1(n3_adj_3597), 
            .I2(n4_adj_3596), .I3(GND_net), .O(n17338));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_930.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n18177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n18176));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n18175));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n18174));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n18173));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n18172));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n18171));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_931 (.I0(\data_in_frame[4] [5]), .I1(n17155), .I2(n4_adj_3596), 
            .I3(GND_net), .O(n16617));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_931.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n18170));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n18169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n18168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n18167));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_932 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n4_adj_3598));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_932.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_933 (.I0(n4_adj_3598), .I1(n34099), .I2(GND_net), 
            .I3(GND_net), .O(n30670));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_in_frame[5] [1]), .I1(n29852), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3599));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n18166));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_27 (.CI(n27515), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27516));
    SB_LUT4 i4_4_lut_adj_935 (.I0(Kp_23__N_833), .I1(\data_in_frame[1] [0]), 
            .I2(n33843), .I3(n6_adj_3599), .O(n33943));   // verilog/coms.v(68[16:69])
    defparam i4_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n18165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n18164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n18163));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13870_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18377));
    defparam i13870_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_936 (.I0(\data_in_frame[5] [5]), .I1(n33792), .I2(\data_in_frame[3] [3]), 
            .I3(\data_in_frame[3] [4]), .O(n16741));   // verilog/coms.v(71[16:34])
    defparam i3_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_2_lut (.I0(n6), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n33352)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34048));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_938 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3600));
    defparam i6_4_lut_adj_938.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_939 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16778));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_940 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_940.LUT_INIT = 16'hfffd;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n18162));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_941 (.I0(n17), .I1(\data_in[1] [6]), .I2(n16_adj_3600), 
            .I3(\data_in[3] [7]), .O(n16397));
    defparam i9_4_lut_adj_941.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n18161));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_942 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n16295), .O(n16_adj_3601));
    defparam i6_4_lut_adj_942.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_943 (.I0(n16397), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_3602));
    defparam i7_4_lut_adj_943.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33804));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_945 (.I0(n17_adj_3602), .I1(\data_in[3] [5]), .I2(n16_adj_3601), 
            .I3(\data_in[3] [3]), .O(n63_c));
    defparam i9_4_lut_adj_945.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n18160));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_946 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n16394), .I3(\data_in[1] [0]), .O(n18_adj_3603));
    defparam i7_4_lut_adj_946.LUT_INIT = 16'hfffd;
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n18159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n18158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n18157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n18156));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_947 (.I0(\data_in[1] [4]), .I1(n18_adj_3603), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [3]), .O(n20_adj_3604));
    defparam i9_4_lut_adj_947.LUT_INIT = 16'hfffd;
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n18155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n18154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n18153));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n18152));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n18151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n18150));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n33843));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n18149));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10_4_lut (.I0(n15_adj_3605), .I1(n20_adj_3604), .I2(n16397), 
            .I3(\data_in[0] [6]), .O(n63_adj_3606));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i20195_4_lut (.I0(n10_adj_3607), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n16466), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i20195_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i2_3_lut_adj_949 (.I0(\FRAME_MATCHER.state [1]), .I1(n16406), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n16420));   // verilog/coms.v(161[5:29])
    defparam i2_3_lut_adj_949.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33898));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n34290));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n34012));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_953 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [7]), 
            .I2(n33898), .I3(n6_adj_3608), .O(Kp_23__N_833));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33929));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [0]), 
            .I2(n3_adj_3597), .I3(n18_adj_3609), .O(n30));   // verilog/coms.v(166[9:87])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_955 (.I0(\data_in_frame[3] [1]), .I1(Kp_23__N_868), 
            .I2(n33898), .I3(n33807), .O(n28));   // verilog/coms.v(166[9:87])
    defparam i11_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_956 (.I0(\data_in_frame[2] [3]), .I1(n33843), 
            .I2(\data_in_frame[2] [6]), .I3(n33804), .O(n29));   // verilog/coms.v(166[9:87])
    defparam i12_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_957 (.I0(n16778), .I1(n34290), .I2(n34048), 
            .I3(n34123), .O(n27));   // verilog/coms.v(166[9:87])
    defparam i10_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n29852));   // verilog/coms.v(166[9:87])
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_958 (.I0(n29852), .I1(\data_in_frame[3] [0]), .I2(n33929), 
            .I3(Kp_23__N_833), .O(n34099));   // verilog/coms.v(68[16:69])
    defparam i3_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_959 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n17155));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_960 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n4_adj_3610));
    defparam i1_3_lut_adj_960.LUT_INIT = 16'heaea;
    SB_LUT4 i32536_2_lut (.I0(byte_transmit_counter[2]), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n38883));
    defparam i32536_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n18148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n18147));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n18146));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_961 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3611));
    defparam i6_4_lut_adj_961.LUT_INIT = 16'h8000;
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n18145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n18144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n18143));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_962 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3612));   // verilog/coms.v(232[13:35])
    defparam i6_4_lut_adj_962.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_963 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13));
    defparam i5_4_lut_adj_963.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_964 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3613));   // verilog/coms.v(232[13:35])
    defparam i5_4_lut_adj_964.LUT_INIT = 16'hfffe;
    SB_LUT4 i20074_4_lut (.I0(n13_adj_3613), .I1(n13), .I2(n14_adj_3612), 
            .I3(n14_adj_3611), .O(n24558));
    defparam i20074_4_lut.LUT_INIT = 16'h32fa;
    SB_LUT4 equal_1134_i15_2_lut (.I0(Kp_23__N_868), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3614));   // verilog/coms.v(230[9:81])
    defparam equal_1134_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_1134_i16_2_lut (.I0(Kp_23__N_871), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3615));   // verilog/coms.v(230[9:81])
    defparam equal_1134_i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_965 (.I0(n30692), .I1(n16741), .I2(n15_adj_3614), 
            .I3(n33943), .O(n28_adj_3616));   // verilog/coms.v(230[9:81])
    defparam i12_4_lut_adj_965.LUT_INIT = 16'hfffb;
    SB_LUT4 i10_4_lut_adj_966 (.I0(n16617), .I1(n17114), .I2(n16_adj_3615), 
            .I3(n17338), .O(n26));   // verilog/coms.v(230[9:81])
    defparam i10_4_lut_adj_966.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_967 (.I0(n16937), .I1(n9), .I2(n17141), .I3(n29784), 
            .O(n27_adj_3617));   // verilog/coms.v(230[9:81])
    defparam i11_4_lut_adj_967.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_968 (.I0(n16789), .I1(n7), .I2(n16715), .I3(n17145), 
            .O(n25));   // verilog/coms.v(230[9:81])
    defparam i9_4_lut_adj_968.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27_adj_3617), .I2(n26), .I3(n28_adj_3616), 
            .O(n31_adj_3618));   // verilog/coms.v(230[9:81])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20076_2_lut (.I0(n31_adj_3618), .I1(n24558), .I2(GND_net), 
            .I3(GND_net), .O(n24560));
    defparam i20076_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_969 (.I0(n25604), .I1(n24585), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [2]), .O(n5_adj_3619));
    defparam i1_4_lut_adj_969.LUT_INIT = 16'haeaa;
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n18142));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_970 (.I0(n5_adj_3619), .I1(n13888), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n4_adj_3620), .O(n19473));
    defparam i3_4_lut_adj_970.LUT_INIT = 16'hbfbb;
    SB_LUT4 i3_4_lut_adj_971 (.I0(byte_transmit_counter[7]), .I1(n25566), 
            .I2(byte_transmit_counter[6]), .I3(byte_transmit_counter[5]), 
            .O(n25598));
    defparam i3_4_lut_adj_971.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n18141));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13871_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18378));
    defparam i13871_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_26_lut (.I0(n6), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27514), .O(n32816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n27491));
    SB_CARRY add_44_26 (.CI(n27514), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27515));
    SB_LUT4 add_44_25_lut (.I0(n6), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27513), .O(n32824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13872_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18379));
    defparam i13872_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13873_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18380));
    defparam i13873_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14970_3_lut (.I0(byte_transmit_counter[3]), .I1(n38993), .I2(n19473), 
            .I3(GND_net), .O(n18540));
    defparam i14970_3_lut.LUT_INIT = 16'hacac;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n18140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n18139));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n18138));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n18137));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n18136));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n18135));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n18134));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_25 (.CI(n27513), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27514));
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n18133));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_24_lut (.I0(n6), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27512), .O(n32832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n18132));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n18131));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut_adj_972 (.I0(n35990), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n16406), .O(n4_adj_3621));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h55d5;
    SB_LUT4 i13811_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n18318));
    defparam i13811_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_3_lut (.I0(n39102), .I1(\byte_transmit_counter[1] ), .I2(n19473), 
            .I3(GND_net), .O(n32898));   // verilog/coms.v(100[12:33])
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n18130));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14981_3_lut (.I0(n19484), .I1(n19473), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n18020));   // verilog/coms.v(100[12:33])
    defparam i14981_3_lut.LUT_INIT = 16'he2e2;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(\FRAME_MATCHER.i [6]), .I3(\FRAME_MATCHER.i [24]), .O(n42));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_973 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [27]), .O(n40));
    defparam i15_4_lut_adj_973.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_974 (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut_adj_974.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n18129));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n18128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n18127));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY add_44_24 (.CI(n27512), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27513));
    SB_LUT4 add_44_23_lut (.I0(n6), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27511), .O(n32846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [19]), .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48), .I2(n37), .I3(n38), .O(n16466));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n18126));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n18125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n18124));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_975 (.I0(\FRAME_MATCHER.state [1]), .I1(n16406), 
            .I2(GND_net), .I3(GND_net), .O(n16403));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_adj_975.LUT_INIT = 16'heeee;
    SB_CARRY add_44_23 (.CI(n27511), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27512));
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n18123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n18122));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n18121));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18403));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_976 (.I0(\data_in[0] [4]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [7]), .I3(\data_in[3] [4]), .O(n10_adj_3622));
    defparam i4_4_lut_adj_976.LUT_INIT = 16'hdfff;
    SB_LUT4 i5_3_lut_adj_977 (.I0(\data_in[1] [1]), .I1(n10_adj_3622), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n16469));
    defparam i5_3_lut_adj_977.LUT_INIT = 16'hefef;
    SB_LUT4 i30894_3_lut (.I0(\data_in[3] [0]), .I1(\data_in[2] [2]), .I2(\data_in[1] [5]), 
            .I3(GND_net), .O(n37145));
    defparam i30894_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_978 (.I0(\data_in[1] [0]), .I1(\data_in[0] [6]), 
            .I2(\data_in[2] [4]), .I3(\data_in[0] [3]), .O(n15_adj_3623));
    defparam i6_4_lut_adj_978.LUT_INIT = 16'hfdff;
    SB_LUT4 i8_4_lut_adj_979 (.I0(n15_adj_3623), .I1(\data_in[1] [4]), .I2(n37145), 
            .I3(n16469), .O(n16295));
    defparam i8_4_lut_adj_979.LUT_INIT = 16'hffef;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3624));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_980 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3625));
    defparam i6_4_lut_adj_980.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_981 (.I0(\data_in[3] [6]), .I1(n14_adj_3625), .I2(n10_adj_3624), 
            .I3(\data_in[2] [1]), .O(n16394));
    defparam i7_4_lut_adj_981.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_982 (.I0(n16394), .I1(\data_in[1] [3]), .I2(n16295), 
            .I3(\data_in[1] [2]), .O(n20_adj_3626));
    defparam i8_4_lut_adj_982.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n18120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n18119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n18118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0] [4]), .C(clk32MHz), 
           .D(n18117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0] [3]), .C(clk32MHz), 
           .D(n18116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0] [2]), .C(clk32MHz), 
           .D(n18115));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_983 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_3627));
    defparam i7_4_lut_adj_983.LUT_INIT = 16'hfeff;
    SB_LUT4 i30924_4_lut (.I0(\data_in[3] [2]), .I1(\data_in[0] [5]), .I2(\data_in[2] [0]), 
            .I3(\data_in[2] [5]), .O(n37178));
    defparam i30924_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_984 (.I0(n37178), .I1(n19_adj_3627), .I2(n20_adj_3626), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut_adj_984.LUT_INIT = 16'hfdfd;
    SB_LUT4 i20253_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_3606), 
            .I2(n63_c), .I3(GND_net), .O(n123));   // verilog/coms.v(139[4] 142[7])
    defparam i20253_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_362_Select_2_i5_4_lut (.I0(n123), .I1(n16404), .I2(n2857), 
            .I3(n63), .O(n5));
    defparam select_362_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 add_44_22_lut (.I0(n6), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27510), .O(n32860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n18114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n18113));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i20256_rep_385_2_lut (.I0(n123), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n42588));   // verilog/coms.v(143[4] 146[7])
    defparam i20256_rep_385_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_44_22 (.CI(n27510), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27511));
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n18112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n18111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n18110));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n18109));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n18108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n18107));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i30887_2_lut_4_lut (.I0(n16256), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3610), .I3(n16405), .O(n37137));   // verilog/coms.v(157[9:60])
    defparam i30887_2_lut_4_lut.LUT_INIT = 16'hff32;
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n18106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n18105));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5529_2_lut_4_lut (.I0(n16256), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3610), .I3(n63), .O(n9783));   // verilog/coms.v(157[9:60])
    defparam i5529_2_lut_4_lut.LUT_INIT = 16'hcd00;
    SB_LUT4 add_44_21_lut (.I0(n6), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27509), .O(n32874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n18104));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n18103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n18102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n18101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n18100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n18099));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n18098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n18097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n18096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n18095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n18094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n18093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n18092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n18091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n18090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n18089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n18088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n18087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n18086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n18085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n18084));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n18083));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n18082));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n18081));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n18080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n18079));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n18078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n18077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n18075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n18074));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_21 (.CI(n27509), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27510));
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n18073));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n18072));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n18071));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n18070));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n18069));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n18068));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n18067));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n18066));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n18065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n18064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n18063));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n18062));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n18061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n18060));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n18059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n18058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n18057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n18056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n18055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n18054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n18053));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14974_3_lut (.I0(byte_transmit_counter[7]), .I1(n38991), .I2(n19473), 
            .I3(GND_net), .O(n18544));
    defparam i14974_3_lut.LUT_INIT = 16'hacac;
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n18020));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), .C(clk32MHz), 
           .D(n32898));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5564_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9818));
    defparam i5564_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_44_20_lut (.I0(n6), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27508), .O(n32892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n17974));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_20 (.CI(n27508), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27509));
    SB_LUT4 add_44_19_lut (.I0(n6), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27507), .O(n32938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_19 (.CI(n27507), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27508));
    SB_LUT4 i14972_3_lut (.I0(byte_transmit_counter[5]), .I1(n38992), .I2(n19473), 
            .I3(GND_net), .O(n18542));
    defparam i14972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_44_18_lut (.I0(n6), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27506), .O(n32956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n17973));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n17972));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n17971));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n17970));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n17969));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n17968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n17967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n17966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n17965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n17964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n17963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n17962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n17961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n17960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n17959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n17958));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n17957));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n17956));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n17955));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n17954));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n17953));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n17952));   // verilog/coms.v(126[12] 289[6])
    SB_DFF LED_3230 (.Q(LED_c), .C(clk32MHz), .D(n34492));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_18 (.CI(n27506), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27507));
    SB_LUT4 i2027_3_lut (.I0(n31), .I1(n31_adj_3618), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n13746));
    defparam i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_4_lut_adj_985 (.I0(n24558), .I1(\FRAME_MATCHER.state_31__N_2467 [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n13746), .O(n6_adj_3630));
    defparam i17_4_lut_adj_985.LUT_INIT = 16'h0c5c;
    SB_LUT4 add_44_17_lut (.I0(n6), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27505), .O(n32978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2020_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3631));
    defparam i2020_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14976_3_lut (.I0(byte_transmit_counter[4]), .I1(n38994), .I2(n19473), 
            .I3(GND_net), .O(n18541));
    defparam i14976_3_lut.LUT_INIT = 16'hacac;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n33372), .S(n3_adj_3632));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i15_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47));
    defparam i15_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n18292));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_17 (.CI(n27505), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27506));
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18315));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18314));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18313));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18312));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18311));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n18310));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n18309));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n18308));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n18307));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n33374), .S(n3_adj_3633));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(n29826), .I1(n35995), .I2(n34018), 
            .I3(\data_in_frame[16] [0]), .O(n34140));
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n33376), .S(n3_adj_3634));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n33378), .S(n3_adj_3635));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n33380), .S(n3_adj_3636));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n33242), .S(n3_adj_3637));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n33192), .S(n3_adj_3638));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n33110), .S(n3_adj_3639));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n33090), .S(n3_adj_3640));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n33076), .S(n3_adj_3641));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n33054), .S(n3_adj_3642));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n33036), .S(n3_adj_3643));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n33018), .S(n3_adj_3644));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n33004), .S(n3_adj_3645));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n32978), .S(n3_adj_3646));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n32956), .S(n3_adj_3647));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n32938), .S(n3_adj_3648));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n32892), .S(n3_adj_3649));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n32874), .S(n3_adj_3650));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n32860), .S(n3_adj_3651));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n32846), .S(n3_adj_3652));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n32832), .S(n3_adj_3653));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n32824), .S(n3_adj_3654));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n32816), .S(n3_adj_3655));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n32810), .S(n3_adj_3656));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n32808), .S(n3_adj_3657));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n32806), .S(n3_adj_3658));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3567), .S(n3_adj_3659));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3660));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3661), .S(n3_adj_3662));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3663), .S(n3_adj_3664));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n17572), .D(n34115));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21]_c [1]), .C(clk32MHz), 
            .E(n17572), .D(n36123));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21]_c [2]), .C(clk32MHz), 
            .E(n17572), .D(n35111));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21]_c [3]), .C(clk32MHz), 
            .E(n17572), .D(n34814));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21]_c [4]), .C(clk32MHz), 
            .E(n17572), .D(n34884));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21]_c [5]), .C(clk32MHz), 
            .E(n17572), .D(n35096));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21]_c [6]), .C(clk32MHz), 
            .E(n17572), .D(n34928));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21]_c [7]), .C(clk32MHz), 
            .E(n17572), .D(n35199));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n17572), .D(n35420));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22]_c [1]), .C(clk32MHz), 
            .E(n17572), .D(n34307));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22]_c [2]), .C(clk32MHz), 
            .E(n17572), .D(n35129));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22]_c [3]), .C(clk32MHz), 
            .E(n17572), .D(n34031));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22]_c [4]), .C(clk32MHz), 
            .E(n17572), .D(n33912));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22]_c [5]), .C(clk32MHz), 
            .E(n17572), .D(n34046));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22]_c [6]), .C(clk32MHz), 
            .E(n17572), .D(n34084));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22]_c [7]), .C(clk32MHz), 
            .E(n17572), .D(n34249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n18306));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n33126), .S(n42066));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n33140), .S(n33382));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n33296), .S(n33142));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n33300), .S(n33190));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n33304), .S(n33188));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n33292), .S(n33198));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n33308), .S(n33186));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n33312), .S(n33184));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n33316), .S(n33182));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n33320), .S(n33180));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n33284), .S(n33218));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n64), .S(n33134));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n24574), .S(n25301));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_3665), .S(n8_adj_3666));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n33324), .S(n33174));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n7_adj_3667), .S(n8_adj_3668));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_3669), .S(n8_adj_3670));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n33328), .S(n33172));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n33332), .S(n33170));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n33336), .S(n33168));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n33340), .S(n33166));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_3671), .S(n8_adj_3672));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n33288), .S(n33200));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n33344), .S(n33164));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n33348), .S(n33162));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_3673), .S(n8_adj_3674));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n33258), .S(n33228));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n33262), .S(n33160));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n33274), .S(n33158));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_3675), .S(n8_adj_3676));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_986 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [8]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n10_adj_3677));
    defparam i4_4_lut_adj_986.LUT_INIT = 16'hfffe;
    SB_LUT4 i28246_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16410));
    defparam i28246_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_44_3_lut (.I0(n6), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27491), .O(n33372)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n18305));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_987 (.I0(\FRAME_MATCHER.state [11]), .I1(n10_adj_3677), 
            .I2(\FRAME_MATCHER.state [12]), .I3(GND_net), .O(n33790));
    defparam i5_3_lut_adj_987.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n18304));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18357));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_337_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_337_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n18303));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3227 (.Q(\r_SM_Main_2__N_3298[0] ), .C(clk32MHz), 
            .D(n39174), .R(n34543));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n18302));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[16] [3]), .I1(n30661), 
            .I2(GND_net), .I3(GND_net), .O(n29928));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h9999;
    SB_LUT4 add_44_16_lut (.I0(n6), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27504), .O(n33004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i35357_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3298[0] ), 
            .I2(n25598), .I3(GND_net), .O(tx_transmit_N_3190));
    defparam i35357_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_adj_989 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34033));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_989.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_990 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[16] [1]), .I3(n34033), .O(n10_adj_3678));
    defparam i4_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18356));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18355));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18354));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18353));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18352));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n18301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n18300));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n18299));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n18298));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18331));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n33144));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_2_lut (.I0(\FRAME_MATCHER.state [25]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3679));   // verilog/coms.v(206[5:16])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_991 (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [28]), 
            .I2(\FRAME_MATCHER.state [19]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n22_adj_3680));   // verilog/coms.v(206[5:16])
    defparam i9_4_lut_adj_991.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [17]), 
            .I2(\FRAME_MATCHER.state [16]), .I3(GND_net), .O(n20_adj_3681));   // verilog/coms.v(206[5:16])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_992 (.I0(\FRAME_MATCHER.state [21]), .I1(n22_adj_3680), 
            .I2(n16_adj_3679), .I3(\FRAME_MATCHER.state [22]), .O(n24_adj_3682));   // verilog/coms.v(206[5:16])
    defparam i11_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_993 (.I0(\FRAME_MATCHER.state [20]), .I1(n24_adj_3682), 
            .I2(n20_adj_3681), .I3(\FRAME_MATCHER.state [29]), .O(n33678));   // verilog/coms.v(206[5:16])
    defparam i12_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_994 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [6]), 
            .I2(\FRAME_MATCHER.state [7]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n33788));
    defparam i3_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_995 (.I0(\data_in_frame[16] [0]), .I1(n10_adj_3678), 
            .I2(n16824), .I3(GND_net), .O(n33811));
    defparam i5_3_lut_adj_995.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_996 (.I0(n30720), .I1(n33971), .I2(\data_in_frame[19] [0]), 
            .I3(\data_in_frame[16] [4]), .O(n29818));
    defparam i3_4_lut_adj_996.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_997 (.I0(Kp_23__N_1444), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[15] [3]), .I3(GND_net), .O(n33823));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_997.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17896));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_2_lut (.I0(\data_in_frame[13] [5]), .I1(n16833), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_3683));   // verilog/coms.v(72[16:43])
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_998 (.I0(n33823), .I1(n30610), .I2(\data_in_frame[15] [6]), 
            .I3(\data_in_frame[17] [5]), .O(n13_adj_3684));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n18291));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_999 (.I0(n13_adj_3684), .I1(n30710), .I2(n12_adj_3683), 
            .I3(\data_in_frame[18] [0]), .O(n34206));   // verilog/coms.v(72[16:43])
    defparam i7_4_lut_adj_999.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[14] [7]), .I3(\data_in_frame[17] [3]), .O(n33983));
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(n17155), .O(Kp_23__N_868));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1001 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(n34099), .O(Kp_23__N_871));
    defparam i1_2_lut_4_lut_adj_1001.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1328));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1002 (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [27]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(GND_net), .O(n211));
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1003 (.I0(n211), .I1(n33788), .I2(n33678), .I3(n6_adj_3685), 
            .O(n16285));   // verilog/coms.v(206[5:16])
    defparam i4_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1004 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n16285), .I3(GND_net), .O(n16406));   // verilog/coms.v(244[5:25])
    defparam i2_3_lut_adj_1004.LUT_INIT = 16'hfbfb;
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 equal_1134_i9_3_lut_4_lut (.I0(\data_in_frame[3] [6]), .I1(n33898), 
            .I2(\data_in_frame[4] [0]), .I3(\data_in_frame[3] [7]), .O(n9));   // verilog/coms.v(83[17:28])
    defparam equal_1134_i9_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34021));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1006 (.I0(\data_in_frame[10] [5]), .I1(n33940), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[8] [5]), .O(n12_adj_3686));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1007 (.I0(n17170), .I1(n12_adj_3686), .I2(n34203), 
            .I3(\data_in_frame[10] [6]), .O(Kp_23__N_1444));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1008 (.I0(\data_in_frame[19] [4]), .I1(n29870), 
            .I2(n34218), .I3(n33983), .O(n34105));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1009 (.I0(Kp_23__N_1444), .I1(\data_in_frame[17] [3]), 
            .I2(\data_in_frame[19] [6]), .I3(GND_net), .O(n14_adj_3687));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1010 (.I0(\data_in_frame[19] [5]), .I1(n33849), 
            .I2(n17037), .I3(n17357), .O(n15_adj_3688));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_CARRY add_44_16 (.CI(n27504), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27505));
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n18297));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17895));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_4_lut_adj_1011 (.I0(n15_adj_3688), .I1(n34021), .I2(n14_adj_3687), 
            .I3(n33886), .O(n34027));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i12_3_lut (.I0(\data_in_frame[18] [2]), .I1(n33859), .I2(\data_in_frame[18] [3]), 
            .I3(GND_net), .O(n60));
    defparam i12_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i22_2_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n70));
    defparam i22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36_4_lut (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[10] [1]), .I3(n16964), .O(n84));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17894));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17893));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n18296));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n18295));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n18294));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n18293));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n17141), .I1(n29900), .I2(n16937), 
            .I3(GND_net), .O(n35093));
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [7]), 
            .I2(n34015), .I3(GND_net), .O(n51));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(n34027), .I1(n29890), .I2(n33801), .I3(n34105), 
            .O(n73));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(n34308), .I1(n34209), .I2(n34263), .I3(n34170), 
            .O(n80));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n34156), .I1(n60), .I2(\data_in_frame[17] [7]), 
            .I3(Kp_23__N_1319), .O(n78));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(\data_in_frame[5] [0]), .I1(n29838), .I2(\data_in_frame[14] [3]), 
            .I3(n34329), .O(n79));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n35093), .I1(n34323), .I2(\data_in_frame[14] [4]), 
            .I3(n34251), .O(n77));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n29571), .I1(n34129), .I2(n34293), .I3(n33917), 
            .O(n76));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(n34140), .I1(Kp_23__N_1328), .I2(n34186), .I3(n33983), 
            .O(n75));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i44_4_lut (.I0(n77), .I1(n79), .I2(n78), .I3(n80), .O(n92));
    defparam i44_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i37_4_lut (.I0(n73), .I1(n51), .I2(n34147), .I3(n34206), 
            .O(n85));
    defparam i37_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34_4_lut (.I0(n33952), .I1(n33836), .I2(n33903), .I3(\data_in_frame[18] [1]), 
            .O(n82));
    defparam i34_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i42_4_lut (.I0(\data_in_frame[13] [0]), .I1(n84), .I2(n70), 
            .I3(n30633), .O(n90));
    defparam i42_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i46_4_lut (.I0(n85), .I1(n92), .I2(n75), .I3(n76), .O(n94));
    defparam i46_4_lut.LUT_INIT = 16'h6996;
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n17793));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17791));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n17892));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n18279));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_15_lut (.I0(n6), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27503), .O(n33018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33_4_lut (.I0(n34133), .I1(n34021), .I2(n34108), .I3(n33974), 
            .O(n81));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_44_15 (.CI(n27503), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27504));
    SB_LUT4 add_44_14_lut (.I0(n6), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27502), .O(n33036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_14 (.CI(n27502), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27503));
    SB_LUT4 i2_2_lut_3_lut (.I0(n63_c), .I1(n63_adj_3606), .I2(n63), .I3(GND_net), 
            .O(n11748));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i20735_2_lut_3_lut (.I0(n63_c), .I1(n63_adj_3606), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n93[1]));
    defparam i20735_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_44_13_lut (.I0(n6), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27501), .O(n33054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_626_9_lut (.I0(n9818), .I1(byte_transmit_counter[7]), .I2(GND_net), 
            .I3(n27528), .O(n38991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i47_4_lut (.I0(n81), .I1(n94), .I2(n90), .I3(n82), .O(n30333));
    defparam i47_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20799_1_lut (.I0(n34510), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n6));
    defparam i20799_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13850_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18357));
    defparam i13850_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_626_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n27527), .O(n2236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13851_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n18358));
    defparam i13851_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_13 (.CI(n27501), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27502));
    SB_LUT4 i13852_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n18359));
    defparam i13852_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13853_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n18360));
    defparam i13853_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13854_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18361));
    defparam i13854_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_626_8 (.CI(n27527), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n27528));
    SB_LUT4 i4_4_lut_adj_1013 (.I0(n34093), .I1(\data_in_frame[14] [6]), 
            .I2(n16648), .I3(n34251), .O(n10_adj_3690));
    defparam i4_4_lut_adj_1013.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(\data_in_frame[19] [1]), .I1(n16748), 
            .I2(n10_adj_3690), .I3(\data_in_frame[16] [7]), .O(n29890));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'h9669;
    SB_LUT4 i13855_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18362));
    defparam i13855_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(n7), .I1(\data_in_frame[7] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3691));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 add_626_7_lut (.I0(n9818), .I1(byte_transmit_counter[5]), .I2(GND_net), 
            .I3(n27526), .O(n38992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_12_lut (.I0(n6), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27500), .O(n33076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1016 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[12] [5]), 
            .I2(n17362), .I3(n6_adj_3691), .O(n34170));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i13856_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18363));
    defparam i13856_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[4] [3]), .I3(n33804), .O(n17114));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13857_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n18364));
    defparam i13857_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34323));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i31016_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n37336));
    defparam i31016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n39058), .I2(n5_adj_3692), .I3(byte_transmit_counter[2]), 
            .O(n41878));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i31017_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n37337));
    defparam i31017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30948_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n37268));
    defparam i30948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30947_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n37267));
    defparam i30947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1018 (.I0(\data_out_frame[14] [4]), .I1(n34060), 
            .I2(n29866), .I3(GND_net), .O(n30663));
    defparam i1_2_lut_3_lut_adj_1018.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1019 (.I0(\data_out_frame[14] [4]), .I1(n34060), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n33965));
    defparam i1_2_lut_3_lut_adj_1019.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1020 (.I0(n16876), .I1(\data_in_frame[10] [3]), 
            .I2(n34170), .I3(n6_adj_3693), .O(n16648));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1021 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n3_adj_3597));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18402));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1022 (.I0(n16648), .I1(n34323), .I2(\data_in_frame[17] [4]), 
            .I3(GND_net), .O(n33849));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1022.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18351));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_2_lut_4_lut (.I0(n17252), .I1(n33948), .I2(n16983), .I3(n1515), 
            .O(n7_adj_3694));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_44_12 (.CI(n27500), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27501));
    SB_LUT4 add_44_11_lut (.I0(n6), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27499), .O(n33090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1023 (.I0(n17338), .I1(n16631), .I2(\data_in_frame[13] [1]), 
            .I3(n34224), .O(n10_adj_3695));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_CARRY add_626_7 (.CI(n27526), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n27527));
    SB_LUT4 i1_2_lut_4_lut_adj_1024 (.I0(n17252), .I1(n33948), .I2(n16983), 
            .I3(\data_out_frame[13] [4]), .O(n34054));
    defparam i1_2_lut_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1025 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(n17307), .I3(n34024), .O(n16923));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1026 (.I0(\data_in_frame[6] [3]), .I1(n10_adj_3695), 
            .I2(\data_in_frame[13] [2]), .I3(GND_net), .O(n34203));   // verilog/coms.v(72[16:43])
    defparam i5_3_lut_adj_1026.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(n10_adj_3696), .O(n17040));   // verilog/coms.v(71[16:34])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1027 (.I0(n34302), .I1(n34320), .I2(\data_out_frame[12] [0]), 
            .I3(n34173), .O(n1716));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_CARRY add_44_11 (.CI(n27499), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27500));
    SB_LUT4 i4_4_lut_adj_1028 (.I0(n16815), .I1(\data_in_frame[12] [7]), 
            .I2(n16796), .I3(n6_adj_3697), .O(n33886));
    defparam i4_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 add_626_6_lut (.I0(n9818), .I1(byte_transmit_counter[4]), .I2(GND_net), 
            .I3(n27525), .O(n38994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_626_6 (.CI(n27525), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n27526));
    SB_LUT4 add_626_5_lut (.I0(n9818), .I1(byte_transmit_counter[3]), .I2(GND_net), 
            .I3(n27524), .O(n38993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18350));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18348));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18347));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1029 (.I0(n34302), .I1(n34320), .I2(\data_out_frame[12] [1]), 
            .I3(GND_net), .O(n17392));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_1029.LUT_INIT = 16'h9696;
    SB_LUT4 add_44_10_lut (.I0(n6), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27498), .O(n33110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_626_5 (.CI(n27524), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n27525));
    SB_CARRY add_44_10 (.CI(n27498), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27499));
    SB_LUT4 i1_2_lut_3_lut_adj_1030 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(\data_out_frame[18] [2]), .I3(GND_net), .O(n14_adj_3698));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 add_626_4_lut (.I0(n9818), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(n27523), .O(n19484)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_626_4 (.CI(n27523), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n27524));
    SB_LUT4 add_44_9_lut (.I0(n6), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27497), .O(n33192)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34212));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1032 (.I0(\data_in_frame[19] [2]), .I1(n34212), 
            .I2(\data_in_frame[14] [7]), .I3(n17354), .O(n10_adj_3699));
    defparam i4_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 add_626_3_lut (.I0(n9818), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n27522), .O(n39102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_adj_1033 (.I0(n33971), .I1(n10_adj_3699), .I2(\data_in_frame[17] [0]), 
            .I3(GND_net), .O(n34015));
    defparam i5_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1034 (.I0(\data_out_frame[15] [7]), .I1(n29832), 
            .I2(n16086), .I3(GND_net), .O(n34087));
    defparam i1_2_lut_3_lut_adj_1034.LUT_INIT = 16'h9696;
    SB_CARRY add_626_3 (.CI(n27522), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n27523));
    SB_LUT4 i5_4_lut_adj_1035 (.I0(n33886), .I1(n34009), .I2(\data_in_frame[16] [7]), 
            .I3(\data_in_frame[14] [5]), .O(n12_adj_3700));
    defparam i5_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_CARRY add_44_9 (.CI(n27497), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27498));
    SB_LUT4 i6_4_lut_adj_1036 (.I0(\data_in_frame[17] [2]), .I1(n12_adj_3700), 
            .I2(n34212), .I3(\data_in_frame[15] [1]), .O(n29870));
    defparam i6_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1037 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10] [5]), 
            .I2(\data_in_frame[13] [0]), .I3(GND_net), .O(n34275));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1037.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1038 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n33974));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1038.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1039 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [1]), 
            .I2(n17145), .I3(GND_net), .O(n34293));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1039.LUT_INIT = 16'h9696;
    SB_LUT4 add_626_2_lut (.I0(GND_net), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3190), .I3(GND_net), .O(n2236[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_626_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_44_8_lut (.I0(n6), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27496), .O(n33242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1040 (.I0(n16668), .I1(n17256), .I2(\data_out_frame[17] [5]), 
            .I3(n33932), .O(n34257));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_CARRY add_626_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), .I1(tx_transmit_N_3190), 
            .CO(n27522));
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18346));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1041 (.I0(n16668), .I1(n17256), .I2(n17425), 
            .I3(\data_out_frame[20] [0]), .O(n34073));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_33_lut (.I0(n6), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27521), .O(n2_adj_3663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_8 (.CI(n27496), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27497));
    SB_LUT4 i1_2_lut_4_lut_adj_1042 (.I0(n35783), .I1(\data_out_frame[20] [3]), 
            .I2(n35798), .I3(n33932), .O(n34046));
    defparam i1_2_lut_4_lut_adj_1042.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18345));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18344));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1043 (.I0(n16715), .I1(n33940), .I2(GND_net), 
            .I3(GND_net), .O(n16815));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18342));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18341));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1044 (.I0(n35783), .I1(\data_out_frame[20] [3]), 
            .I2(n35798), .I3(\data_out_frame[20] [2]), .O(n33911));
    defparam i1_2_lut_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1045 (.I0(\data_in_frame[6] [0]), .I1(n33974), 
            .I2(n16624), .I3(n17145), .O(n10_adj_3701));   // verilog/coms.v(70[16:41])
    defparam i4_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1046 (.I0(n16715), .I1(n10_adj_3701), .I2(n7), 
            .I3(GND_net), .O(n16876));   // verilog/coms.v(70[16:41])
    defparam i5_3_lut_adj_1046.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34133));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18340));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1048 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[8] [4]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n33859));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1049 (.I0(n16876), .I1(\data_in_frame[12] [6]), 
            .I2(n16815), .I3(GND_net), .O(n34159));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1049.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1050 (.I0(n16748), .I1(n16624), .I2(n33859), 
            .I3(n16789), .O(n10_adj_3702));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1051 (.I0(\data_in_frame[6] [3]), .I1(n10_adj_3702), 
            .I2(n34159), .I3(GND_net), .O(n17354));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_1051.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1052 (.I0(n34133), .I1(n34159), .I2(\data_in_frame[10] [7]), 
            .I3(n33817), .O(n12_adj_3703));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(n93[1]), .I1(n63), .I2(n19), .I3(n33787), 
            .O(n33126));   // verilog/coms.v(143[4] 146[7])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hb0bb;
    SB_LUT4 add_44_32_lut (.I0(n6), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27520), .O(n2_adj_3661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1053 (.I0(\data_in_frame[11] [0]), .I1(n12_adj_3703), 
            .I2(n34275), .I3(n17338), .O(n17357));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [20]), 
            .I3(n9_adj_3705), .O(n33170));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1054 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [21]), 
            .I3(n9_adj_3705), .O(n33168));
    defparam i1_2_lut_3_lut_4_lut_adj_1054.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1055 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [10]), 
            .I3(n9_adj_3705), .O(n33182));
    defparam i1_2_lut_3_lut_4_lut_adj_1055.LUT_INIT = 16'hf020;
    SB_LUT4 i1_3_lut_4_lut_adj_1056 (.I0(n11748), .I1(n33787), .I2(n224_c), 
            .I3(\FRAME_MATCHER.state [3]), .O(n33140));
    defparam i1_3_lut_4_lut_adj_1056.LUT_INIT = 16'hf200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1057 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [11]), 
            .I3(n9_adj_3705), .O(n33180));
    defparam i1_2_lut_3_lut_4_lut_adj_1057.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\data_in_frame[16] [1]), .I1(n30677), 
            .I2(GND_net), .I3(GND_net), .O(n34076));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16631));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1060 (.I0(\data_in_frame[7] [1]), .I1(n17114), 
            .I2(Kp_23__N_871), .I3(n17338), .O(n34156));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1061 (.I0(n33856), .I1(n34156), .I2(\data_in_frame[11] [3]), 
            .I3(\data_in_frame[4] [7]), .O(n12_adj_3706));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1062 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [26]), 
            .I3(n9_adj_3705), .O(n33162));
    defparam i1_2_lut_3_lut_4_lut_adj_1062.LUT_INIT = 16'hf020;
    SB_LUT4 i6_4_lut_adj_1063 (.I0(\data_in_frame[6] [5]), .I1(n12_adj_3706), 
            .I2(n34272), .I3(\data_in_frame[9] [2]), .O(n30393));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1064 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [9]), 
            .I3(n9_adj_3705), .O(n33184));
    defparam i1_2_lut_3_lut_4_lut_adj_1064.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1065 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [28]), 
            .I3(n9_adj_3705), .O(n33228));
    defparam i1_2_lut_3_lut_4_lut_adj_1065.LUT_INIT = 16'hf020;
    SB_LUT4 i4_4_lut_adj_1066 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[6] [6]), 
            .I2(n33817), .I3(n6_adj_3707), .O(n16824));   // verilog/coms.v(76[16:50])
    defparam i4_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1067 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [16]), 
            .I3(n9_adj_3705), .O(n33174));
    defparam i1_2_lut_3_lut_4_lut_adj_1067.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34209));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1069 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [24]), 
            .I3(n9_adj_3705), .O(n33200));
    defparam i1_2_lut_3_lut_4_lut_adj_1069.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1070 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [7]), 
            .I3(n9_adj_3705), .O(n33198));
    defparam i1_2_lut_3_lut_4_lut_adj_1070.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1071 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [29]), 
            .I3(n9_adj_3705), .O(n33160));
    defparam i1_2_lut_3_lut_4_lut_adj_1071.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n34147));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1073 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [12]), 
            .I3(n9_adj_3705), .O(n33218));
    defparam i1_2_lut_3_lut_4_lut_adj_1073.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n33836));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1075 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [25]), 
            .I3(n9_adj_3705), .O(n33164));
    defparam i1_2_lut_3_lut_4_lut_adj_1075.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(n16741), .I1(n9), .I2(GND_net), .I3(GND_net), 
            .O(n17362));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1077 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [8]), 
            .I3(n9_adj_3705), .O(n33186));
    defparam i1_2_lut_3_lut_4_lut_adj_1077.LUT_INIT = 16'hf020;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(\data_in_frame[8] [0]), .I1(n16741), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[10] [3]), .O(n10_adj_3708));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1079 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [30]), 
            .I3(n9_adj_3705), .O(n33158));
    defparam i1_2_lut_3_lut_4_lut_adj_1079.LUT_INIT = 16'hf020;
    SB_LUT4 i5_3_lut_adj_1080 (.I0(\data_in_frame[6] [0]), .I1(n10_adj_3708), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n33917));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_in_frame[12] [3]), .I1(n16093), 
            .I2(GND_net), .I3(GND_net), .O(n34009));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1082 (.I0(n17141), .I1(Kp_23__N_1058), .I2(n33917), 
            .I3(n6_adj_3709), .O(n16748));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1083 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [19]), 
            .I3(n9_adj_3705), .O(n33172));
    defparam i1_2_lut_3_lut_4_lut_adj_1083.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1084 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [22]), 
            .I3(n9_adj_3705), .O(n33166));
    defparam i1_2_lut_3_lut_4_lut_adj_1084.LUT_INIT = 16'hf020;
    SB_LUT4 i5_4_lut_3_lut_4_lut (.I0(n35783), .I1(n33923), .I2(n16668), 
            .I3(\data_out_frame[17] [4]), .O(n12_adj_3710));
    defparam i5_4_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3692));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1085 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [6]), 
            .I3(n9_adj_3705), .O(n33188));
    defparam i1_2_lut_3_lut_4_lut_adj_1085.LUT_INIT = 16'hf020;
    SB_LUT4 i33060_2_lut (.I0(\data_out_frame[5] [4]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n39058));
    defparam i33060_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n41872));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(n35995), .I1(n34018), .I2(GND_net), 
            .I3(GND_net), .O(n30720));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1087 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [5]), 
            .I3(n9_adj_3705), .O(n33190));
    defparam i1_2_lut_3_lut_4_lut_adj_1087.LUT_INIT = 16'hf020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1088 (.I0(n11748), .I1(n33787), .I2(\FRAME_MATCHER.state [4]), 
            .I3(n9_adj_3705), .O(n33142));
    defparam i1_2_lut_3_lut_4_lut_adj_1088.LUT_INIT = 16'hf020;
    SB_LUT4 i2_3_lut_adj_1089 (.I0(n30692), .I1(n4_c), .I2(\data_in_frame[6] [7]), 
            .I3(GND_net), .O(n34272));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1089.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1090 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [7]), 
            .I2(n30201), .I3(GND_net), .O(n30655));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_1090.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3711));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1092 (.I0(n34272), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[7] [2]), .I3(n6_adj_3711), .O(n34254));
    defparam i4_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1093 (.I0(\data_in_frame[0] [7]), .I1(n34123), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n17141));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1093.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(\data_in_frame[12] [0]), .I1(n29915), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n34186));
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(\data_in_frame[13] [7]), .I1(n33895), 
            .I2(n34227), .I3(n6_adj_3712), .O(n35254));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(n29838), .I1(n16952), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3713));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1097 (.I0(n33968), .I1(n34209), .I2(\data_in_frame[14] [2]), 
            .I3(n6_adj_3713), .O(n34018));
    defparam i4_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1098 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n33767), .O(n33775));
    defparam i1_2_lut_3_lut_4_lut_adj_1098.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_4_lut_adj_1099 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[14] [4]), 
            .I2(n34060), .I3(\data_out_frame[16] [5]), .O(n17259));
    defparam i1_2_lut_4_lut_adj_1099.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1100 (.I0(\data_in_frame[14] [1]), .I1(n34018), 
            .I2(n35254), .I3(GND_net), .O(n30661));
    defparam i2_3_lut_adj_1100.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1101 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n33758), .O(n33766));
    defparam i1_2_lut_3_lut_4_lut_adj_1101.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_1102 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[14] [0]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[16] [2]), 
            .O(n16989));
    defparam i2_3_lut_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1103 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [1]), .O(n34177));
    defparam i2_3_lut_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 equal_119_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_3689));   // verilog/coms.v(154[7:23])
    defparam equal_119_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1104 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(n34180), .O(n34));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1105 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n33908));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1106 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n33948));
    defparam i1_2_lut_3_lut_adj_1106.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1107 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n34278));
    defparam i1_2_lut_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1108 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n33880));
    defparam i1_2_lut_3_lut_adj_1108.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1109 (.I0(n29836), .I1(\data_out_frame[18] [3]), 
            .I2(\data_out_frame[18] [4]), .I3(GND_net), .O(n15_adj_3714));
    defparam i2_2_lut_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1110 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [31]), .O(n7_adj_3675));
    defparam i1_2_lut_4_lut_adj_1110.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1111 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [30]), .O(n33274));
    defparam i1_2_lut_4_lut_adj_1111.LUT_INIT = 16'hdc00;
    SB_LUT4 i2_2_lut_4_lut_adj_1112 (.I0(n33961), .I1(\data_out_frame[12] [3]), 
            .I2(n17128), .I3(\data_out_frame[13] [0]), .O(n10_adj_3715));
    defparam i2_2_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i21044_2_lut_3_lut_4_lut (.I0(n16280), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n34510), .O(n2540));   // verilog/coms.v(148[5:9])
    defparam i21044_2_lut_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_3_lut_4_lut_adj_1113 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[6] [1]), .I3(\data_out_frame[6] [6]), .O(n33945));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1114 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [29]), .O(n33262));
    defparam i1_2_lut_4_lut_adj_1114.LUT_INIT = 16'hdc00;
    SB_LUT4 i2_3_lut_4_lut_adj_1115 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[9] [0]), .I3(\data_out_frame[11] [1]), .O(n34266));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1116 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[8] [0]), .O(n33993));
    defparam i2_3_lut_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i9_3_lut_4_lut (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [1]), .I3(n34057), .O(n26_adj_3716));
    defparam i9_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1117 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [28]), .O(n33258));
    defparam i1_2_lut_4_lut_adj_1117.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1118 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [27]), .O(n7_adj_3673));
    defparam i1_2_lut_4_lut_adj_1118.LUT_INIT = 16'hdc00;
    SB_LUT4 i2_3_lut_4_lut_adj_1119 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[17] [3]), .I3(\data_out_frame[17] [7]), 
            .O(n33923));
    defparam i2_3_lut_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1120 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [6]), .I3(\data_out_frame[7] [7]), .O(n6_adj_3717));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1121 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n17307));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1122 (.I0(\data_out_frame[13] [5]), .I1(n1515), 
            .I2(n16066), .I3(\data_out_frame[13] [6]), .O(n29832));
    defparam i2_3_lut_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1123 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [26]), .O(n33348));
    defparam i1_2_lut_4_lut_adj_1123.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(n16906), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n34215));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1125 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(n17040), .I3(\data_out_frame[15] [3]), .O(n16668));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1126 (.I0(\data_out_frame[13] [0]), .I1(n16929), 
            .I2(\data_out_frame[12] [5]), .I3(n16923), .O(n6_adj_3718));
    defparam i2_2_lut_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(n30663), .I1(\data_out_frame[16] [6]), 
            .I2(n29810), .I3(GND_net), .O(n33795));
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1128 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [25]), .O(n33344));
    defparam i1_2_lut_4_lut_adj_1128.LUT_INIT = 16'hdc00;
    SB_LUT4 i2_3_lut_4_lut_adj_1129 (.I0(n34320), .I1(n34326), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[14] [1]), .O(n34003));
    defparam i2_3_lut_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1130 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [24]), .O(n33288));
    defparam i1_2_lut_4_lut_adj_1130.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(\data_out_frame[17] [0]), .I1(n16585), 
            .I2(\data_out_frame[17] [1]), .I3(GND_net), .O(n34120));
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1132 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[6] [4]), .O(n14_adj_3719));   // verilog/coms.v(71[16:34])
    defparam i5_3_lut_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n16_adj_3720));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1133 (.I0(\data_out_frame[20] [1]), .I1(n16668), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n34242));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1133.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(n16066), .I1(\data_out_frame[12] [0]), 
            .I2(n34003), .I3(GND_net), .O(n34006));
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1135 (.I0(n30663), .I1(n34111), .I2(n34245), 
            .I3(n29836), .O(n30686));
    defparam i2_3_lut_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1136 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [23]), .O(n7_adj_3671));
    defparam i1_2_lut_4_lut_adj_1136.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1137 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [22]), .O(n33340));
    defparam i1_2_lut_4_lut_adj_1137.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1138 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [21]), .O(n33336));
    defparam i1_2_lut_4_lut_adj_1138.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1139 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [20]), .O(n33332));
    defparam i1_2_lut_4_lut_adj_1139.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1140 (.I0(tx_active), .I1(\r_SM_Main_2__N_3298[0] ), 
            .I2(n25598), .I3(n11748), .O(n14163));
    defparam i1_2_lut_4_lut_adj_1140.LUT_INIT = 16'hef00;
    SB_LUT4 i1_2_lut_4_lut_adj_1141 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [19]), .O(n33328));
    defparam i1_2_lut_4_lut_adj_1141.LUT_INIT = 16'hdc00;
    SB_LUT4 i33421_2_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n39105));
    defparam i33421_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1142 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(n16741), .I3(n9), .O(n6_adj_3709));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1143 (.I0(\data_in_frame[14] [5]), .I1(n29571), 
            .I2(n29826), .I3(\data_in_frame[16] [6]), .O(n33971));
    defparam i1_2_lut_3_lut_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 mux_664_i1_3_lut_4_lut (.I0(n31_adj_3618), .I1(n24558), .I2(tx_transmit_N_3190), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n25608));   // verilog/coms.v(147[4] 288[11])
    defparam mux_664_i1_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 i1_2_lut_4_lut_adj_1144 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [18]), .O(n7_adj_3669));
    defparam i1_2_lut_4_lut_adj_1144.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1145 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [17]), .O(n7_adj_3667));
    defparam i1_2_lut_4_lut_adj_1145.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1146 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [16]), .O(n33324));
    defparam i1_2_lut_4_lut_adj_1146.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1147 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [15]), .O(n7_adj_3665));
    defparam i1_2_lut_4_lut_adj_1147.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_3_lut_adj_1148 (.I0(n16748), .I1(\data_in_frame[12] [3]), 
            .I2(n16093), .I3(GND_net), .O(n29571));
    defparam i1_2_lut_3_lut_adj_1148.LUT_INIT = 16'h9696;
    SB_LUT4 i20089_2_lut_4_lut (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [14]), .O(n24574));
    defparam i20089_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1149 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [13]), .O(n64));
    defparam i1_2_lut_4_lut_adj_1149.LUT_INIT = 16'hdc00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21]_c [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3721));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33091_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n39413));   // verilog/coms.v(104[34:55])
    defparam i33091_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3722));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1150 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [12]), .O(n33284));
    defparam i1_2_lut_4_lut_adj_1150.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1151 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [11]), .O(n33320));
    defparam i1_2_lut_4_lut_adj_1151.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_3_lut_adj_1152 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[4] [6]), 
            .I2(n34129), .I3(GND_net), .O(n6_adj_3707));   // verilog/coms.v(76[16:50])
    defparam i1_2_lut_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i31014_4_lut (.I0(n19_adj_3721), .I1(\data_out_frame[22]_c [7]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37334));
    defparam i31014_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1153 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [10]), .O(n33316));
    defparam i1_2_lut_4_lut_adj_1153.LUT_INIT = 16'hdc00;
    SB_LUT4 i31015_3_lut (.I0(n41821), .I1(n37334), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37335));
    defparam i31015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30983_4_lut (.I0(n5_adj_3722), .I1(n39413), .I2(n38883), 
            .I3(\byte_transmit_counter[0] ), .O(n37303));
    defparam i30983_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i30985_4_lut (.I0(n37303), .I1(n37335), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37305));
    defparam i30985_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30984_3_lut (.I0(n41839), .I1(n41833), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37304));
    defparam i30984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1154 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(n16789), .I3(\data_in_frame[8] [6]), .O(n33817));   // verilog/coms.v(76[16:50])
    defparam i2_3_lut_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1155 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [9]), .O(n33312));
    defparam i1_2_lut_4_lut_adj_1155.LUT_INIT = 16'hdc00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21]_c [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3723));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1156 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [8]), .O(n33308));
    defparam i1_2_lut_4_lut_adj_1156.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1157 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [7]), .O(n33292));
    defparam i1_2_lut_4_lut_adj_1157.LUT_INIT = 16'hdc00;
    SB_LUT4 i33084_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n39406));   // verilog/coms.v(104[34:55])
    defparam i33084_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3724));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31011_4_lut (.I0(n19_adj_3723), .I1(\data_out_frame[22]_c [6]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37331));
    defparam i31011_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1158 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [6]), .O(n33304));
    defparam i1_2_lut_4_lut_adj_1158.LUT_INIT = 16'hdc00;
    SB_LUT4 i31012_3_lut (.I0(n41815), .I1(n37331), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37332));
    defparam i31012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30980_4_lut (.I0(n5_adj_3724), .I1(n39406), .I2(n38883), 
            .I3(\byte_transmit_counter[0] ), .O(n37300));
    defparam i30980_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i30982_4_lut (.I0(n37300), .I1(n37332), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37302));
    defparam i30982_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30981_3_lut (.I0(n41851), .I1(n41845), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37301));
    defparam i30981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1159 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [5]), .O(n33300));
    defparam i1_2_lut_4_lut_adj_1159.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1160 (.I0(n16417), .I1(n224_c), .I2(n14163), 
            .I3(\FRAME_MATCHER.state [4]), .O(n33296));
    defparam i1_2_lut_4_lut_adj_1160.LUT_INIT = 16'hdc00;
    SB_LUT4 mux_1027_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n4423));
    defparam mux_1027_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21]_c [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3725));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n41872_bdd_4_lut (.I0(n41872), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n41875));
    defparam n41872_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13842_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n18349));
    defparam i13842_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13843_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n18350));
    defparam i13843_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13844_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n18351));
    defparam i13844_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(\byte_transmit_counter[1] ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n39401));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 mux_1027_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14] [7]), .O(n4446));
    defparam mux_1027_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3727));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1161 (.I0(n17357), .I1(\data_in_frame[6] [3]), 
            .I2(n10_adj_3702), .I3(n34159), .O(n34218));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i13845_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n18352));
    defparam i13845_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31008_4_lut (.I0(n19_adj_3725), .I1(\data_out_frame[22]_c [5]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37328));
    defparam i31008_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13846_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n18353));
    defparam i13846_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31009_3_lut (.I0(n41809), .I1(n37328), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37329));
    defparam i31009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13847_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n18354));
    defparam i13847_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30977_4_lut (.I0(n5_adj_3727), .I1(\byte_transmit_counter[0] ), 
            .I2(n38883), .I3(n39401), .O(n37297));
    defparam i30977_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35527 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n41866));
    defparam byte_transmit_counter_0__bdd_4_lut_35527.LUT_INIT = 16'he4aa;
    SB_LUT4 i30979_4_lut (.I0(n37297), .I1(n37329), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37299));
    defparam i30979_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n41866_bdd_4_lut (.I0(n41866), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n41869));
    defparam n41866_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13848_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n18355));
    defparam i13848_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35522 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n41860));
    defparam byte_transmit_counter_0__bdd_4_lut_35522.LUT_INIT = 16'he4aa;
    SB_LUT4 n41860_bdd_4_lut (.I0(n41860), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n41863));
    defparam n41860_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13849_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n18356));
    defparam i13849_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35517 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n41854));
    defparam byte_transmit_counter_0__bdd_4_lut_35517.LUT_INIT = 16'he4aa;
    SB_LUT4 i13786_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n18293));
    defparam i13786_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41854_bdd_4_lut (.I0(n41854), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n41857));
    defparam n41854_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35512 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n41848));
    defparam byte_transmit_counter_0__bdd_4_lut_35512.LUT_INIT = 16'he4aa;
    SB_LUT4 n41848_bdd_4_lut (.I0(n41848), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n41851));
    defparam n41848_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35507 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n41842));
    defparam byte_transmit_counter_0__bdd_4_lut_35507.LUT_INIT = 16'he4aa;
    SB_LUT4 i30978_3_lut (.I0(n41863), .I1(n41857), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37298));
    defparam i30978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1162 (.I0(n4025), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2467 [3]), 
            .O(n13950));
    defparam i1_2_lut_3_lut_4_lut_adj_1162.LUT_INIT = 16'h2000;
    SB_LUT4 i13787_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n18294));
    defparam i13787_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13788_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n18295));
    defparam i13788_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41842_bdd_4_lut (.I0(n41842), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n41845));
    defparam n41842_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35502 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n41836));
    defparam byte_transmit_counter_0__bdd_4_lut_35502.LUT_INIT = 16'he4aa;
    SB_LUT4 n41836_bdd_4_lut (.I0(n41836), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n41839));
    defparam n41836_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35497 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n41830));
    defparam byte_transmit_counter_0__bdd_4_lut_35497.LUT_INIT = 16'he4aa;
    SB_LUT4 i13789_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n18296));
    defparam i13789_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41830_bdd_4_lut (.I0(n41830), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n41833));
    defparam n41830_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13790_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n18297));
    defparam i13790_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35492 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n41824));
    defparam byte_transmit_counter_0__bdd_4_lut_35492.LUT_INIT = 16'he4aa;
    SB_LUT4 i13791_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n18298));
    defparam i13791_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41824_bdd_4_lut (.I0(n41824), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n41827));
    defparam n41824_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35487 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n41818));
    defparam byte_transmit_counter_0__bdd_4_lut_35487.LUT_INIT = 16'he4aa;
    SB_LUT4 i13792_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n18299));
    defparam i13792_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41818_bdd_4_lut (.I0(n41818), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n41821));
    defparam n41818_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35482 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n41812));
    defparam byte_transmit_counter_0__bdd_4_lut_35482.LUT_INIT = 16'he4aa;
    SB_LUT4 n41812_bdd_4_lut (.I0(n41812), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n41815));
    defparam n41812_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21]_c [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3728));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31005_4_lut (.I0(n19_adj_3728), .I1(\data_out_frame[22]_c [4]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37325));
    defparam i31005_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i34290_3_lut (.I0(n41827), .I1(n41743), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40612));
    defparam i34290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31006_3_lut (.I0(n41803), .I1(n37325), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37326));
    defparam i31006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34294_3_lut (.I0(n41881), .I1(n40612), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n40616));   // verilog/coms.v(104[34:55])
    defparam i34294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13793_3_lut_4_lut (.I0(n8_adj_3689), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n18300));
    defparam i13793_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35477 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n41806));
    defparam byte_transmit_counter_0__bdd_4_lut_35477.LUT_INIT = 16'he4aa;
    SB_LUT4 i34295_4_lut (.I0(n40616), .I1(n37326), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i34295_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33020_2_lut (.I0(\data_out_frame[0] [3]), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n39029));   // verilog/coms.v(104[34:55])
    defparam i33020_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21]_c [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3729));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1027_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14] [6]), .O(n4445));
    defparam mux_1027_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n39029), .I2(byte_transmit_counter[2]), .I3(\byte_transmit_counter[0] ), 
            .O(n6_adj_3730));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3731));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31002_4_lut (.I0(n19_adj_3729), .I1(\data_out_frame[22]_c [3]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37322));
    defparam i31002_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31003_3_lut (.I0(n41797), .I1(n37322), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37323));
    defparam i31003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30974_3_lut (.I0(n5_adj_3731), .I1(n6_adj_3730), .I2(n38883), 
            .I3(GND_net), .O(n37294));
    defparam i30974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30976_4_lut (.I0(n37294), .I1(n37323), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37296));
    defparam i30976_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30975_3_lut (.I0(n41875), .I1(n41869), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37295));
    defparam i30975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34666_2_lut_3_lut_3_lut_3_lut (.I0(n4025), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n17572));
    defparam i34666_2_lut_3_lut_3_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1163 (.I0(n35783), .I1(\data_out_frame[18] [0]), 
            .I2(n16102), .I3(n33911), .O(n33912));
    defparam i1_2_lut_3_lut_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1027_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14] [5]), .O(n4444));
    defparam mux_1027_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i33126_2_lut (.I0(\data_out_frame[0] [2]), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n39026));   // verilog/coms.v(104[34:55])
    defparam i33126_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21]_c [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3732));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1027_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[14] [4]), .O(n4443));
    defparam mux_1027_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(n39026), .I2(byte_transmit_counter[2]), .I3(\byte_transmit_counter[0] ), 
            .O(n6_adj_3733));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3734));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30999_4_lut (.I0(n19_adj_3732), .I1(\data_out_frame[22]_c [2]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37319));
    defparam i30999_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31000_3_lut (.I0(n41791), .I1(n37319), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37320));
    defparam i31000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30971_3_lut (.I0(n5_adj_3734), .I1(n6_adj_3733), .I2(n38883), 
            .I3(GND_net), .O(n37291));
    defparam i30971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30973_4_lut (.I0(n37291), .I1(n37320), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37293));
    defparam i30973_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30972_3_lut (.I0(n41749), .I1(n41737), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37292));
    defparam i30972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1164 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [1]), .I3(n17145), .O(n33940));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21]_c [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_3735));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1165 (.I0(\data_out_frame[15] [7]), .I1(n29832), 
            .I2(n16086), .I3(\data_out_frame[14] [0]), .O(n34043));
    defparam i1_2_lut_3_lut_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i33061_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n39382));   // verilog/coms.v(104[34:55])
    defparam i33061_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1166 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(\data_out_frame[20] [1]), .I3(n17279), .O(n6_adj_3736));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1167 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[13] [0]), .O(n6_adj_3697));
    defparam i1_2_lut_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_3737));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30996_4_lut (.I0(n19_adj_3735), .I1(\data_out_frame[22]_c [1]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n37316));
    defparam i30996_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30997_3_lut (.I0(n41785), .I1(n37316), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37317));
    defparam i30997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30968_4_lut (.I0(n5_adj_3737), .I1(n39382), .I2(n38883), 
            .I3(\byte_transmit_counter[0] ), .O(n37288));
    defparam i30968_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i30970_4_lut (.I0(n37288), .I1(n37317), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n37290));
    defparam i30970_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30969_3_lut (.I0(n41761), .I1(n41755), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n37289));
    defparam i30969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1168 (.I0(n17141), .I1(n29784), .I2(\data_in_frame[12] [0]), 
            .I3(n34153), .O(n29838));
    defparam i2_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(n17141), .I1(n29784), .I2(n34186), 
            .I3(GND_net), .O(n6_adj_3712));
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1170 (.I0(n33943), .I1(\data_in_frame[11] [4]), 
            .I2(n30393), .I3(n34254), .O(n30610));
    defparam i2_3_lut_4_lut_adj_1170.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1171 (.I0(n33943), .I1(\data_in_frame[11] [4]), 
            .I2(n35254), .I3(GND_net), .O(n34108));
    defparam i1_2_lut_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1172 (.I0(Kp_23__N_1537), .I1(n34140), .I2(n30710), 
            .I3(\data_in_frame[15] [5]), .O(n34906));
    defparam i2_3_lut_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1027_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14] [3]), .O(n4442));
    defparam mux_1027_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1173 (.I0(n17265), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(n34199), .O(n16066));
    defparam i1_2_lut_3_lut_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n13914));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'heeee;
    SB_LUT4 i28299_4_lut (.I0(n25604), .I1(\FRAME_MATCHER.state [3]), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n13914), .O(n34543));
    defparam i28299_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_1175 (.I0(\FRAME_MATCHER.state [1]), .I1(n25604), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n4_adj_3738));
    defparam i1_3_lut_adj_1175.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_713_i1_4_lut (.I0(n24585), .I1(n25608), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n25610));   // verilog/coms.v(147[4] 288[11])
    defparam mux_713_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i32854_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n25610), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n4_adj_3738), .O(n39174));   // verilog/coms.v(147[4] 288[11])
    defparam i32854_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 mux_1027_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14] [2]), .O(n4441));
    defparam mux_1027_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n17265), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[13] [6]), .I3(n34236), .O(n7_adj_3739));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1176 (.I0(Kp_23__N_1537), .I1(n34140), .I2(n34206), 
            .I3(n10_adj_3590), .O(n36064));
    defparam i5_3_lut_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 n41806_bdd_4_lut (.I0(n41806), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n41809));
    defparam n41806_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1027_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14] [1]), .O(n4440));
    defparam mux_1027_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35472 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n41800));
    defparam byte_transmit_counter_0__bdd_4_lut_35472.LUT_INIT = 16'he4aa;
    SB_LUT4 n41800_bdd_4_lut (.I0(n41800), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n41803));
    defparam n41800_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30939_4_lut (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[1] [1]), .O(n37194));
    defparam i30939_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1177 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(n17145), .I3(GND_net), .O(n6_adj_3693));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i13834_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n18341));
    defparam i13834_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13835_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n18342));
    defparam i13835_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35467 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n41794));
    defparam byte_transmit_counter_0__bdd_4_lut_35467.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1027_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14] [0]), .O(n4439));
    defparam mux_1027_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13836_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n18343));
    defparam i13836_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13837_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n18344));
    defparam i13837_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1178 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [4]), .O(n38_adj_3741));
    defparam i14_4_lut_adj_1178.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut_adj_1179 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [4]), .O(n39_adj_3742));
    defparam i15_4_lut_adj_1179.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\FRAME_MATCHER.state [31]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3676));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h8888;
    SB_LUT4 n41794_bdd_4_lut (.I0(n41794), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n41797));
    defparam n41794_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1181 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[16] [5]), 
            .I2(n35995), .I3(n29826), .O(n34093));
    defparam i2_3_lut_4_lut_adj_1181.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1182 (.I0(\data_in_frame[14] [5]), .I1(n29571), 
            .I2(\data_in_frame[17] [0]), .I3(GND_net), .O(n34251));
    defparam i1_2_lut_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1183 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n29818), .I3(GND_net), .O(n34070));
    defparam i1_2_lut_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\FRAME_MATCHER.state [27]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3674));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1185 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n33792), .O(n18_adj_3609));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1186 (.I0(\data_in_frame[15] [5]), .I1(n16824), 
            .I2(n30393), .I3(\data_in_frame[17] [6]), .O(n34263));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_4_lut_adj_1186.LUT_INIT = 16'h9669;
    SB_LUT4 i20419_2_lut_3_lut (.I0(n34510), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n24905));
    defparam i20419_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\FRAME_MATCHER.state [23]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3672));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h8888;
    SB_LUT4 i13838_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n18345));
    defparam i13838_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13839_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n18346));
    defparam i13839_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1188 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [3]), .O(n37_adj_3743));
    defparam i13_4_lut_adj_1188.LUT_INIT = 16'h2000;
    SB_LUT4 i30935_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [1]), .I3(\data_in_frame[0] [6]), .O(n37190));
    defparam i30935_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\FRAME_MATCHER.state [18]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3670));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h8888;
    SB_LUT4 i22_4_lut (.I0(n37_adj_3743), .I1(n39_adj_3742), .I2(n38_adj_3741), 
            .I3(n37194), .O(n46));
    defparam i22_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\FRAME_MATCHER.state [17]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3668));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(\FRAME_MATCHER.state [15]), .I1(n220_c), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3666));
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h8888;
    SB_LUT4 i30937_4_lut (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[2] [2]), .O(n37192));
    defparam i30937_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30926_4_lut (.I0(n11748), .I1(n37137), .I2(n37135), .I3(n33787), 
            .O(n220_c));
    defparam i30926_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 i23_3_lut (.I0(n37192), .I1(n46), .I2(n37190), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2467 [3]));
    defparam i23_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i20814_2_lut (.I0(\FRAME_MATCHER.state [14]), .I1(n220_c), .I2(GND_net), 
            .I3(GND_net), .O(n25301));
    defparam i20814_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30885_2_lut (.I0(n16404), .I1(n2857), .I2(GND_net), .I3(GND_net), 
            .O(n37135));
    defparam i30885_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1192 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n35805));
    defparam i2_3_lut_adj_1192.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1193 (.I0(\FRAME_MATCHER.state [13]), .I1(n11748), 
            .I2(n37188), .I3(GND_net), .O(n33134));
    defparam i1_3_lut_adj_1193.LUT_INIT = 16'h0808;
    SB_LUT4 i1_4_lut_adj_1194 (.I0(n25604), .I1(n39105), .I2(n35805), 
            .I3(\FRAME_MATCHER.state [3]), .O(n4025));
    defparam i1_4_lut_adj_1194.LUT_INIT = 16'h0544;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35462 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n41788));
    defparam byte_transmit_counter_0__bdd_4_lut_35462.LUT_INIT = 16'he4aa;
    SB_LUT4 i13840_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n18347));
    defparam i13840_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13841_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n18348));
    defparam i13841_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state_31__N_2467 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33747));
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h4444;
    SB_LUT4 i216_3_lut (.I0(n16420), .I1(n3761), .I2(n11748), .I3(GND_net), 
            .O(n224_c));   // verilog/coms.v(113[11:12])
    defparam i216_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1196 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(n34147), .I3(n33836), .O(Kp_23__N_1537));
    defparam i2_3_lut_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i28324_4_lut (.I0(n16256), .I1(n4_adj_3610), .I2(n6_adj_3631), 
            .I3(\FRAME_MATCHER.state [2]), .O(n34572));
    defparam i28324_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i2_3_lut_4_lut_adj_1197 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[18] [5]), .I3(\data_in_frame[18] [4]), .O(n33801));
    defparam i2_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1198 (.I0(\FRAME_MATCHER.i [31]), .I1(n16403), 
            .I2(n34572), .I3(n11748), .O(n9_adj_3705));
    defparam i2_4_lut_adj_1198.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1199 (.I0(\FRAME_MATCHER.state [3]), .I1(n14163), 
            .I2(n9_adj_3705), .I3(n4_adj_3744), .O(n14_adj_3745));
    defparam i1_4_lut_adj_1199.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_4_lut_adj_1200 (.I0(\FRAME_MATCHER.state [1]), .I1(n14_adj_3745), 
            .I2(n33747), .I3(n16280), .O(n33382));
    defparam i1_4_lut_adj_1200.LUT_INIT = 16'hccec;
    SB_LUT4 n41878_bdd_4_lut_4_lut (.I0(\data_out_frame[0] [4]), .I1(\byte_transmit_counter[0] ), 
            .I2(byte_transmit_counter[2]), .I3(n41878), .O(n41881));
    defparam n41878_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_LUT4 n41788_bdd_4_lut (.I0(n41788), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n41791));
    defparam n41788_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i28215_2_lut (.I0(n16420), .I1(n3761), .I2(GND_net), .I3(GND_net), 
            .O(n34455));
    defparam i28215_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 select_362_Select_1_i5_4_lut (.I0(n63), .I1(n16404), .I2(n2857), 
            .I3(n93[1]), .O(n5_adj_3746));
    defparam select_362_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i20764_2_lut (.I0(n93[1]), .I1(n9783), .I2(GND_net), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2435 [1]));   // verilog/coms.v(157[6] 159[9])
    defparam i20764_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut_adj_1201 (.I0(n93[1]), .I1(n5_adj_3746), .I2(n34455), 
            .I3(n63), .O(n6_adj_3747));
    defparam i2_4_lut_adj_1201.LUT_INIT = 16'hcecf;
    SB_LUT4 i3_4_lut_adj_1202 (.I0(n35990), .I1(n6_adj_3747), .I2(\FRAME_MATCHER.state_31__N_2435 [1]), 
            .I3(n16405), .O(n42066));
    defparam i3_4_lut_adj_1202.LUT_INIT = 16'hddfd;
    SB_LUT4 i13802_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n18309));
    defparam i13802_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13803_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n18310));
    defparam i13803_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1027_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n4438));
    defparam mux_1027_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13804_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18311));
    defparam i13804_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35457 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n41782));
    defparam byte_transmit_counter_0__bdd_4_lut_35457.LUT_INIT = 16'he4aa;
    SB_LUT4 i13805_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18312));
    defparam i13805_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1027_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n4437));
    defparam mux_1027_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13806_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18313));
    defparam i13806_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13807_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18314));
    defparam i13807_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13808_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18315));
    defparam i13808_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[20] [6]), .I1(n34248), 
            .I2(GND_net), .I3(GND_net), .O(n34249));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(n33932), .I1(n34082), .I2(GND_net), 
            .I3(GND_net), .O(n34084));
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 n41782_bdd_4_lut (.I0(n41782), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n41785));
    defparam n41782_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[20] [2]), .I1(n34030), 
            .I2(GND_net), .I3(GND_net), .O(n34031));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i13809_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18316));
    defparam i13809_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1027_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n4436));
    defparam mux_1027_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1206 (.I0(\data_out_frame[19] [6]), .I1(n16102), 
            .I2(n34073), .I3(n6_adj_3736), .O(n35129));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1206.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_out_frame[17] [6]), .I1(n34281), 
            .I2(GND_net), .I3(GND_net), .O(n16102));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i13833_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n18340));
    defparam i13833_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1208 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n6_adj_3630), .I3(n4025), .O(n17568));
    defparam i2_3_lut_4_lut_adj_1208.LUT_INIT = 16'he000;
    SB_LUT4 i6_4_lut_adj_1209 (.I0(n30686), .I1(n12_adj_3710), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[20] [1]), .O(n34030));
    defparam i6_4_lut_adj_1209.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1210 (.I0(n34257), .I1(n34030), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3749));
    defparam i2_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1211 (.I0(n34305), .I1(n34051), .I2(n34114), 
            .I3(n33911), .O(n14_adj_3750));
    defparam i6_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1212 (.I0(n30703), .I1(n14_adj_3750), .I2(n10_adj_3749), 
            .I3(n34082), .O(n34307));
    defparam i7_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1213 (.I0(n34043), .I1(n34284), .I2(\data_out_frame[12] [1]), 
            .I3(n34003), .O(n12_adj_3751));
    defparam i5_4_lut_adj_1213.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1214 (.I0(n16677), .I1(n12_adj_3751), .I2(\data_out_frame[20] [5]), 
            .I3(n34173), .O(n34082));
    defparam i6_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\data_out_frame[18] [5]), .I1(n34082), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3752));
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h6666;
    SB_LUT4 i13826_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n18333));
    defparam i13826_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1216 (.I0(n1716), .I1(n16989), .I2(n34006), .I3(n6_adj_3752), 
            .O(n34248));
    defparam i4_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1217 (.I0(n35798), .I1(n34087), .I2(\data_out_frame[16] [2]), 
            .I3(\data_out_frame[16] [1]), .O(n12_adj_3753));
    defparam i5_4_lut_adj_1217.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1218 (.I0(\data_out_frame[18] [3]), .I1(n12_adj_3753), 
            .I2(\data_out_frame[20] [4]), .I3(n34006), .O(n33932));
    defparam i6_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i13827_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n18334));
    defparam i13827_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1219 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16406), .I3(GND_net), .O(n16404));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_3_lut_adj_1219.LUT_INIT = 16'hfdfd;
    SB_LUT4 i3_4_lut_adj_1220 (.I0(\data_out_frame[18] [2]), .I1(n29879), 
            .I2(n34043), .I3(\data_out_frame[16] [1]), .O(n35798));
    defparam i3_4_lut_adj_1220.LUT_INIT = 16'h9669;
    SB_LUT4 i13828_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n18335));
    defparam i13828_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1221 (.I0(n30316), .I1(n35798), .I2(n34242), 
            .I3(\data_out_frame[17] [3]), .O(n18_adj_3754));
    defparam i7_4_lut_adj_1221.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1222 (.I0(\data_out_frame[19] [5]), .I1(n18_adj_3754), 
            .I2(\data_out_frame[20] [3]), .I3(n34257), .O(n20_adj_3755));
    defparam i9_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i13829_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n18336));
    defparam i13829_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1223 (.I0(n34248), .I1(n20_adj_3755), .I2(n16_adj_3720), 
            .I3(\data_out_frame[20] [2]), .O(n35199));
    defparam i10_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i13830_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n18337));
    defparam i13830_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13831_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n18338));
    defparam i13831_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(n16668), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17279));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i13832_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n18339));
    defparam i13832_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20193_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n16256), .O(n2857));   // verilog/coms.v(221[9:54])
    defparam i20193_3_lut_4_lut.LUT_INIT = 16'h0f08;
    SB_LUT4 i3_4_lut_adj_1225 (.I0(n17279), .I1(n34233), .I2(n34036), 
            .I3(\data_out_frame[19] [5]), .O(n34928));
    defparam i3_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1226 (.I0(n34230), .I1(\data_out_frame[15] [2]), 
            .I2(n16565), .I3(n34024), .O(n15_adj_3756));   // verilog/coms.v(71[16:34])
    defparam i6_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i13772_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n18279));
    defparam i13772_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1227 (.I0(n15_adj_3756), .I1(n33875), .I2(n14_adj_3719), 
            .I3(\data_out_frame[13] [0]), .O(n17425));   // verilog/coms.v(71[16:34])
    defparam i8_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i13773_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n18280));
    defparam i13773_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1228 (.I0(\data_out_frame[19] [4]), .I1(n17425), 
            .I2(n16585), .I3(\data_out_frame[17] [2]), .O(n34036));
    defparam i3_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1229 (.I0(\data_out_frame[17] [3]), .I1(n34036), 
            .I2(n29828), .I3(\data_out_frame[19] [3]), .O(n35096));
    defparam i3_4_lut_adj_1229.LUT_INIT = 16'h9669;
    SB_LUT4 i13774_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n18281));
    defparam i13774_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1027_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n4435));
    defparam mux_1027_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(n29828), .I1(n34120), .I2(n33883), 
            .I3(n30665), .O(n34884));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i13775_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n18282));
    defparam i13775_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1231 (.I0(\data_out_frame[19] [2]), .I1(n34120), 
            .I2(n33795), .I3(\data_out_frame[19] [1]), .O(n34814));
    defparam i3_4_lut_adj_1231.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(n1716), .I1(n34102), .I2(GND_net), 
            .I3(GND_net), .O(n34051));
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1233 (.I0(n30665), .I1(n34051), .I2(\data_out_frame[18] [6]), 
            .I3(\data_out_frame[19] [1]), .O(n35111));
    defparam i3_4_lut_adj_1233.LUT_INIT = 16'h9669;
    SB_LUT4 i13776_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n18283));
    defparam i13776_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1234 (.I0(n33977), .I1(n34215), .I2(n16923), 
            .I3(GND_net), .O(n16585));
    defparam i2_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i13777_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n18284));
    defparam i13777_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\data_out_frame[17] [0]), .I1(n16585), 
            .I2(GND_net), .I3(GND_net), .O(n17051));
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3757));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1237 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(n33833), .I3(n6_adj_3757), .O(n33977));
    defparam i4_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1238 (.I0(n16929), .I1(n33977), .I2(\data_out_frame[12] [5]), 
            .I3(\data_out_frame[14] [7]), .O(n12_adj_3758));
    defparam i5_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1239 (.I0(\data_out_frame[16] [7]), .I1(n12_adj_3758), 
            .I2(n17051), .I3(n29866), .O(n34305));
    defparam i6_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_out_frame[12] [0]), .I1(n34003), 
            .I2(GND_net), .I3(GND_net), .O(n17085));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1027_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n4434));
    defparam mux_1027_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(n30663), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30665));
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16406), .I3(GND_net), .O(n16405));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34024));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(n30663), .I1(n34111), .I2(GND_net), 
            .I3(GND_net), .O(n34079));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1027_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n4433));
    defparam mux_1027_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1245 (.I0(n16906), .I1(\data_out_frame[14] [6]), 
            .I2(\data_out_frame[18] [7]), .I3(n34079), .O(n10_adj_3759));
    defparam i4_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1246 (.I0(n29910), .I1(n10_adj_3759), .I2(\data_out_frame[16] [5]), 
            .I3(GND_net), .O(n29810));
    defparam i5_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1247 (.I0(n16929), .I1(\data_out_frame[12] [5]), 
            .I2(n16923), .I3(GND_net), .O(n29910));
    defparam i2_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i13770_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n18277));
    defparam i13770_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1248 (.I0(\data_out_frame[15] [1]), .I1(n34299), 
            .I2(n6_adj_3718), .I3(\data_out_frame[14] [7]), .O(n34233));
    defparam i1_4_lut_adj_1248.LUT_INIT = 16'h9669;
    SB_LUT4 i13771_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n18278));
    defparam i13771_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1249 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [0]), 
            .I2(n29810), .I3(\data_out_frame[16] [4]), .O(n34102));
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33883));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16809));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1027_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n4432));
    defparam mux_1027_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1252 (.I0(\data_out_frame[11] [5]), .I1(n33880), 
            .I2(n34278), .I3(n33914), .O(n34326));
    defparam i3_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 equal_121_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3740));   // verilog/coms.v(154[7:23])
    defparam equal_121_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_120_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3726));   // verilog/coms.v(154[7:23])
    defparam equal_120_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i4_4_lut_adj_1253 (.I0(n7_adj_3739), .I1(n34054), .I2(n34326), 
            .I3(n29830), .O(n29879));
    defparam i4_4_lut_adj_1253.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_4_lut (.I0(n34510), .I1(n16410), .I2(n4_adj_3621), 
            .I3(n16280), .O(n33787));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'hf5fd;
    SB_LUT4 i4_4_lut_adj_1254 (.I0(\data_out_frame[16] [0]), .I1(n29848), 
            .I2(\data_out_frame[18] [1]), .I3(n34087), .O(n10_adj_3760));
    defparam i4_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1255 (.I0(\data_out_frame[17] [7]), .I1(n10_adj_3760), 
            .I2(n16066), .I3(GND_net), .O(n35783));
    defparam i5_3_lut_adj_1255.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1256 (.I0(\data_out_frame[15] [5]), .I1(n34054), 
            .I2(n1509), .I3(\data_out_frame[13] [3]), .O(n29848));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1257 (.I0(n17392), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n34111));
    defparam i2_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1258 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n34236));
    defparam i2_3_lut_adj_1258.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16677));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1260 (.I0(n33814), .I1(n17002), .I2(\data_out_frame[6] [6]), 
            .I3(n34126), .O(n10_adj_3761));
    defparam i4_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1261 (.I0(\data_out_frame[7] [2]), .I1(n10_adj_3761), 
            .I2(\data_out_frame[11] [5]), .I3(GND_net), .O(n16086));
    defparam i5_3_lut_adj_1261.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1027_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n4431));
    defparam mux_1027_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(n16086), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34042));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1263 (.I0(\data_out_frame[14] [2]), .I1(n17465), 
            .I2(n17265), .I3(GND_net), .O(n34173));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34317));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1265 (.I0(n16066), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n29830));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1266 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[5] [7]), .O(n33833));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1027_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n4430));
    defparam mux_1027_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1267 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[10] [7]), .I3(\data_out_frame[11] [0]), 
            .O(n34230));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1268 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n33814));
    defparam i2_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16594));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33889));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1271 (.I0(n33889), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[10] [3]), .I3(n6_adj_3717), .O(n16929));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(n16929), .I1(n33961), .I2(\data_out_frame[12] [4]), 
            .I3(GND_net), .O(n16906));
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n33820), .I1(\data_out_frame[14] [5]), 
            .I2(n16906), .I3(GND_net), .O(n29866));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35452 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n41764));
    defparam byte_transmit_counter_0__bdd_4_lut_35452.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1027_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n4429));
    defparam mux_1027_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_4_lut_adj_1274 (.I0(\data_out_frame[13] [3]), .I1(n34066), 
            .I2(n1664), .I3(n16594), .O(n12_adj_3762));
    defparam i5_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n33814), .I1(\data_out_frame[5] [0]), .I2(\data_out_frame[10] [3]), 
            .I3(\data_out_frame[11] [7]), .O(n54));   // verilog/coms.v(72[16:27])
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13762_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n18269));
    defparam i13762_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19_4_lut (.I0(n34162), .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[5] [1]), 
            .I3(\data_out_frame[12] [0]), .O(n52));   // verilog/coms.v(72[16:27])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n34311), .I1(n34177), .I2(n34230), .I3(n34060), 
            .O(n53));   // verilog/coms.v(72[16:27])
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13763_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n18270));
    defparam i13763_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13764_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n18271));
    defparam i13764_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1275 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[11] [3]), 
            .I2(n33993), .I3(n34266), .O(n51_adj_3763));   // verilog/coms.v(72[16:27])
    defparam i18_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i13765_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n18272));
    defparam i13765_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i25_4_lut_adj_1276 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[8] [0]), 
            .I2(n17307), .I3(n34), .O(n58));   // verilog/coms.v(72[16:27])
    defparam i25_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1277 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[7] [3]), 
            .I2(n33908), .I3(\data_out_frame[7] [7]), .O(n56));   // verilog/coms.v(72[16:27])
    defparam i23_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1278 (.I0(n33999), .I1(n33889), .I2(n33945), 
            .I3(n33833), .O(n57));   // verilog/coms.v(72[16:27])
    defparam i24_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1279 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[12] [1]), .I3(n33862), .O(n55));   // verilog/coms.v(72[16:27])
    defparam i22_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut_adj_1280 (.I0(n55), .I1(n57), .I2(n56), .I3(n58), 
            .O(n64_adj_3764));   // verilog/coms.v(72[16:27])
    defparam i31_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1281 (.I0(n51_adj_3763), .I1(n53), .I2(n52), 
            .I3(n54), .O(n63_adj_3765));   // verilog/coms.v(72[16:27])
    defparam i30_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i13766_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n18273));
    defparam i13766_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13767_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n18274));
    defparam i13767_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13768_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n18275));
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1282 (.I0(n29832), .I1(n12_adj_3762), .I2(\data_out_frame[13] [0]), 
            .I3(n30663), .O(n35671));
    defparam i6_4_lut_adj_1282.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1283 (.I0(n35671), .I1(n34317), .I2(n34173), 
            .I3(n34215), .O(n12_adj_3766));
    defparam i5_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1284 (.I0(n34042), .I1(n63_adj_3765), .I2(n34302), 
            .I3(n64_adj_3764), .O(n11));
    defparam i4_4_lut_adj_1284.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1285 (.I0(n11), .I1(n26_adj_3716), .I2(\data_out_frame[15] [2]), 
            .I3(n12_adj_3766), .O(n30_adj_3767));
    defparam i13_4_lut_adj_1285.LUT_INIT = 16'h9669;
    SB_LUT4 n41764_bdd_4_lut (.I0(n41764), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n41767));
    defparam n41764_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11_4_lut_adj_1286 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [0]), 
            .I2(n17252), .I3(\data_out_frame[15] [5]), .O(n28_adj_3768));
    defparam i11_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1287 (.I0(n34236), .I1(n29866), .I2(n33935), 
            .I3(\data_out_frame[15] [3]), .O(n29_adj_3769));
    defparam i12_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i13769_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n18276));
    defparam i13769_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13824_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n18331));
    defparam i13824_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1288 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[15] [1]), 
            .I2(n17091), .I3(n17110), .O(n27_adj_3770));
    defparam i10_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i13825_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n18332));
    defparam i13825_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1289 (.I0(n27_adj_3770), .I1(n29_adj_3769), .I2(n28_adj_3768), 
            .I3(n30_adj_3767), .O(n34245));
    defparam i16_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_out_frame[17] [5]), .I1(n33923), 
            .I2(GND_net), .I3(GND_net), .O(n17174));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i13818_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n18325));
    defparam i13818_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34284));
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1292 (.I0(n17174), .I1(n34245), .I2(\data_out_frame[17] [6]), 
            .I3(n30663), .O(n12_adj_3771));
    defparam i5_4_lut_adj_1292.LUT_INIT = 16'h9669;
    SB_LUT4 i13819_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n18326));
    defparam i13819_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1293 (.I0(\data_out_frame[17] [4]), .I1(n12_adj_3771), 
            .I2(n34111), .I3(n29848), .O(n29836));
    defparam i6_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i13820_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n18327));
    defparam i13820_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1027_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n4428));
    defparam mux_1027_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n13888));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h4406;
    SB_LUT4 i13821_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n18328));
    defparam i13821_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1294 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n34183));
    defparam i2_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1295 (.I0(\data_out_frame[9] [7]), .I1(n34183), 
            .I2(n33993), .I3(\data_out_frame[5] [3]), .O(n17128));
    defparam i3_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16661));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33914));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i13822_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n18329));
    defparam i13822_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13823_3_lut_4_lut (.I0(n8), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n18330));
    defparam i13823_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1298 (.I0(\data_out_frame[9] [6]), .I1(n33914), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[5] [2]), .O(n12_adj_3772));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1299 (.I0(n16661), .I1(n12_adj_3772), .I2(\data_out_frame[11] [7]), 
            .I3(\data_out_frame[5] [3]), .O(n34320));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1300 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n24905), .O(n33758));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1300.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_adj_1301 (.I0(\data_out_frame[14] [3]), .I1(n17128), 
            .I2(\data_out_frame[12] [2]), .I3(GND_net), .O(n34302));
    defparam i2_3_lut_adj_1301.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1302 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n24905), .O(n33767));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1302.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(n31_adj_3618), .I1(n24558), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n4_adj_3620));
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1304 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16406), .I3(GND_net), .O(n4_adj_3744));
    defparam i1_2_lut_3_lut_adj_1304.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_1305 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16406), .I3(GND_net), .O(n16417));
    defparam i1_2_lut_3_lut_adj_1305.LUT_INIT = 16'hf7f7;
    SB_LUT4 i28268_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n16406), .I3(GND_net), .O(n34510));
    defparam i28268_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i5_3_lut_adj_1306 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n14_adj_3773));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 equal_123_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_123_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_122_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3748));   // verilog/coms.v(154[7:23])
    defparam equal_122_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1307 (.I0(n33830), .I1(n34143), .I2(\data_out_frame[6] [2]), 
            .I3(\data_out_frame[6] [6]), .O(n15_adj_3774));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1308 (.I0(n15_adj_3774), .I1(\data_out_frame[13] [2]), 
            .I2(n14_adj_3773), .I3(\data_out_frame[13] [3]), .O(n17256));   // verilog/coms.v(72[16:27])
    defparam i8_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34066));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1310 (.I0(\data_out_frame[15] [6]), .I1(n34066), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[17] [7]), .O(n12_adj_3775));
    defparam i5_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1311 (.I0(n17256), .I1(n12_adj_3775), .I2(n34166), 
            .I3(n16983), .O(n34281));
    defparam i6_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i13812_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n18319));
    defparam i13812_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21076_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(\byte_transmit_counter[1] ), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[3]), 
            .O(n25566));
    defparam i21076_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n34057));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1313 (.I0(n33862), .I1(\data_out_frame[9] [3]), 
            .I2(n34057), .I3(\data_out_frame[11] [4]), .O(n34166));
    defparam i3_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1027_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n4427));
    defparam mux_1027_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1314 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n6_adj_3608));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16565));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34143));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i28251_3_lut_4_lut (.I0(n16280), .I1(n16410), .I2(LED_c), 
            .I3(n11748), .O(n34492));   // verilog/coms.v(148[5:9])
    defparam i28251_3_lut_4_lut.LUT_INIT = 16'he0ee;
    SB_LUT4 mux_1027_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n4426));
    defparam mux_1027_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17110));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34311));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1319 (.I0(\data_out_frame[10] [7]), .I1(n34311), 
            .I2(n17110), .I3(\data_out_frame[6] [3]), .O(n33830));
    defparam i3_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_out_frame[8] [7]), .I1(n33830), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3776));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35439 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n41758));
    defparam byte_transmit_counter_0__bdd_4_lut_35439.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1321 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(n6_adj_3776), .O(n1509));
    defparam i4_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1027_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n4425));
    defparam mux_1027_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n33792));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1323 (.I0(n33945), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[10] [5]), .I3(n34266), .O(n10_adj_3696));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n33788), .I3(GND_net), .O(n6_adj_3593));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1325 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33999));
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1027_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n24560), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16] [1]), .O(n4424));
    defparam mux_1027_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1326 (.I0(\data_out_frame[11] [2]), .I1(n33999), 
            .I2(\data_out_frame[9] [0]), .I3(\data_out_frame[9] [2]), .O(n16983));
    defparam i3_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n33790), .I3(GND_net), .O(n6_adj_3685));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17252));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1329 (.I0(\data_out_frame[7] [0]), .I1(n34166), 
            .I2(n17252), .I3(\data_out_frame[7] [1]), .O(n1515));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16803));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'h6666;
    SB_LUT4 i939_2_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1695));   // verilog/coms.v(69[16:27])
    defparam i939_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1331 (.I0(n7_adj_3694), .I1(n17040), .I2(n34199), 
            .I3(n1509), .O(n34299));
    defparam i4_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1332 (.I0(n33961), .I1(\data_out_frame[12] [3]), 
            .I2(n17128), .I3(GND_net), .O(n33820));
    defparam i2_3_lut_adj_1332.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1333 (.I0(n34299), .I1(\data_out_frame[16] [7]), 
            .I2(n1695), .I3(n16803), .O(n14_adj_3777));
    defparam i6_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1334 (.I0(\data_out_frame[14] [5]), .I1(n14_adj_3777), 
            .I2(n10_adj_3715), .I3(\data_out_frame[15] [1]), .O(n29828));
    defparam i7_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1335 (.I0(n17392), .I1(n33965), .I2(n34281), 
            .I3(\data_out_frame[18] [6]), .O(n22_adj_3778));
    defparam i9_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i2023_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(\FRAME_MATCHER.i [3]), .O(n10_adj_3607));
    defparam i2023_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i11_4_lut_adj_1336 (.I0(n15_adj_3714), .I1(n22_adj_3778), .I2(\data_out_frame[18] [5]), 
            .I3(n35783), .O(n24_adj_3779));
    defparam i11_4_lut_adj_1336.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1337 (.I0(n16668), .I1(n29879), .I2(\data_out_frame[18] [7]), 
            .I3(n14_adj_3698), .O(n23));
    defparam i10_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1338 (.I0(\data_out_frame[19] [4]), .I1(n16809), 
            .I2(\data_out_frame[19] [5]), .I3(n33883), .O(n10_adj_3780));
    defparam i4_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1339 (.I0(\data_out_frame[19] [1]), .I1(n10_adj_3780), 
            .I2(n23), .I3(n24_adj_3779), .O(n30703));
    defparam i5_4_lut_adj_1339.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1340 (.I0(n34102), .I1(n34233), .I2(\data_out_frame[18] [5]), 
            .I3(n17259), .O(n12_adj_3781));
    defparam i5_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1341 (.I0(n17085), .I1(n12_adj_3781), .I2(n34305), 
            .I3(n30703), .O(n30316));
    defparam i6_4_lut_adj_1341.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1342 (.I0(n30316), .I1(n30703), .I2(\data_out_frame[20] [7]), 
            .I3(n29828), .O(n12_adj_3782));
    defparam i5_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1343 (.I0(n16803), .I1(n12_adj_3782), .I2(n33795), 
            .I3(\data_out_frame[17] [0]), .O(n36123));
    defparam i6_4_lut_adj_1343.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34126));
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1345 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n34180));
    defparam i2_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34162));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1347 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33862));
    defparam i1_2_lut_adj_1347.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1348 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [1]), .O(n6_adj_3571));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1349 (.I0(\FRAME_MATCHER.state[0] ), .I1(n16285), 
            .I2(n16410), .I3(\FRAME_MATCHER.state [3]), .O(n35990));   // verilog/coms.v(195[5:24])
    defparam i2_3_lut_4_lut_adj_1349.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(\FRAME_MATCHER.state[0] ), .I1(n16285), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n16280));   // verilog/coms.v(195[5:24])
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17002));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1352 (.I0(n34278), .I1(\data_out_frame[11] [4]), 
            .I2(n33862), .I3(GND_net), .O(n33935));
    defparam i2_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i908_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1664));   // verilog/coms.v(83[17:28])
    defparam i908_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in[1] [1]), .I1(n10_adj_3622), .I2(\data_in[2] [7]), 
            .I3(\data_in[3] [0]), .O(n15_adj_3605));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i3_4_lut_adj_1353 (.I0(\data_out_frame[5] [3]), .I1(n34180), 
            .I2(n33880), .I3(n33862), .O(n17265));
    defparam i3_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1354 (.I0(n33935), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[9] [2]), .I3(n33948), .O(n34199));
    defparam i3_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 n41758_bdd_4_lut (.I0(n41758), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n41761));
    defparam n41758_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33875));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34287));
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3783));
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1358 (.I0(n34177), .I1(\data_out_frame[8] [0]), 
            .I2(n34287), .I3(n6_adj_3783), .O(n33961));
    defparam i4_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1359 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n8_adj_3784));   // verilog/coms.v(83[17:28])
    defparam i3_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1360 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3785));   // verilog/coms.v(83[17:28])
    defparam i2_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1361 (.I0(n33908), .I1(\data_out_frame[9] [6]), 
            .I2(n7_adj_3785), .I3(n8_adj_3784), .O(n17465));   // verilog/coms.v(83[17:28])
    defparam i2_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1362 (.I0(n17465), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[12] [2]), .I3(n33961), .O(n34060));
    defparam i3_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n33807));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i13813_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n18320));
    defparam i13813_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1364 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17091));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_1364.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_adj_1365 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[0] [6]), .I3(n4_adj_3598), .O(n6_adj_3573));   // verilog/coms.v(68[16:69])
    defparam i2_2_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i13911_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n18418));
    defparam i13911_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13910_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n18417));
    defparam i13910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35434 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n41752));
    defparam byte_transmit_counter_0__bdd_4_lut_35434.LUT_INIT = 16'he4aa;
    SB_LUT4 i13814_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n18321));
    defparam i13814_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16812));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h6666;
    SB_LUT4 i13608_3_lut_4_lut (.I0(n4025), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17568), .I3(\data_out_frame[0] [2]), .O(n18115));
    defparam i13608_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 n41752_bdd_4_lut (.I0(n41752), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n41755));
    defparam n41752_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35429 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n41746));
    defparam byte_transmit_counter_0__bdd_4_lut_35429.LUT_INIT = 16'he4aa;
    SB_LUT4 i13909_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n18416));
    defparam i13909_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(n33929), .I3(\data_in_frame[3] [2]), .O(n34123));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 n41746_bdd_4_lut (.I0(n41746), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n41749));
    defparam n41746_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13609_3_lut_4_lut (.I0(n4025), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17568), .I3(\data_out_frame[0] [3]), .O(n18116));
    defparam i13609_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(n4_adj_3598), .I1(n34099), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n30692));
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1369 (.I0(n16066), .I1(n16812), .I2(n17259), 
            .I3(n16989), .O(n34114));
    defparam i3_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i13610_3_lut_4_lut (.I0(n4025), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17568), .I3(\data_out_frame[0] [4]), .O(n18117));
    defparam i13610_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i13908_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n18415));
    defparam i13908_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13907_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n18414));
    defparam i13907_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1370 (.I0(\data_out_frame[18] [6]), .I1(n34114), 
            .I2(GND_net), .I3(GND_net), .O(n34115));
    defparam i1_2_lut_adj_1370.LUT_INIT = 16'h9999;
    SB_LUT4 select_337_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3664));
    defparam select_337_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3662));
    defparam select_337_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3660));
    defparam select_337_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3659));
    defparam select_337_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3658));
    defparam select_337_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3657));
    defparam select_337_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3656));
    defparam select_337_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3655));
    defparam select_337_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3654));
    defparam select_337_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3653));
    defparam select_337_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3652));
    defparam select_337_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3651));
    defparam select_337_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3650));
    defparam select_337_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3649));
    defparam select_337_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3648));
    defparam select_337_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3647));
    defparam select_337_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3646));
    defparam select_337_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3645));
    defparam select_337_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3644));
    defparam select_337_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3643));
    defparam select_337_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3642));
    defparam select_337_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3641));
    defparam select_337_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3640));
    defparam select_337_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13815_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n18322));
    defparam i13815_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_337_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3639));
    defparam select_337_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3638));
    defparam select_337_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13906_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n18413));
    defparam i13906_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13754_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n18261));
    defparam i13754_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13913_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n18420));
    defparam i13913_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_337_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3637));
    defparam select_337_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3636));
    defparam select_337_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3635));
    defparam select_337_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3634));
    defparam select_337_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_337_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3633));
    defparam select_337_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13755_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n18262));
    defparam i13755_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1371 (.I0(n31), .I1(n31_adj_3618), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n25604), .O(n7_adj_3592));
    defparam i2_2_lut_4_lut_adj_1371.LUT_INIT = 16'hffca;
    SB_LUT4 i13756_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n18263));
    defparam i13756_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13757_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n18264));
    defparam i13757_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13758_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n18265));
    defparam i13758_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13912_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n18419));
    defparam i13912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35424 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n41740));
    defparam byte_transmit_counter_0__bdd_4_lut_35424.LUT_INIT = 16'he4aa;
    SB_LUT4 i13898_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18405));
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13759_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n18266));
    defparam i13759_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n41740_bdd_4_lut (.I0(n41740), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n41743));
    defparam n41740_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13760_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n18267));
    defparam i13760_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13761_3_lut_4_lut (.I0(n8), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n18268));
    defparam i13761_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut_adj_1372 (.I0(n19473), .I1(n9818), .I2(n2236[0]), 
            .I3(\byte_transmit_counter[0] ), .O(n18521));
    defparam i1_4_lut_4_lut_adj_1372.LUT_INIT = 16'hea40;
    SB_LUT4 i5_3_lut_4_lut_adj_1373 (.I0(\data_in_frame[16] [3]), .I1(n30661), 
            .I2(n10_adj_3586), .I3(\data_in_frame[20] [7]), .O(n34944));
    defparam i5_3_lut_4_lut_adj_1373.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_4_lut_adj_1374 (.I0(n19473), .I1(n9818), .I2(n2236[6]), 
            .I3(byte_transmit_counter[6]), .O(n18543));
    defparam i1_4_lut_4_lut_adj_1374.LUT_INIT = 16'hea40;
    SB_LUT4 i13746_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n18253));
    defparam i13746_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13747_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n18254));
    defparam i13747_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13748_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n18255));
    defparam i13748_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13749_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n18256));
    defparam i13749_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(n30677), .I1(\data_in_frame[17] [7]), 
            .I2(n35995), .I3(n29826), .O(n6_adj_3578));
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'h9669;
    SB_LUT4 select_337_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2540), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3632));
    defparam select_337_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[16] [1]), 
            .I2(n30677), .I3(GND_net), .O(n6_adj_3587));
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'h9696;
    SB_LUT4 i13750_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n18257));
    defparam i13750_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_35419 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n41734));
    defparam byte_transmit_counter_0__bdd_4_lut_35419.LUT_INIT = 16'he4aa;
    SB_LUT4 n41734_bdd_4_lut (.I0(n41734), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n41737));
    defparam n41734_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35532 (.I0(\byte_transmit_counter[1] ), 
            .I1(n37267), .I2(n37268), .I3(byte_transmit_counter[2]), .O(n41728));
    defparam byte_transmit_counter_1__bdd_4_lut_35532.LUT_INIT = 16'he4aa;
    SB_LUT4 n41728_bdd_4_lut (.I0(n41728), .I1(n37337), .I2(n37336), .I3(byte_transmit_counter[2]), 
            .O(n41731));
    defparam n41728_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13900_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18407));
    defparam i13900_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13816_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n18323));
    defparam i13816_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13899_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18406));
    defparam i13899_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13751_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n18258));
    defparam i13751_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13752_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n18259));
    defparam i13752_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13905_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18412));
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13753_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n18260));
    defparam i13753_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13904_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18411));
    defparam i13904_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13903_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18410));
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13902_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18409));
    defparam i13902_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1377 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[7] [6]), .I3(GND_net), .O(n33990));
    defparam i1_2_lut_3_lut_adj_1377.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[7] [5]), 
            .I2(\data_in_frame[7] [4]), .I3(GND_net), .O(n34153));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1379 (.I0(n33943), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[7] [3]), .I3(Kp_23__N_871), .O(n35103));
    defparam i2_3_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 equal_109_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3594));   // verilog/coms.v(154[7:23])
    defparam equal_109_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13901_3_lut_4_lut (.I0(n8_adj_3740), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18408));
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_108_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3576));   // verilog/coms.v(154[7:23])
    defparam equal_108_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i13784_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n18291));
    defparam i13784_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13785_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n18292));
    defparam i13785_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13778_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n18285));
    defparam i13778_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13779_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n18286));
    defparam i13779_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13817_3_lut_4_lut (.I0(n8_adj_3576), .I1(n33767), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n18324));
    defparam i13817_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13780_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n18287));
    defparam i13780_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13781_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n18288));
    defparam i13781_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13782_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n18289));
    defparam i13782_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13783_3_lut_4_lut (.I0(n8_adj_3726), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n18290));
    defparam i13783_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13895_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18402));
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37305), .I3(n37304), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13896_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18403));
    defparam i13896_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13894_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18401));
    defparam i13894_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13897_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18404));
    defparam i13897_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13890_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18397));
    defparam i13890_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37302), .I3(n37301), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13891_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18398));
    defparam i13891_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37299), .I3(n37298), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13892_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18399));
    defparam i13892_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_2_lut_3_lut (.I0(n33943), .I1(n4_adj_3598), .I2(n34099), 
            .I3(GND_net), .O(n12_adj_3570));   // verilog/coms.v(77[16:35])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13893_3_lut_4_lut (.I0(n8_adj_3748), .I1(n33776), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18400));
    defparam i13893_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37296), .I3(n37295), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i2_3_lut_4_lut_adj_1380 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n16466), .I3(\FRAME_MATCHER.i [4]), .O(n16256));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1380.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1381 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n24905), .O(n33776));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1381.LUT_INIT = 16'hefff;
    SB_LUT4 i13387_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n17894));
    defparam i13387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13739_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n18246));
    defparam i13739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13740_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n18247));
    defparam i13740_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(\data_in_frame[15] [7]), .I1(n35103), 
            .I2(n10_adj_3569), .I3(\data_in_frame[9] [5]), .O(n34329));
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37287), .I3(n41731), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i2_3_lut_4_lut_adj_1383 (.I0(Kp_23__N_868), .I1(Kp_23__N_871), 
            .I2(\data_in_frame[5] [0]), .I3(n29784), .O(n29900));
    defparam i2_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37290), .I3(n37289), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n37293), .I3(n37292), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13741_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n18248));
    defparam i13741_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1384 (.I0(n16824), .I1(n30393), .I2(n17187), 
            .I3(\data_in_frame[13] [4]), .O(n30710));
    defparam i2_3_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i13742_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n18249));
    defparam i13742_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13743_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n18250));
    defparam i13743_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13744_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n18251));
    defparam i13744_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13745_3_lut_4_lut (.I0(n8_adj_3594), .I1(n33758), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n18252));
    defparam i13745_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1385 (.I0(n33986), .I1(n34221), .I2(\data_in_frame[6] [3]), 
            .I3(\data_in_frame[10] [7]), .O(n17170));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(\data_in_frame[14] [0]), .I1(n33943), 
            .I2(\data_in_frame[11] [4]), .I3(n35254), .O(n6_adj_3566));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    uart_tx tx (.n18509(n18509), .r_SM_Main({r_SM_Main}), .clk32MHz(clk32MHz), 
            .n17827(n17827), .r_Bit_Index({r_Bit_Index}), .n17830(n17830), 
            .\r_SM_Main_2__N_3298[0] (\r_SM_Main_2__N_3298[0] ), .GND_net(GND_net), 
            .tx_data({tx_data}), .\r_SM_Main_2__N_3295[1] (\r_SM_Main_2__N_3295[1] ), 
            .n17625(n17625), .n17748(n17748), .n4706(n4706), .n17989(n17989), 
            .VCC_net(VCC_net), .tx_active(tx_active), .tx_o(tx_o), .tx_enable(tx_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.n18539(n18539), .VCC_net(VCC_net), .r_Clock_Count({Open_14, 
            Open_15, Open_16, Open_17, Open_18, \r_Clock_Count[2] , 
            \r_Clock_Count[1] , \r_Clock_Count[0] }), .clk32MHz(clk32MHz), 
            .n17836(n17836), .r_Bit_Index({r_Bit_Index_adj_10}), .n17833(n17833), 
            .r_SM_Main({\r_SM_Main[2]_adj_7 , \r_SM_Main[1]_adj_6 , Open_19}), 
            .n2346(n2346), .GND_net(GND_net), .r_Rx_Data(r_Rx_Data), .PIN_13_N_106(PIN_13_N_106), 
            .\r_Clock_Count[6] (\r_Clock_Count[6] ), .\r_Clock_Count[4] (\r_Clock_Count[4] ), 
            .n16429(n16429), .n4(n4), .n35922(n35922), .n4684(n4684), 
            .n17619(n17619), .n17746(n17746), .n17931(n17931), .n17936(n17936), 
            .n17942(n17942), .n17980(n17980), .n17992(n17992), .n18003(n18003), 
            .rx_data({rx_data}), .n33396(n33396), .rx_data_ready(rx_data_ready), 
            .n220(n220), .n222(n222), .n224(n224), .n225(n225), .n226(n226), 
            .n24632(n24632), .n4_adj_1(n4_adj_8), .n4_adj_2(n4_adj_9), 
            .n16424(n16424), .n17843(n17843), .n17842(n17842), .n17841(n17841), 
            .n17840(n17840), .n17839(n17839), .n17838(n17838), .n17837(n17837), 
            .n17522(n17522)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n18509, r_SM_Main, clk32MHz, n17827, r_Bit_Index, 
            n17830, \r_SM_Main_2__N_3298[0] , GND_net, tx_data, \r_SM_Main_2__N_3295[1] , 
            n17625, n17748, n4706, n17989, VCC_net, tx_active, tx_o, 
            tx_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18509;
    output [2:0]r_SM_Main;
    input clk32MHz;
    input n17827;
    output [2:0]r_Bit_Index;
    input n17830;
    input \r_SM_Main_2__N_3298[0] ;
    input GND_net;
    input [7:0]tx_data;
    output \r_SM_Main_2__N_3295[1] ;
    output n17625;
    output n17748;
    output n4706;
    input n17989;
    input VCC_net;
    output tx_active;
    output tx_o;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [8:0]n312;
    
    wire n17604;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n17731, n104, n14127;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n27543, n27542, n25370, n35491, n10, n19975, n27541, 
        n27540, n27539, n27538, n27537, n27536, n17910, n20001, 
        n10_adj_3565, n37306, n37307, n37370, n37369, n42264, n11836, 
        n41770, o_Tx_Serial_N_3326, n12, n17535;
    
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n18509));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17827));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17830));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .E(n17604), 
            .D(n312[8]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .E(n17604), 
            .D(n312[7]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .E(n17604), 
            .D(n312[6]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .E(n17604), 
            .D(n312[5]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .E(n17604), 
            .D(n312[4]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .E(n17604), 
            .D(n312[3]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .E(n17604), 
            .D(n312[2]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .E(n17604), 
            .D(n312[1]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3298[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n27543), .O(n312[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n27542), .O(n312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n25370));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3295[1] ), .O(n17625));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i13241_3_lut (.I0(n17625), .I1(n25370), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17748));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13241_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1253_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4706));   // verilog/uart_tx.v(98[36:51])
    defparam i1253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_59_9 (.CI(n27542), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n27543));
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[2]), .O(n35491));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[6]), .I2(n35491), 
            .I3(r_Clock_Count[7]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[5]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3295[1] ));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_862 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3295[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n19975));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h8888;
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n27541), .O(n312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n27541), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n27542));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n27540), .O(n312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n27540), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n27541));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n27539), .O(n312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n27539), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n27540));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n27538), .O(n312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n27538), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n27539));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27537), .O(n312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n27537), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27538));
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17989));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27536), .O(n312[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n27536), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27537));
    SB_LUT4 add_59_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n312[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n27536));
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n17910));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n20001));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n10_adj_3565));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(n17604), 
            .D(n312[0]), .R(n17731));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n14127), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30986_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n37306));
    defparam i30986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30987_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n37307));
    defparam i30987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31050_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n37370));
    defparam i31050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31049_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n37369));
    defparam i31049_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n42264));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(n11836), .I2(\r_SM_Main_2__N_3295[1] ), 
            .I3(r_SM_Main[0]), .O(n17910));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_4_lut_4_lut_adj_863 (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3295[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n17731));
    defparam i1_4_lut_4_lut_adj_863.LUT_INIT = 16'h4445;
    SB_LUT4 i15444_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17604));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i15444_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3295[1] ), .O(n42264));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n37369), 
            .I2(n37370), .I3(r_Bit_Index[2]), .O(n41770));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n41770_bdd_4_lut (.I0(n41770), .I1(n37307), .I2(n37306), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3326));
    defparam n41770_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i26_3_lut (.I0(o_Tx_Serial_N_3326), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10_adj_3565));
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_4_lut_adj_864 (.I0(n104), .I1(n17604), .I2(r_SM_Main[1]), 
            .I3(n19975), .O(n17535));
    defparam i2_4_lut_adj_864.LUT_INIT = 16'hc808;
    SB_LUT4 i15498_3_lut (.I0(n17535), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n20001));   // verilog/uart_tx.v(31[16:25])
    defparam i15498_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i7438_4_lut (.I0(\r_SM_Main_2__N_3298[0] ), .I1(n25370), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3295[1] ), .O(n11836));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7438_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3298[0] ), .O(n14127));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n18539, VCC_net, r_Clock_Count, clk32MHz, n17836, 
            r_Bit_Index, n17833, r_SM_Main, n2346, GND_net, r_Rx_Data, 
            PIN_13_N_106, \r_Clock_Count[6] , \r_Clock_Count[4] , n16429, 
            n4, n35922, n4684, n17619, n17746, n17931, n17936, 
            n17942, n17980, n17992, n18003, rx_data, n33396, rx_data_ready, 
            n220, n222, n224, n225, n226, n24632, n4_adj_1, n4_adj_2, 
            n16424, n17843, n17842, n17841, n17840, n17839, n17838, 
            n17837, n17522) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18539;
    input VCC_net;
    output [7:0]r_Clock_Count;
    input clk32MHz;
    input n17836;
    output [2:0]r_Bit_Index;
    input n17833;
    output [2:0]r_SM_Main;
    output n2346;
    input GND_net;
    output r_Rx_Data;
    input PIN_13_N_106;
    output \r_Clock_Count[6] ;
    output \r_Clock_Count[4] ;
    output n16429;
    output n4;
    output n35922;
    output n4684;
    output n17619;
    output n17746;
    input n17931;
    input n17936;
    input n17942;
    input n17980;
    input n17992;
    input n18003;
    output [7:0]rx_data;
    input n33396;
    output rx_data_ready;
    output n220;
    output n222;
    output n224;
    output n225;
    output n226;
    output n24632;
    output n4_adj_1;
    output n4_adj_2;
    output n16424;
    input n17843;
    input n17842;
    input n17841;
    input n17840;
    input n17839;
    input n17838;
    input n17837;
    output n17522;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n25556;
    wire [2:0]r_SM_Main_2__N_3224;
    
    wire n33744, n17555;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n39034, n39033, r_Rx_Data_R, n3;
    wire [7:0]r_Clock_Count_c;   // verilog/uart_rx.v(32[17:30])
    
    wire n24, n33743, n44, n16377, n46, n36246, n6, n16265, 
        n4_adj_3561, n19, n4_adj_3562, n33196;
    wire [31:0]n194;
    
    wire n32, n26, n18014, n25159, n27535, n27534, n27533, n17901, 
        n27532, n27531, n27530, n27529, n1, n25444;
    
    SB_DFFE r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18539));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17836));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17833));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n25556));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3224[2]), 
            .R(n33744));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1068_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n17555));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1068_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32873_2_lut (.I0(r_SM_Main_2__N_3224[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39034));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32873_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35353_4_lut (.I0(r_SM_Main[2]), .I1(n39033), .I2(n39034), 
            .I3(r_SM_Main[1]), .O(n25556));
    defparam i35353_4_lut.LUT_INIT = 16'h0511;
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_106));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i2_3_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[0]), 
            .I3(GND_net), .O(n3));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count_c[3]), .I1(n3), .I2(GND_net), 
            .I3(GND_net), .O(n24));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_850 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33743));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_850.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count_c[7]), .I1(n44), .I2(n33743), 
            .I3(n24), .O(n16377));
    defparam i3_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_adj_851 (.I0(r_Clock_Count_c[5]), .I1(\r_Clock_Count[6] ), 
            .I2(\r_Clock_Count[4] ), .I3(GND_net), .O(n44));
    defparam i2_3_lut_adj_851.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_852 (.I0(r_Clock_Count[0]), .I1(n46), .I2(r_Clock_Count[2]), 
            .I3(r_Clock_Count[1]), .O(n36246));
    defparam i3_4_lut_adj_852.LUT_INIT = 16'hdfff;
    SB_LUT4 i2_2_lut (.I0(n36246), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i28209_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n2346));
    defparam i28209_4_lut.LUT_INIT = 16'hbaaa;
    SB_LUT4 i3_4_lut_adj_853 (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_3224[2]), .O(n16265));
    defparam i3_4_lut_adj_853.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_854 (.I0(r_Bit_Index[0]), .I1(n16265), .I2(GND_net), 
            .I3(GND_net), .O(n16429));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_854.LUT_INIT = 16'heeee;
    SB_LUT4 equal_140_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_140_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(n2346), .I1(n16377), .I2(n36246), .I3(n4_adj_3561), 
            .O(n35922));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_4_lut (.I0(n36246), .I1(n16377), .I2(r_SM_Main[1]), .I3(r_SM_Main_c[0]), 
            .O(n19));
    defparam i1_4_lut.LUT_INIT = 16'hcecc;
    SB_LUT4 i1_4_lut_adj_855 (.I0(n19), .I1(r_Clock_Count_c[7]), .I2(n4_adj_3562), 
            .I3(n2346), .O(n33196));
    defparam i1_4_lut_adj_855.LUT_INIT = 16'heca0;
    SB_LUT4 i34654_4_lut (.I0(n194[5]), .I1(r_Clock_Count_c[5]), .I2(n2346), 
            .I3(n32), .O(n26));
    defparam i34654_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_4_lut_adj_856 (.I0(n35922), .I1(r_Clock_Count_c[3]), .I2(n194[3]), 
            .I3(n2346), .O(n18014));
    defparam i1_4_lut_adj_856.LUT_INIT = 16'h4450;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_Clock_Count_c[7]), .I1(n44), .I2(r_Clock_Count_c[3]), 
            .I3(GND_net), .O(n46));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(n36246), 
            .I3(n16377), .O(n32));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h00bf;
    SB_LUT4 i1_2_lut_3_lut_adj_857 (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), 
            .I2(r_SM_Main[2]), .I3(GND_net), .O(n4_adj_3561));
    defparam i1_2_lut_3_lut_adj_857.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1231_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4684));   // verilog/uart_rx.v(102[36:51])
    defparam i1231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_858 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n25159));
    defparam i2_3_lut_adj_858.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_859 (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3224[2]), 
            .I2(r_SM_Main_c[0]), .I3(r_SM_Main[1]), .O(n17619));
    defparam i2_4_lut_adj_859.LUT_INIT = 16'h0405;
    SB_LUT4 i13239_3_lut (.I0(n17619), .I1(n25159), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17746));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13239_3_lut.LUT_INIT = 16'h8a8a;
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n17931));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17936));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count_c[3]), .C(clk32MHz), .D(n18014));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(\r_Clock_Count[4] ), .C(clk32MHz), .D(n17942));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count_c[5]), .C(clk32MHz), .D(n26));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(clk32MHz), .D(n17980));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count_c[7]), .C(clk32MHz), .D(n33196));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17992));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18003));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n33396));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(n17555), .I1(r_Clock_Count_c[7]), .I2(GND_net), 
            .I3(n27535), .O(n4_adj_3562)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(\r_Clock_Count[6] ), .I2(GND_net), 
            .I3(n27534), .O(n220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n27534), .I0(\r_Clock_Count[6] ), .I1(GND_net), 
            .CO(n27535));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count_c[5]), .I2(GND_net), 
            .I3(n27533), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n27533), .I0(r_Clock_Count_c[5]), .I1(GND_net), 
            .CO(n27534));
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n17901));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(\r_Clock_Count[4] ), .I2(GND_net), 
            .I3(n27532), .O(n222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_6 (.CI(n27532), .I0(\r_Clock_Count[4] ), .I1(GND_net), 
            .CO(n27533));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count_c[3]), .I2(GND_net), 
            .I3(n27531), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n27531), .I0(r_Clock_Count_c[3]), .I1(GND_net), 
            .CO(n27532));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27530), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n27530), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27531));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27529), .O(n225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n27529), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27530));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n27529));
    SB_LUT4 i20147_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n24632));
    defparam i20147_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_136_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_136_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_138_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_138_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_860 (.I0(n16265), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n16424));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17843));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17842));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17841));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17840));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17839));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17838));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17837));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i35360_2_lut_3_lut (.I0(r_SM_Main_c[0]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(GND_net), .O(n33744));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i35360_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i20691_2_lut_3_lut_4_lut (.I0(r_Clock_Count_c[7]), .I1(n44), 
            .I2(r_Clock_Count_c[3]), .I3(n3), .O(r_SM_Main_2__N_3224[2]));
    defparam i20691_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_c[0]), 
            .I3(r_SM_Main_2__N_3224[2]), .O(n17522));
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_4_lut (.I0(n3), .I1(n46), 
            .I2(r_SM_Main_c[0]), .I3(r_Rx_Data), .O(n1));
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_4_lut.LUT_INIT = 16'hd0df;
    SB_LUT4 i33089_3_lut_4_lut (.I0(n3), .I1(n46), .I2(r_Rx_Data), .I3(r_SM_Main_c[0]), 
            .O(n39033));
    defparam i33089_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n25159), .I1(r_SM_Main_2__N_3224[2]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n25444));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i1_4_lut_adj_861 (.I0(r_SM_Main[2]), .I1(n1), .I2(n25444), 
            .I3(r_SM_Main[1]), .O(n17901));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_861.LUT_INIT = 16'h0544;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n2731, encoder0_position, GND_net, 
            n18466, clk32MHz, n18467, n18468, n18469, n18470, n18471, 
            n18451, n18452, n18472, n18473, n18462, n18463, n18464, 
            n18465, n18453, n18454, n18455, n18456, n18457, n18458, 
            n18459, n18460, n18461, data_o, count_enable, n17897, 
            n18498, n34976, reg_B, n17900, PIN_2_c_0, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2731;
    output [23:0]encoder0_position;
    input GND_net;
    input n18466;
    input clk32MHz;
    input n18467;
    input n18468;
    input n18469;
    input n18470;
    input n18471;
    input n18451;
    input n18452;
    input n18472;
    input n18473;
    input n18462;
    input n18463;
    input n18464;
    input n18465;
    input n18453;
    input n18454;
    input n18455;
    input n18456;
    input n18457;
    input n18458;
    input n18459;
    input n18460;
    input n18461;
    output [1:0]data_o;
    output count_enable;
    input n17897;
    input n18498;
    output n34976;
    output [1:0]reg_B;
    input n17900;
    input PIN_2_c_0;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n2727, n27551, n27552, n27550, n27549, n27548, n27547, 
        n27546, B_delayed, A_delayed, n27545, count_direction, n27544, 
        n27567, n27566, n27565, n27564, n27563, n27562, n27561, 
        n27560, n27559, n27558, n27557, n27556, n27555, n27554, 
        n27553;
    
    SB_LUT4 add_619_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2727), 
            .I3(n27551), .O(n2731[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_9 (.CI(n27551), .I0(encoder0_position[7]), .I1(n2727), 
            .CO(n27552));
    SB_LUT4 add_619_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2727), 
            .I3(n27550), .O(n2731[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_8 (.CI(n27550), .I0(encoder0_position[6]), .I1(n2727), 
            .CO(n27551));
    SB_LUT4 add_619_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2727), 
            .I3(n27549), .O(n2731[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_7 (.CI(n27549), .I0(encoder0_position[5]), .I1(n2727), 
            .CO(n27550));
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n18466));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n18467));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n18468));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n18469));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n18470));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n18471));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n18451));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n18452));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n18472));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n18473));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n18462));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n18463));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n18464));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n18465));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n18453));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n18454));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n18455));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n18456));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n18457));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n18458));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n18459));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n18460));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n18461));   // quad.v(35[10] 41[6])
    SB_LUT4 add_619_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2727), 
            .I3(n27548), .O(n2731[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_6 (.CI(n27548), .I0(encoder0_position[4]), .I1(n2727), 
            .CO(n27549));
    SB_LUT4 add_619_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2727), 
            .I3(n27547), .O(n2731[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_5 (.CI(n27547), .I0(encoder0_position[3]), .I1(n2727), 
            .CO(n27548));
    SB_LUT4 add_619_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2727), 
            .I3(n27546), .O(n2731[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_619_4 (.CI(n27546), .I0(encoder0_position[2]), .I1(n2727), 
            .CO(n27547));
    SB_LUT4 add_619_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2727), 
            .I3(n27545), .O(n2731[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_619_3 (.CI(n27545), .I0(encoder0_position[1]), .I1(n2727), 
            .CO(n27546));
    SB_LUT4 add_619_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27544), .O(n2731[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_2 (.CI(n27544), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27545));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_619_1 (.CI(GND_net), .I0(n2727), .I1(n2727), .CO(n27544));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17897));   // quad.v(35[10] 41[6])
    SB_LUT4 add_619_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2727), 
            .I3(n27567), .O(n2731[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_619_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2727), 
            .I3(n27566), .O(n2731[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_24 (.CI(n27566), .I0(encoder0_position[22]), .I1(n2727), 
            .CO(n27567));
    SB_LUT4 add_619_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2727), 
            .I3(n27565), .O(n2731[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_23 (.CI(n27565), .I0(encoder0_position[21]), .I1(n2727), 
            .CO(n27566));
    SB_LUT4 add_619_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2727), 
            .I3(n27564), .O(n2731[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_22 (.CI(n27564), .I0(encoder0_position[20]), .I1(n2727), 
            .CO(n27565));
    SB_LUT4 add_619_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2727), 
            .I3(n27563), .O(n2731[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_21 (.CI(n27563), .I0(encoder0_position[19]), .I1(n2727), 
            .CO(n27564));
    SB_LUT4 add_619_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2727), 
            .I3(n27562), .O(n2731[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_20 (.CI(n27562), .I0(encoder0_position[18]), .I1(n2727), 
            .CO(n27563));
    SB_LUT4 add_619_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2727), 
            .I3(n27561), .O(n2731[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_19 (.CI(n27561), .I0(encoder0_position[17]), .I1(n2727), 
            .CO(n27562));
    SB_LUT4 add_619_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2727), 
            .I3(n27560), .O(n2731[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_18 (.CI(n27560), .I0(encoder0_position[16]), .I1(n2727), 
            .CO(n27561));
    SB_LUT4 add_619_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2727), 
            .I3(n27559), .O(n2731[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_17 (.CI(n27559), .I0(encoder0_position[15]), .I1(n2727), 
            .CO(n27560));
    SB_LUT4 add_619_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2727), 
            .I3(n27558), .O(n2731[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_16 (.CI(n27558), .I0(encoder0_position[14]), .I1(n2727), 
            .CO(n27559));
    SB_LUT4 add_619_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2727), 
            .I3(n27557), .O(n2731[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_15 (.CI(n27557), .I0(encoder0_position[13]), .I1(n2727), 
            .CO(n27558));
    SB_LUT4 add_619_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2727), 
            .I3(n27556), .O(n2731[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_14 (.CI(n27556), .I0(encoder0_position[12]), .I1(n2727), 
            .CO(n27557));
    SB_LUT4 add_619_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2727), 
            .I3(n27555), .O(n2731[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_13 (.CI(n27555), .I0(encoder0_position[11]), .I1(n2727), 
            .CO(n27556));
    SB_LUT4 add_619_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2727), 
            .I3(n27554), .O(n2731[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_12 (.CI(n27554), .I0(encoder0_position[10]), .I1(n2727), 
            .CO(n27555));
    SB_LUT4 add_619_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2727), 
            .I3(n27553), .O(n2731[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_11 (.CI(n27553), .I0(encoder0_position[9]), .I1(n2727), 
            .CO(n27554));
    SB_LUT4 add_619_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2727), 
            .I3(n27552), .O(n2731[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_619_10 (.CI(n27552), .I0(encoder0_position[8]), .I1(n2727), 
            .CO(n27553));
    SB_LUT4 i894_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2727));   // quad.v(37[5] 40[8])
    defparam i894_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n18498(n18498), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .n34976(n34976), .GND_net(GND_net), .reg_B({reg_B}), 
            .n17900(n17900), .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18498, data_o, clk32MHz, n34976, GND_net, 
            reg_B, n17900, PIN_2_c_0, PIN_1_c_1) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18498;
    output [1:0]data_o;
    input clk32MHz;
    output n34976;
    input GND_net;
    output [1:0]reg_B;
    input n17900;
    input PIN_2_c_0;
    input PIN_1_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3459;
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18498));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n34976));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34976), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22817_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22817_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1140__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17900));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1140__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1140__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i22826_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22826_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22819_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22819_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (VCC_net, PIN_19_c_0, CLK_c, 
            \half_duty_new[0] , n18513, \half_duty[0][2] , n18514, \half_duty[0][3] , 
            n18515, \half_duty[0][4] , n18517, \half_duty[0][6] , n18518, 
            \half_duty[0][7] , n18512, \half_duty[0][1] , GND_net, n1035, 
            n17932, \half_duty[0][0] , \half_duty_new[1] , \half_duty_new[2] , 
            \half_duty_new[3] , \half_duty_new[4] , \half_duty_new[6] , 
            \half_duty_new[7] , pwm_setpoint) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input VCC_net;
    output PIN_19_c_0;
    input CLK_c;
    output \half_duty_new[0] ;
    input n18513;
    output \half_duty[0][2] ;
    input n18514;
    output \half_duty[0][3] ;
    input n18515;
    output \half_duty[0][4] ;
    input n18517;
    output \half_duty[0][6] ;
    input n18518;
    output \half_duty[0][7] ;
    input n18512;
    output \half_duty[0][1] ;
    input GND_net;
    output n1035;
    input n17932;
    output \half_duty[0][0] ;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input [22:0]pwm_setpoint;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n10, n27487;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire pwm_out_0__N_557, n17544;
    wire [9:0]half_duty_new_9__N_639;
    
    wire n23054;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n27488, n40977, n27486;
    wire [10:0]n49;
    
    wire pause_counter_0__N_587, n8;
    wire [10:0]pwm_out_0__N_562;
    
    wire n27485, n40979, n27484, n40981, n27483, n27489, pwm_out_0__N_561, 
        n5, n27482, n34475, pause_counter_0, n4, n27481, n3, n27480, 
        n2, n27479, n28353, n28352, n28351, n28350, n28349, n1, 
        n28348, n28347, n28346, n28345;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n37057, n12, n18, n19, n28344, n20, n13, n22, n37176, 
        n14, n18_adj_3560, n16, n17, n15;
    wire [22:0]n5649;
    
    wire n27756, n27755, n27754, n27753, n27752, n27751, n27750, 
        n27749, n27748, n27747, n27746, n27745, n27744, n27743, 
        n27742, n27741, n27740, n27739, n27738, n27737, n27736, 
        n27735, n27734, n27733, n27732, n27731, n27730, n27729, 
        n27728, n27727, n27726, n27725, n27724, n27723, n27722, 
        n27721, n27720, n27719, n27718, n27717, n27716, n27715, 
        n27714;
    
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n27487), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n17544), .D(pwm_out_0__N_557));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_639[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n18513));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n18514));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n18515));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0] [5]), .C(CLK_c), .D(n23054));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n18517));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n18518));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n18512));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_20_11 (.CI(n27487), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27488));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n27486), .O(n40977)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_DFFESR count_0__1139__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[10]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_10 (.CI(n27486), .I0(GND_net), .I1(VCC_net), 
            .CO(n27487));
    SB_DFFESR count_0__1139__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[9]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[8]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[7]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[6]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_562[7]), 
            .I3(n27485), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_DFFESR count_0__1139__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[5]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[4]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[3]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[2]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1139__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[1]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_9 (.CI(n27485), .I0(GND_net), .I1(pwm_out_0__N_562[7]), 
            .CO(n27486));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_562[6]), 
            .I3(n27484), .O(n40979)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n27484), .I0(VCC_net), .I1(pwm_out_0__N_562[6]), 
            .CO(n27485));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_562[5]), 
            .I3(n27483), .O(n40981)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_13 (.CI(n27489), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_561));
    SB_DFFESR count_0__1139__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_587), 
            .D(n49[0]), .R(n1035));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_7 (.CI(n27483), .I0(GND_net), .I1(pwm_out_0__N_562[5]), 
            .CO(n27484));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_562[4]), 
            .I3(n27482), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n34475));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_20_6 (.CI(n27482), .I0(GND_net), .I1(pwm_out_0__N_562[4]), 
            .CO(n27483));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_562[3]), 
            .I3(n27481), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n27481), .I0(GND_net), .I1(pwm_out_0__N_562[3]), 
            .CO(n27482));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_562[2]), 
            .I3(n27480), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n27480), .I0(GND_net), .I1(pwm_out_0__N_562[2]), 
            .CO(n27481));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_562[1]), 
            .I3(n27479), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 count_0__1139_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n28353), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1139_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n28352), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_11 (.CI(n28352), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n28353));
    SB_LUT4 count_0__1139_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n28351), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_10 (.CI(n28351), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n28352));
    SB_CARRY pwm_out_0__I_20_3 (.CI(n27479), .I0(GND_net), .I1(pwm_out_0__N_562[1]), 
            .CO(n27480));
    SB_LUT4 count_0__1139_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n28350), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_9 (.CI(n28350), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n28351));
    SB_LUT4 count_0__1139_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n28349), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_562[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY count_0__1139_add_4_8 (.CI(n28349), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n28350));
    SB_LUT4 count_0__1139_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n28348), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_7 (.CI(n28348), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n28349));
    SB_LUT4 count_0__1139_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n28347), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_6 (.CI(n28347), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n28348));
    SB_LUT4 count_0__1139_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n28346), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_5 (.CI(n28346), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n28347));
    SB_LUT4 count_0__1139_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n28345), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18555_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1035), .I3(GND_net), .O(n23054));
    defparam i18555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30809_2_lut (.I0(\count[0] [8]), .I1(\count[0] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n37057));
    defparam i30809_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(\count[0] [4]), .I1(\count[0] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n12));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY count_0__1139_add_4_4 (.CI(n28345), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n28346));
    SB_LUT4 i7_4_lut (.I0(n37057), .I1(\count[0] [3]), .I2(\count[0] [10]), 
            .I3(pause_counter_0), .O(n18));
    defparam i7_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i8_4_lut (.I0(\count[0] [9]), .I1(\count[0] [0]), .I2(\count[0] [1]), 
            .I3(\count[0] [2]), .O(n19));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut (.I0(n19), .I1(\count[0] [7]), .I2(n18), .I3(n12), 
            .O(n1035));
    defparam i10_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 count_0__1139_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n28344), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_562[0]), 
            .CO(n27479));
    SB_CARRY count_0__1139_add_4_3 (.CI(n28344), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n28345));
    SB_LUT4 count_0__1139_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1139_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1139_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n28344));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n27488), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27489));
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n17932));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35380_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_557), .I2(GND_net), 
            .I3(GND_net), .O(n34475));
    defparam i35380_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_639[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_639[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_639[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_639[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(half_duty_new[5]), .C(CLK_c), .D(half_duty_new_9__N_639[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_639[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_639[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i8_4_lut_adj_845 (.I0(n4), .I1(n40977), .I2(n40979), .I3(pwm_out_0__N_561), 
            .O(n20));
    defparam i8_4_lut_adj_845.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\count[0] [10]), .I1(n5), .I2(GND_net), 
            .I3(GND_net), .O(n13));
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h2222;
    SB_LUT4 i10_4_lut_adj_847 (.I0(n13), .I1(n20), .I2(n8), .I3(n40981), 
            .O(n22));
    defparam i10_4_lut_adj_847.LUT_INIT = 16'h0008;
    SB_LUT4 i30922_4_lut (.I0(n2), .I1(n3), .I2(n10), .I3(n1), .O(n37176));
    defparam i30922_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n37176), .I1(pause_counter_0), .I2(pwm_out_0__N_557), 
            .I3(n22), .O(n17544));
    defparam i1_4_lut.LUT_INIT = 16'h1303;
    SB_LUT4 i3_4_lut (.I0(\half_duty[0][4] ), .I1(\half_duty[0][1] ), .I2(\count[0] [4]), 
            .I3(\count[0] [1]), .O(n14));   // vhdl/pwm.vhd(80[8:31])
    defparam i3_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_848 (.I0(\count[0] [0]), .I1(n14), .I2(\count[0] [10]), 
            .I3(\half_duty[0][0] ), .O(n18_adj_3560));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_4_lut_adj_848.LUT_INIT = 16'hfdfe;
    SB_LUT4 i5_4_lut (.I0(\half_duty[0][3] ), .I1(\half_duty[0][2] ), .I2(\count[0] [3]), 
            .I3(\count[0] [2]), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i6_4_lut (.I0(\count[0] [6]), .I1(\count[0] [9]), .I2(\half_duty[0][6] ), 
            .I3(\count[0] [8]), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i4_4_lut (.I0(\half_duty[0][7] ), .I1(\count[0] [5]), .I2(\count[0] [7]), 
            .I3(\half_duty[0] [5]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10_4_lut_adj_849 (.I0(n15), .I1(n17), .I2(n16), .I3(n18_adj_3560), 
            .O(pwm_out_0__N_557));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_849.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2015_24_lut (.I0(GND_net), .I1(n5649[22]), .I2(pwm_setpoint[22]), 
            .I3(n27756), .O(half_duty_new_9__N_639[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2015_23_lut (.I0(GND_net), .I1(n5649[21]), .I2(pwm_setpoint[21]), 
            .I3(n27755), .O(half_duty_new_9__N_639[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_23 (.CI(n27755), .I0(n5649[21]), .I1(pwm_setpoint[21]), 
            .CO(n27756));
    SB_LUT4 add_2015_22_lut (.I0(GND_net), .I1(n5649[20]), .I2(pwm_setpoint[20]), 
            .I3(n27754), .O(half_duty_new_9__N_639[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_22 (.CI(n27754), .I0(n5649[20]), .I1(pwm_setpoint[20]), 
            .CO(n27755));
    SB_LUT4 add_2015_21_lut (.I0(GND_net), .I1(n5649[19]), .I2(pwm_setpoint[19]), 
            .I3(n27753), .O(half_duty_new_9__N_639[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_21 (.CI(n27753), .I0(n5649[19]), .I1(pwm_setpoint[19]), 
            .CO(n27754));
    SB_LUT4 add_2015_20_lut (.I0(GND_net), .I1(n5649[18]), .I2(pwm_setpoint[18]), 
            .I3(n27752), .O(half_duty_new_9__N_639[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_20 (.CI(n27752), .I0(n5649[18]), .I1(pwm_setpoint[18]), 
            .CO(n27753));
    SB_LUT4 add_2015_19_lut (.I0(GND_net), .I1(n5649[17]), .I2(pwm_setpoint[17]), 
            .I3(n27751), .O(half_duty_new_9__N_639[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_19 (.CI(n27751), .I0(n5649[17]), .I1(pwm_setpoint[17]), 
            .CO(n27752));
    SB_LUT4 add_2015_18_lut (.I0(GND_net), .I1(n5649[16]), .I2(pwm_setpoint[16]), 
            .I3(n27750), .O(half_duty_new_9__N_639[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_18 (.CI(n27750), .I0(n5649[16]), .I1(pwm_setpoint[16]), 
            .CO(n27751));
    SB_LUT4 add_2015_17_lut (.I0(GND_net), .I1(n5649[15]), .I2(pwm_setpoint[15]), 
            .I3(n27749), .O(half_duty_new_9__N_639[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2015_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2015_17 (.CI(n27749), .I0(n5649[15]), .I1(pwm_setpoint[15]), 
            .CO(n27750));
    SB_CARRY add_2015_16 (.CI(n27748), .I0(n5649[14]), .I1(pwm_setpoint[14]), 
            .CO(n27749));
    SB_CARRY add_2015_15 (.CI(n27747), .I0(n5649[13]), .I1(pwm_setpoint[13]), 
            .CO(n27748));
    SB_CARRY add_2015_14 (.CI(n27746), .I0(n5649[12]), .I1(pwm_setpoint[12]), 
            .CO(n27747));
    SB_CARRY add_2015_13 (.CI(n27745), .I0(n5649[11]), .I1(pwm_setpoint[11]), 
            .CO(n27746));
    SB_CARRY add_2015_12 (.CI(n27744), .I0(n5649[10]), .I1(pwm_setpoint[10]), 
            .CO(n27745));
    SB_CARRY add_2015_11 (.CI(n27743), .I0(n5649[9]), .I1(pwm_setpoint[9]), 
            .CO(n27744));
    SB_CARRY add_2015_10 (.CI(n27742), .I0(n5649[8]), .I1(pwm_setpoint[8]), 
            .CO(n27743));
    SB_CARRY add_2015_9 (.CI(n27741), .I0(n5649[7]), .I1(pwm_setpoint[7]), 
            .CO(n27742));
    SB_CARRY add_2015_8 (.CI(n27740), .I0(n5649[6]), .I1(pwm_setpoint[6]), 
            .CO(n27741));
    SB_CARRY add_2015_7 (.CI(n27739), .I0(n5649[5]), .I1(pwm_setpoint[5]), 
            .CO(n27740));
    SB_CARRY add_2015_6 (.CI(n27738), .I0(n5649[4]), .I1(pwm_setpoint[4]), 
            .CO(n27739));
    SB_CARRY add_2015_5 (.CI(n27737), .I0(n5649[3]), .I1(pwm_setpoint[3]), 
            .CO(n27738));
    SB_CARRY add_2015_4 (.CI(n27736), .I0(n5649[2]), .I1(pwm_setpoint[2]), 
            .CO(n27737));
    SB_CARRY add_2015_3 (.CI(n27735), .I0(n5649[1]), .I1(pwm_setpoint[1]), 
            .CO(n27736));
    SB_CARRY add_2015_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n27735));
    SB_LUT4 add_2023_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n27734), .O(n5649[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2023_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n27733), .O(n5649[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_22 (.CI(n27733), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n27734));
    SB_LUT4 add_2023_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n27732), .O(n5649[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_21 (.CI(n27732), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n27733));
    SB_LUT4 add_2023_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n27731), .O(n5649[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_20 (.CI(n27731), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n27732));
    SB_LUT4 add_2023_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n27730), .O(n5649[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_19 (.CI(n27730), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n27731));
    SB_LUT4 add_2023_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n27729), .O(n5649[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_18 (.CI(n27729), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n27730));
    SB_LUT4 add_2023_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n27728), .O(n5649[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_17 (.CI(n27728), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n27729));
    SB_LUT4 add_2023_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n27727), .O(n5649[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_16 (.CI(n27727), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n27728));
    SB_LUT4 add_2023_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n27726), .O(n5649[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_15 (.CI(n27726), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n27727));
    SB_LUT4 add_2023_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n27725), .O(n5649[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_14 (.CI(n27725), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n27726));
    SB_LUT4 add_2023_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n27724), .O(n5649[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_13 (.CI(n27724), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n27725));
    SB_LUT4 add_2023_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n27723), .O(n5649[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_12 (.CI(n27723), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n27724));
    SB_LUT4 add_2023_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n27722), .O(n5649[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_11 (.CI(n27722), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n27723));
    SB_LUT4 add_2023_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n27721), .O(n5649[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_10 (.CI(n27721), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n27722));
    SB_LUT4 add_2023_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n27720), .O(n5649[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_9 (.CI(n27720), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n27721));
    SB_LUT4 add_2023_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n27719), .O(n5649[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_8 (.CI(n27719), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n27720));
    SB_LUT4 add_2023_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n27718), .O(n5649[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_7 (.CI(n27718), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n27719));
    SB_LUT4 add_2023_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n27717), .O(n5649[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_6 (.CI(n27717), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n27718));
    SB_LUT4 add_2023_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n27716), .O(n5649[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_5 (.CI(n27716), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n27717));
    SB_LUT4 add_2023_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n27715), .O(n5649[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_4 (.CI(n27715), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n27716));
    SB_LUT4 add_2023_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n27714), .O(n5649[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_3 (.CI(n27714), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n27715));
    SB_LUT4 add_2023_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5649[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2023_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2023_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n27714));
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0] [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18563_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_out_0__N_562[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i18563_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_562[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_587));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[6] , motor_state, \Kp[1] , \Kp[0] , 
            setpoint, \Kp[2] , \Kp[7] , duty, VCC_net, PWMLimit, 
            clk32MHz, \Kp[3] , \Kp[4] , \Kp[5] , n41708) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input \Kp[6] ;
    input [23:0]motor_state;
    input \Kp[1] ;
    input \Kp[0] ;
    input [23:0]setpoint;
    input \Kp[2] ;
    input \Kp[7] ;
    output [23:0]duty;
    input VCC_net;
    input [23:0]PWMLimit;
    input clk32MHz;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    output n41708;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [14:0]n8715;
    wire [13:0]n8732;
    
    wire n29104, n29103;
    wire [23:0]n103;
    wire [23:0]n1;
    
    wire n27593, n27594, n27592, n29102, n29101, n27591, n29100, 
        n29099;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n460, n29098, n29097, n536, n29096;
    wire [23:0]\PID_CONTROLLER.err_23__N_3354 ;
    wire [23:0]n1_adj_3559;
    
    wire n27635, n463, n29095, n390, n29094, n317, n29093, n244, 
        n29092, n27634, n27590, n171, n29091, n29, n98, n83, 
        n14, n156, n533;
    wire [15:0]n8697;
    
    wire n29090, n29089, n39701, n6, n29088, n29087, n39, n41, 
        n45, n29086, n29085, n37, n29084;
    wire [23:0]duty_23__N_3330;
    
    wire n29_adj_3461, n31, n29083, n29082, n43, n23_adj_3462, n25_adj_3463, 
        n35, n33, n29081, n11, n229, n15, n27, n29080, n9, 
        n17, n19_adj_3464, n21_adj_3465, n387, n29079, n314, n29078, 
        n13, n39202, n39111, n241, n29077, n27633, n168, n29076, 
        n26, n95, n27632;
    wire [16:0]n8678;
    
    wire n29075, n29074, n27631, n27630, n27629, n27628, n12, 
        n30, n39357, n39890, n29073, n27627, n39862, n40700, n27626, 
        n40252, n29072, n40844, n27625, n6_adj_3470, n40692, n40693, 
        n29071, n16, n24_adj_3471, n39711, n29070, n27624, n29069, 
        n29068, n29067, n8_adj_3473, n39705, n40324, n40530, n4_adj_3474, 
        n40541, n29066, n530, n29065, n40542, n39746, n457, n29064, 
        n384, n29063, n311, n29062, n238, n29061, n165, n29060, 
        n23_adj_3475, n92;
    wire [17:0]n8658;
    
    wire n29059, n29058, n10_adj_3476, n39741, n40820, n29057, n39911, 
        n29056;
    wire [21:0]n8568;
    wire [20:0]n8592;
    
    wire n28595, n28594, n28593, n29055, n28592, n29054, n28591, 
        n29053, n40931, n29052, n28590, n302, n375, n448, n40932, 
        n40906, n29051, n28589, n521, n28588, n28587, n29050, 
        n39717, n28586, n29049, n527, n29048, n28585, n454, n29047, 
        n40730, n28584, n39917, n381, n29046, n28583, n40852, 
        n27623, n28582, duty_23__N_3402, n308, n29045, n41_adj_3478, 
        n39_adj_3479, n45_adj_3480, n235, n29044, n43_adj_3481, n37_adj_3482, 
        n28581, n29_adj_3483, n27622, n515, n28580, n31_adj_3485, 
        n23_adj_3486, n25_adj_3487, n162, n29043, n442, n28579, 
        n11_adj_3488, n27_adj_3489, n35_adj_3490, n369, n28578, n296, 
        n28577, n223, n28576, n20, n89, n150, n28575;
    wire [18:0]n8637;
    
    wire n29042, n29041, n8_adj_3491, n77, n29040, n29039, n27621, 
        n29038, n29037, n29036, n29035, n29034, n29033, n29032, 
        n13_adj_3493, n29031, n15_adj_3494, n524, n29030, n451, 
        n29029, n27620, n378, n29028, n33_adj_3496, n305, n29027, 
        n232, n29026, n86, n17_adj_3497, n9_adj_3498, n17_adj_3499, 
        n19_adj_3500, n159, n29025, n21_adj_3501;
    wire [19:0]n8615;
    
    wire n29024, n29023, n39675, n39661, n27619, n12_adj_3502, n10_adj_3503, 
        n30_adj_3504, n40202, n40196, n40794, n40425, n29022, n40867, 
        n16_adj_3505, n29021, n29020, n29019, n29018, n29017, n29016, 
        n29015, n40537, n29014, n40538, n29013, n29012, n29011, 
        n29010, n29009, n29008, n29007, n29006, n27618, n29005, 
        n29004, n29003, n27617, n29002, n29001, n29000, n8_adj_3507, 
        n24_adj_3508, n39621, n39593, n40326, n39919, n4_adj_3509, 
        n40533, n40534, n39649, n39641, n40822, n39921, n40933, 
        n40934, n40904, n39623, n40732, n28999, n28998, n27616, 
        n28997, n28996, n28995, n39927, n28994, n28993, n27615, 
        n27614, n28992, n518, n28991, n445, n28990, n372, n28989, 
        n299, n28988, n226, n28987, n153, n28986, n11_adj_3513, 
        n80, n39021, n28985;
    wire [47:0]n28;
    
    wire n28984, n28983, n28982, n27613, n28981, n28980, n40854, 
        n28979, n102, n28978, n28977, n28976;
    wire [23:0]duty_23__N_3378;
    
    wire n28975, n28974, n28973, n28972, n28971, n28970;
    wire [5:0]n8832;
    
    wire n35928, n490, n29185;
    wire [4:0]n8840;
    
    wire n417, n29184, n512, n28969, n344, n29183, n439, n28968, 
        n366, n28967, n271, n29182, n198, n29181, n293, n28966, 
        n220, n28965, n27612, n147, n28964, n56_adj_3517, n125_adj_3518, 
        n5_adj_3519, n74_adj_3520;
    wire [6:0]n8823;
    
    wire n560, n29180, n487, n29179, n414, n29178, n341, n29177, 
        n268, n29176, n195, n29175, n53_adj_3521, n122_adj_3522;
    wire [7:0]n8813;
    
    wire n29174, n557, n29173, n484, n29172, n411, n29171, n338, 
        n29170, n27611, n265, n29169, n192, n29168, n50, n119_adj_3524;
    wire [8:0]n8802;
    
    wire n29167, n29166, n554, n29165, n481, n29164, n27610, n408, 
        n29163, n335, n29162, n262, n29161, n27609, n189, n29160, 
        n47, n116_adj_3527;
    wire [9:0]n8790;
    
    wire n29159, n29158, n27608, n29157, n551, n29156, n478, n29155, 
        n405, n29154, n27607, n332, n29153, n27606, n259, n29152, 
        n186, n29151, n44, n113_adj_3531;
    wire [10:0]n8777;
    
    wire n29150, n29149, n29148, n29147, n548, n29146, n27605, 
        n101, n475, n29145, n32, n402, n29144, n329, n29143, 
        n256, n29142, n174, n247, n183, n29141, n41_adj_3535, 
        n110_adj_3536;
    wire [11:0]n8763;
    
    wire n29140, n29139, n320, n29138, n393, n27604, n29137, n466, 
        n29136, n545, n29135, n539, n472, n29134, n27603, n399, 
        n29133, n27602, n27601, n27600, n104_adj_3543, n35_adj_3544, 
        n177, n326, n29132, n253, n29131, n180, n29130, n250, 
        n38, n107_adj_3545, n323, n396;
    wire [12:0]n8748;
    
    wire n29129, n29128, n27599, n29127, n29126, n27598, n29125, 
        n29124, n542, n29123, n469, n29122, n27597, n29121, n29120, 
        n29119, n29118, n29117, n29116, n29115, n29114, n29113, 
        n29112, n29111, n29110, n27596, n29109, n29108, n29107, 
        n27595, n29106, n29105, n6_adj_3549;
    wire [3:0]n8847;
    
    wire n4_adj_3550;
    wire [2:0]n8853;
    
    wire n207;
    wire [1:0]n8858;
    
    wire n27395, n6_adj_3551, n27420, n14_adj_3552, n8_adj_3553, n12_adj_3554, 
        n11_adj_3555, n15_adj_3556, n17_adj_3557, n27361, n4_adj_3558, 
        n27318;
    
    SB_LUT4 add_4604_16_lut (.I0(GND_net), .I1(n8732[13]), .I2(GND_net), 
            .I3(n29104), .O(n8715[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_15_lut (.I0(GND_net), .I1(n8732[12]), .I2(GND_net), 
            .I3(n29103), .O(n8715[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n27593), .O(n103[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_15 (.CI(n29103), .I0(n8732[12]), .I1(GND_net), .CO(n29104));
    SB_CARRY unary_minus_8_add_3_6 (.CI(n27593), .I0(GND_net), .I1(n1[4]), 
            .CO(n27594));
    SB_LUT4 unary_minus_8_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n27592), .O(n103[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_14_lut (.I0(GND_net), .I1(n8732[11]), .I2(GND_net), 
            .I3(n29102), .O(n8715[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_14 (.CI(n29102), .I0(n8732[11]), .I1(GND_net), .CO(n29103));
    SB_LUT4 add_4604_13_lut (.I0(GND_net), .I1(n8732[10]), .I2(GND_net), 
            .I3(n29101), .O(n8715[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_5 (.CI(n27592), .I0(GND_net), .I1(n1[3]), 
            .CO(n27593));
    SB_CARRY add_4604_13 (.CI(n29101), .I0(n8732[10]), .I1(GND_net), .CO(n29102));
    SB_LUT4 unary_minus_8_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n27591), .O(n103[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_12_lut (.I0(GND_net), .I1(n8732[9]), .I2(GND_net), 
            .I3(n29100), .O(n8715[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_12 (.CI(n29100), .I0(n8732[9]), .I1(GND_net), .CO(n29101));
    SB_LUT4 add_4604_11_lut (.I0(GND_net), .I1(n8732[8]), .I2(GND_net), 
            .I3(n29099), .O(n8715[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4604_11 (.CI(n29099), .I0(n8732[8]), .I1(GND_net), .CO(n29100));
    SB_LUT4 add_4604_10_lut (.I0(GND_net), .I1(n8732[7]), .I2(GND_net), 
            .I3(n29098), .O(n8715[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_10 (.CI(n29098), .I0(n8732[7]), .I1(GND_net), .CO(n29099));
    SB_LUT4 add_4604_9_lut (.I0(GND_net), .I1(n8732[6]), .I2(GND_net), 
            .I3(n29097), .O(n8715[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_9 (.CI(n29097), .I0(n8732[6]), .I1(GND_net), .CO(n29098));
    SB_LUT4 add_4604_8_lut (.I0(GND_net), .I1(n8732[5]), .I2(n536), .I3(n29096), 
            .O(n8715[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_3559[23]), .I3(n27635), .O(\PID_CONTROLLER.err_23__N_3354 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_8 (.CI(n29096), .I0(n8732[5]), .I1(n536), .CO(n29097));
    SB_LUT4 add_4604_7_lut (.I0(GND_net), .I1(n8732[4]), .I2(n463), .I3(n29095), 
            .O(n8715[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_7 (.CI(n29095), .I0(n8732[4]), .I1(n463), .CO(n29096));
    SB_LUT4 add_4604_6_lut (.I0(GND_net), .I1(n8732[3]), .I2(n390), .I3(n29094), 
            .O(n8715[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_6 (.CI(n29094), .I0(n8732[3]), .I1(n390), .CO(n29095));
    SB_LUT4 add_4604_5_lut (.I0(GND_net), .I1(n8732[2]), .I2(n317), .I3(n29093), 
            .O(n8715[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_5 (.CI(n29093), .I0(n8732[2]), .I1(n317), .CO(n29094));
    SB_LUT4 add_4604_4_lut (.I0(GND_net), .I1(n8732[1]), .I2(n244), .I3(n29092), 
            .O(n8715[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_3559[22]), .I3(n27634), .O(\PID_CONTROLLER.err_23__N_3354 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_4 (.CI(n27591), .I0(GND_net), .I1(n1[2]), 
            .CO(n27592));
    SB_CARRY add_4604_4 (.CI(n29092), .I0(n8732[1]), .I1(n244), .CO(n29093));
    SB_LUT4 unary_minus_8_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n27590), .O(n103[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_3_lut (.I0(GND_net), .I1(n8732[0]), .I2(n171), .I3(n29091), 
            .O(n8715[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_3 (.CI(n27590), .I0(GND_net), .I1(n1[1]), 
            .CO(n27591));
    SB_CARRY add_4604_3 (.CI(n29091), .I0(n8732[0]), .I1(n171), .CO(n29092));
    SB_LUT4 add_4604_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n8715[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n29091));
    SB_LUT4 mult_4_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[6]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4603_17_lut (.I0(GND_net), .I1(n8715[14]), .I2(GND_net), 
            .I3(n29090), .O(n8697[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4603_16_lut (.I0(GND_net), .I1(n8715[13]), .I2(GND_net), 
            .I3(n29089), .O(n8697[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33379_3_lut_4_lut (.I0(duty[3]), .I1(n103[3]), .I2(n103[2]), 
            .I3(duty[2]), .O(n39701));   // verilog/motorControl.v(45[19:35])
    defparam i33379_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_8_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n103[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_7_i6_3_lut_3_lut (.I0(duty[3]), .I1(n103[3]), .I2(n103[2]), 
            .I3(GND_net), .O(n6));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_4603_16 (.CI(n29089), .I0(n8715[13]), .I1(GND_net), .CO(n29090));
    SB_LUT4 add_4603_15_lut (.I0(GND_net), .I1(n8715[12]), .I2(GND_net), 
            .I3(n29088), .O(n8697[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_15 (.CI(n29088), .I0(n8715[12]), .I1(GND_net), .CO(n29089));
    SB_LUT4 add_4603_14_lut (.I0(GND_net), .I1(n8715[11]), .I2(GND_net), 
            .I3(n29087), .O(n8697[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4603_14 (.CI(n29087), .I0(n8715[11]), .I1(GND_net), .CO(n29088));
    SB_LUT4 add_4603_13_lut (.I0(GND_net), .I1(n8715[10]), .I2(GND_net), 
            .I3(n29086), .O(n8697[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_13 (.CI(n29086), .I0(n8715[10]), .I1(GND_net), .CO(n29087));
    SB_LUT4 add_4603_12_lut (.I0(GND_net), .I1(n8715[9]), .I2(GND_net), 
            .I3(n29085), .O(n8697[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4603_12 (.CI(n29085), .I0(n8715[9]), .I1(GND_net), .CO(n29086));
    SB_LUT4 add_4603_11_lut (.I0(GND_net), .I1(n8715[8]), .I2(GND_net), 
            .I3(n29084), .O(n8697[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_11 (.CI(n29084), .I0(n8715[8]), .I1(GND_net), .CO(n29085));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3330[0]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [0]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3461));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4603_10_lut (.I0(GND_net), .I1(n8715[7]), .I2(GND_net), 
            .I3(n29083), .O(n8697[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_10 (.CI(n29083), .I0(n8715[7]), .I1(GND_net), .CO(n29084));
    SB_LUT4 add_4603_9_lut (.I0(GND_net), .I1(n8715[6]), .I2(GND_net), 
            .I3(n29082), .O(n8697[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_9 (.CI(n29082), .I0(n8715[6]), .I1(GND_net), .CO(n29083));
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3462));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3463));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4603_8_lut (.I0(GND_net), .I1(n8715[5]), .I2(n533), .I3(n29081), 
            .O(n8697[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_4_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4603_8 (.CI(n29081), .I0(n8715[5]), .I1(n533), .CO(n29082));
    SB_LUT4 add_4603_7_lut (.I0(GND_net), .I1(n8715[4]), .I2(n460), .I3(n29080), 
            .O(n8697[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_7 (.CI(n29080), .I0(n8715[4]), .I1(n460), .CO(n29081));
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3464));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3465));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_8_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n27590));
    SB_LUT4 add_4603_6_lut (.I0(GND_net), .I1(n8715[3]), .I2(n387), .I3(n29079), 
            .O(n8697[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_6 (.CI(n29079), .I0(n8715[3]), .I1(n387), .CO(n29080));
    SB_CARRY state_23__I_0_add_2_24 (.CI(n27634), .I0(motor_state[22]), 
            .I1(n1_adj_3559[22]), .CO(n27635));
    SB_LUT4 add_4603_5_lut (.I0(GND_net), .I1(n8715[2]), .I2(n314), .I3(n29078), 
            .O(n8697[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_5 (.CI(n29078), .I0(n8715[2]), .I1(n314), .CO(n29079));
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32882_4_lut (.I0(n21_adj_3465), .I1(n19_adj_3464), .I2(n17), 
            .I3(n9), .O(n39202));
    defparam i32882_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32791_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n39111));
    defparam i32791_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4603_4_lut (.I0(GND_net), .I1(n8715[1]), .I2(n241), .I3(n29077), 
            .O(n8697[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_3559[21]), .I3(n27633), .O(\PID_CONTROLLER.err_23__N_3354 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_4 (.CI(n29077), .I0(n8715[1]), .I1(n241), .CO(n29078));
    SB_LUT4 add_4603_3_lut (.I0(GND_net), .I1(n8715[0]), .I2(n168), .I3(n29076), 
            .O(n8697[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_3 (.CI(n29076), .I0(n8715[0]), .I1(n168), .CO(n29077));
    SB_CARRY state_23__I_0_add_2_23 (.CI(n27633), .I0(motor_state[21]), 
            .I1(n1_adj_3559[21]), .CO(n27634));
    SB_LUT4 add_4603_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n8697[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n29076));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_3559[20]), .I3(n27632), .O(\PID_CONTROLLER.err_23__N_3354 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_18_lut (.I0(GND_net), .I1(n8697[15]), .I2(GND_net), 
            .I3(n29075), .O(n8678[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_17_lut (.I0(GND_net), .I1(n8697[14]), .I2(GND_net), 
            .I3(n29074), .O(n8678[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_17 (.CI(n29074), .I0(n8697[14]), .I1(GND_net), .CO(n29075));
    SB_CARRY state_23__I_0_add_2_22 (.CI(n27632), .I0(motor_state[20]), 
            .I1(n1_adj_3559[20]), .CO(n27633));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_3559[19]), .I3(n27631), .O(\PID_CONTROLLER.err_23__N_3354 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n27631), .I0(motor_state[19]), 
            .I1(n1_adj_3559[19]), .CO(n27632));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_3559[18]), .I3(n27630), .O(\PID_CONTROLLER.err_23__N_3354 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n27630), .I0(motor_state[18]), 
            .I1(n1_adj_3559[18]), .CO(n27631));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_3559[17]), .I3(n27629), .O(\PID_CONTROLLER.err_23__N_3354 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n27629), .I0(motor_state[17]), 
            .I1(n1_adj_3559[17]), .CO(n27630));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_3559[16]), .I3(n27628), .O(\PID_CONTROLLER.err_23__N_3354 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(duty[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n27628), .I0(motor_state[16]), 
            .I1(n1_adj_3559[16]), .CO(n27629));
    SB_LUT4 i33568_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n39357), 
            .O(n39890));
    defparam i33568_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_4602_16_lut (.I0(GND_net), .I1(n8697[13]), .I2(GND_net), 
            .I3(n29073), .O(n8678[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_16 (.CI(n29073), .I0(n8697[13]), .I1(GND_net), .CO(n29074));
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_3559[15]), .I3(n27627), .O(\PID_CONTROLLER.err_23__N_3354 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n27627), .I0(motor_state[15]), 
            .I1(n1_adj_3559[15]), .CO(n27628));
    SB_LUT4 unary_minus_8_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33540_4_lut (.I0(n19_adj_3464), .I1(n17), .I2(n15), .I3(n39890), 
            .O(n39862));
    defparam i33540_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34378_4_lut (.I0(n25_adj_3463), .I1(n23_adj_3462), .I2(n21_adj_3465), 
            .I3(n39862), .O(n40700));
    defparam i34378_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_3559[14]), .I3(n27626), .O(\PID_CONTROLLER.err_23__N_3354 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33930_4_lut (.I0(n31), .I1(n29_adj_3461), .I2(n27), .I3(n40700), 
            .O(n40252));
    defparam i33930_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_4602_15_lut (.I0(GND_net), .I1(n8697[12]), .I2(GND_net), 
            .I3(n29072), .O(n8678[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n27626), .I0(motor_state[14]), 
            .I1(n1_adj_3559[14]), .CO(n27627));
    SB_LUT4 i34522_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n40252), 
            .O(n40844));
    defparam i34522_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_4602_15 (.CI(n29072), .I0(n8697[12]), .I1(GND_net), .CO(n29073));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_3559[13]), .I3(n27625), .O(\PID_CONTROLLER.err_23__N_3354 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34370_3_lut (.I0(n6_adj_3470), .I1(duty[10]), .I2(n21_adj_3465), 
            .I3(GND_net), .O(n40692));   // verilog/motorControl.v(43[10:25])
    defparam i34370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34371_3_lut (.I0(n40692), .I1(duty[11]), .I2(n23_adj_3462), 
            .I3(GND_net), .O(n40693));   // verilog/motorControl.v(43[10:25])
    defparam i34371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4602_14_lut (.I0(GND_net), .I1(n8697[11]), .I2(GND_net), 
            .I3(n29071), .O(n8678[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(duty[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_3471));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n27625), .I0(motor_state[13]), 
            .I1(n1_adj_3559[13]), .CO(n27626));
    SB_LUT4 i33389_4_lut (.I0(n43), .I1(n25_adj_3463), .I2(n23_adj_3462), 
            .I3(n39202), .O(n39711));
    defparam i33389_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4602_14 (.CI(n29071), .I0(n8697[11]), .I1(GND_net), .CO(n29072));
    SB_LUT4 add_4602_13_lut (.I0(GND_net), .I1(n8697[10]), .I2(GND_net), 
            .I3(n29070), .O(n8678[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_13 (.CI(n29070), .I0(n8697[10]), .I1(GND_net), .CO(n29071));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_3559[12]), .I3(n27624), .O(\PID_CONTROLLER.err_23__N_3354 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_12_lut (.I0(GND_net), .I1(n8697[9]), .I2(GND_net), 
            .I3(n29069), .O(n8678[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_12 (.CI(n29069), .I0(n8697[9]), .I1(GND_net), .CO(n29070));
    SB_LUT4 add_4602_11_lut (.I0(GND_net), .I1(n8697[8]), .I2(GND_net), 
            .I3(n29068), .O(n8678[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_11 (.CI(n29068), .I0(n8697[8]), .I1(GND_net), .CO(n29069));
    SB_LUT4 add_4602_10_lut (.I0(GND_net), .I1(n8697[7]), .I2(GND_net), 
            .I3(n29067), .O(n8678[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34002_4_lut (.I0(n24_adj_3471), .I1(n8_adj_3473), .I2(n45), 
            .I3(n39705), .O(n40324));   // verilog/motorControl.v(43[10:25])
    defparam i34002_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34208_3_lut (.I0(n40693), .I1(duty[12]), .I2(n25_adj_3463), 
            .I3(GND_net), .O(n40530));   // verilog/motorControl.v(43[10:25])
    defparam i34208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34219_3_lut (.I0(n4_adj_3474), .I1(duty[13]), .I2(n27), .I3(GND_net), 
            .O(n40541));   // verilog/motorControl.v(43[10:25])
    defparam i34219_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4602_10 (.CI(n29067), .I0(n8697[7]), .I1(GND_net), .CO(n29068));
    SB_LUT4 add_4602_9_lut (.I0(GND_net), .I1(n8697[6]), .I2(GND_net), 
            .I3(n29066), .O(n8678[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_9 (.CI(n29066), .I0(n8697[6]), .I1(GND_net), .CO(n29067));
    SB_LUT4 add_4602_8_lut (.I0(GND_net), .I1(n8697[5]), .I2(n530), .I3(n29065), 
            .O(n8678[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_8 (.CI(n29065), .I0(n8697[5]), .I1(n530), .CO(n29066));
    SB_LUT4 i34220_3_lut (.I0(n40541), .I1(duty[14]), .I2(n29_adj_3461), 
            .I3(GND_net), .O(n40542));   // verilog/motorControl.v(43[10:25])
    defparam i34220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33424_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_3461), .I3(n39111), 
            .O(n39746));
    defparam i33424_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4602_7_lut (.I0(GND_net), .I1(n8697[4]), .I2(n457), .I3(n29064), 
            .O(n8678[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_7 (.CI(n29064), .I0(n8697[4]), .I1(n457), .CO(n29065));
    SB_LUT4 add_4602_6_lut (.I0(GND_net), .I1(n8697[3]), .I2(n384), .I3(n29063), 
            .O(n8678[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_6 (.CI(n29063), .I0(n8697[3]), .I1(n384), .CO(n29064));
    SB_LUT4 add_4602_5_lut (.I0(GND_net), .I1(n8697[2]), .I2(n311), .I3(n29062), 
            .O(n8678[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_5 (.CI(n29062), .I0(n8697[2]), .I1(n311), .CO(n29063));
    SB_LUT4 add_4602_4_lut (.I0(GND_net), .I1(n8697[1]), .I2(n238), .I3(n29061), 
            .O(n8678[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_4 (.CI(n29061), .I0(n8697[1]), .I1(n238), .CO(n29062));
    SB_LUT4 add_4602_3_lut (.I0(GND_net), .I1(n8697[0]), .I2(n165), .I3(n29060), 
            .O(n8678[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n27624), .I0(motor_state[12]), 
            .I1(n1_adj_3559[12]), .CO(n27625));
    SB_CARRY add_4602_3 (.CI(n29060), .I0(n8697[0]), .I1(n165), .CO(n29061));
    SB_LUT4 add_4602_2_lut (.I0(GND_net), .I1(n23_adj_3475), .I2(n92), 
            .I3(GND_net), .O(n8678[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_2 (.CI(GND_net), .I0(n23_adj_3475), .I1(n92), .CO(n29060));
    SB_LUT4 add_4601_19_lut (.I0(GND_net), .I1(n8678[16]), .I2(GND_net), 
            .I3(n29059), .O(n8658[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4601_18_lut (.I0(GND_net), .I1(n8678[15]), .I2(GND_net), 
            .I3(n29058), .O(n8658[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34498_4_lut (.I0(n30), .I1(n10_adj_3476), .I2(n35), .I3(n39741), 
            .O(n40820));   // verilog/motorControl.v(43[10:25])
    defparam i34498_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4601_18 (.CI(n29058), .I0(n8678[15]), .I1(GND_net), .CO(n29059));
    SB_LUT4 add_4601_17_lut (.I0(GND_net), .I1(n8678[14]), .I2(GND_net), 
            .I3(n29057), .O(n8658[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33589_3_lut (.I0(n40542), .I1(duty[15]), .I2(n31), .I3(GND_net), 
            .O(n39911));   // verilog/motorControl.v(43[10:25])
    defparam i33589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4601_17 (.CI(n29057), .I0(n8678[14]), .I1(GND_net), .CO(n29058));
    SB_LUT4 add_4601_16_lut (.I0(GND_net), .I1(n8678[13]), .I2(GND_net), 
            .I3(n29056), .O(n8658[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_16 (.CI(n29056), .I0(n8678[13]), .I1(GND_net), .CO(n29057));
    SB_LUT4 add_4597_23_lut (.I0(GND_net), .I1(n8592[20]), .I2(GND_net), 
            .I3(n28595), .O(n8568[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4597_22_lut (.I0(GND_net), .I1(n8592[19]), .I2(GND_net), 
            .I3(n28594), .O(n8568[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_22 (.CI(n28594), .I0(n8592[19]), .I1(GND_net), .CO(n28595));
    SB_LUT4 add_4597_21_lut (.I0(GND_net), .I1(n8592[18]), .I2(GND_net), 
            .I3(n28593), .O(n8568[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4601_15_lut (.I0(GND_net), .I1(n8678[12]), .I2(GND_net), 
            .I3(n29055), .O(n8658[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_15 (.CI(n29055), .I0(n8678[12]), .I1(GND_net), .CO(n29056));
    SB_CARRY add_4597_21 (.CI(n28593), .I0(n8592[18]), .I1(GND_net), .CO(n28594));
    SB_LUT4 add_4597_20_lut (.I0(GND_net), .I1(n8592[17]), .I2(GND_net), 
            .I3(n28592), .O(n8568[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_20 (.CI(n28592), .I0(n8592[17]), .I1(GND_net), .CO(n28593));
    SB_LUT4 add_4601_14_lut (.I0(GND_net), .I1(n8678[11]), .I2(GND_net), 
            .I3(n29054), .O(n8658[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4597_19_lut (.I0(GND_net), .I1(n8592[16]), .I2(GND_net), 
            .I3(n28591), .O(n8568[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_14 (.CI(n29054), .I0(n8678[11]), .I1(GND_net), .CO(n29055));
    SB_LUT4 add_4601_13_lut (.I0(GND_net), .I1(n8678[10]), .I2(GND_net), 
            .I3(n29053), .O(n8658[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34609_4_lut (.I0(n39911), .I1(n40820), .I2(n35), .I3(n39746), 
            .O(n40931));   // verilog/motorControl.v(43[10:25])
    defparam i34609_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4601_13 (.CI(n29053), .I0(n8678[10]), .I1(GND_net), .CO(n29054));
    SB_CARRY add_4597_19 (.CI(n28591), .I0(n8592[16]), .I1(GND_net), .CO(n28592));
    SB_LUT4 add_4601_12_lut (.I0(GND_net), .I1(n8678[9]), .I2(GND_net), 
            .I3(n29052), .O(n8658[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4597_18_lut (.I0(GND_net), .I1(n8592[15]), .I2(GND_net), 
            .I3(n28590), .O(n8568[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4597_18 (.CI(n28590), .I0(n8592[15]), .I1(GND_net), .CO(n28591));
    SB_LUT4 mult_4_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34610_3_lut (.I0(n40931), .I1(duty[18]), .I2(n37), .I3(GND_net), 
            .O(n40932));   // verilog/motorControl.v(43[10:25])
    defparam i34610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34584_3_lut (.I0(n40932), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n40906));   // verilog/motorControl.v(43[10:25])
    defparam i34584_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4601_12 (.CI(n29052), .I0(n8678[9]), .I1(GND_net), .CO(n29053));
    SB_LUT4 add_4601_11_lut (.I0(GND_net), .I1(n8678[8]), .I2(GND_net), 
            .I3(n29051), .O(n8658[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4597_17_lut (.I0(GND_net), .I1(n8592[14]), .I2(GND_net), 
            .I3(n28589), .O(n8568[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4597_17 (.CI(n28589), .I0(n8592[14]), .I1(GND_net), .CO(n28590));
    SB_LUT4 add_4597_16_lut (.I0(GND_net), .I1(n8592[13]), .I2(GND_net), 
            .I3(n28588), .O(n8568[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_11 (.CI(n29051), .I0(n8678[8]), .I1(GND_net), .CO(n29052));
    SB_CARRY add_4597_16 (.CI(n28588), .I0(n8592[13]), .I1(GND_net), .CO(n28589));
    SB_LUT4 add_4597_15_lut (.I0(GND_net), .I1(n8592[12]), .I2(GND_net), 
            .I3(n28587), .O(n8568[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4601_10_lut (.I0(GND_net), .I1(n8678[7]), .I2(GND_net), 
            .I3(n29050), .O(n8658[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_10 (.CI(n29050), .I0(n8678[7]), .I1(GND_net), .CO(n29051));
    SB_LUT4 i33395_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n40844), 
            .O(n39717));
    defparam i33395_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4597_15 (.CI(n28587), .I0(n8592[12]), .I1(GND_net), .CO(n28588));
    SB_LUT4 add_4597_14_lut (.I0(GND_net), .I1(n8592[11]), .I2(GND_net), 
            .I3(n28586), .O(n8568[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_14 (.CI(n28586), .I0(n8592[11]), .I1(GND_net), .CO(n28587));
    SB_LUT4 add_4601_9_lut (.I0(GND_net), .I1(n8678[6]), .I2(GND_net), 
            .I3(n29049), .O(n8658[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_9 (.CI(n29049), .I0(n8678[6]), .I1(GND_net), .CO(n29050));
    SB_LUT4 add_4601_8_lut (.I0(GND_net), .I1(n8678[5]), .I2(n527), .I3(n29048), 
            .O(n8658[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_8 (.CI(n29048), .I0(n8678[5]), .I1(n527), .CO(n29049));
    SB_LUT4 add_4597_13_lut (.I0(GND_net), .I1(n8592[10]), .I2(GND_net), 
            .I3(n28585), .O(n8568[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4601_7_lut (.I0(GND_net), .I1(n8678[4]), .I2(n454), .I3(n29047), 
            .O(n8658[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34408_4_lut (.I0(n40530), .I1(n40324), .I2(n45), .I3(n39711), 
            .O(n40730));   // verilog/motorControl.v(43[10:25])
    defparam i34408_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4597_13 (.CI(n28585), .I0(n8592[10]), .I1(GND_net), .CO(n28586));
    SB_LUT4 add_4597_12_lut (.I0(GND_net), .I1(n8592[9]), .I2(GND_net), 
            .I3(n28584), .O(n8568[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_7 (.CI(n29047), .I0(n8678[4]), .I1(n454), .CO(n29048));
    SB_LUT4 i33595_3_lut (.I0(n40906), .I1(duty[20]), .I2(n41), .I3(GND_net), 
            .O(n39917));   // verilog/motorControl.v(43[10:25])
    defparam i33595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4601_6_lut (.I0(GND_net), .I1(n8678[3]), .I2(n381), .I3(n29046), 
            .O(n8658[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_12 (.CI(n28584), .I0(n8592[9]), .I1(GND_net), .CO(n28585));
    SB_LUT4 add_4597_11_lut (.I0(GND_net), .I1(n8592[8]), .I2(GND_net), 
            .I3(n28583), .O(n8568[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34530_4_lut (.I0(n39917), .I1(n40730), .I2(n45), .I3(n39717), 
            .O(n40852));   // verilog/motorControl.v(43[10:25])
    defparam i34530_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_3559[11]), .I3(n27623), .O(\PID_CONTROLLER.err_23__N_3354 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_6 (.CI(n29046), .I0(n8678[3]), .I1(n381), .CO(n29047));
    SB_CARRY add_4597_11 (.CI(n28583), .I0(n8592[8]), .I1(GND_net), .CO(n28584));
    SB_LUT4 add_4597_10_lut (.I0(GND_net), .I1(n8592[7]), .I2(GND_net), 
            .I3(n28582), .O(n8568[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34531_3_lut (.I0(n40852), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3402));   // verilog/motorControl.v(43[10:25])
    defparam i34531_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4601_5_lut (.I0(GND_net), .I1(n8678[2]), .I2(n308), .I3(n29045), 
            .O(n8658[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_10 (.CI(n28582), .I0(n8592[7]), .I1(GND_net), .CO(n28583));
    SB_CARRY state_23__I_0_add_2_13 (.CI(n27623), .I0(motor_state[11]), 
            .I1(n1_adj_3559[11]), .CO(n27624));
    SB_LUT4 LessThan_7_i41_2_lut (.I0(duty[20]), .I1(n103[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3478));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i39_2_lut (.I0(duty[19]), .I1(n103[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3479));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4601_5 (.CI(n29045), .I0(n8678[2]), .I1(n308), .CO(n29046));
    SB_LUT4 LessThan_7_i45_2_lut (.I0(duty[22]), .I1(n103[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3480));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4601_4_lut (.I0(GND_net), .I1(n8678[1]), .I2(n235), .I3(n29044), 
            .O(n8658[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[7]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_7_i43_2_lut (.I0(duty[21]), .I1(n103[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3481));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4601_4 (.CI(n29044), .I0(n8678[1]), .I1(n235), .CO(n29045));
    SB_LUT4 LessThan_7_i37_2_lut (.I0(duty[18]), .I1(n103[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3482));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4597_9_lut (.I0(GND_net), .I1(n8592[6]), .I2(GND_net), 
            .I3(n28581), .O(n8568[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_7_i29_2_lut (.I0(duty[14]), .I1(n103[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3483));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_3559[10]), .I3(n27622), .O(\PID_CONTROLLER.err_23__N_3354 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_9 (.CI(n28581), .I0(n8592[6]), .I1(GND_net), .CO(n28582));
    SB_LUT4 add_4597_8_lut (.I0(GND_net), .I1(n8592[5]), .I2(n515), .I3(n28580), 
            .O(n8568[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_7_i31_2_lut (.I0(duty[15]), .I1(n103[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3485));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i23_2_lut (.I0(duty[11]), .I1(n103[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3486));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4597_8 (.CI(n28580), .I0(n8592[5]), .I1(n515), .CO(n28581));
    SB_LUT4 LessThan_7_i25_2_lut (.I0(duty[12]), .I1(n103[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3487));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4601_3_lut (.I0(GND_net), .I1(n8678[0]), .I2(n162), .I3(n29043), 
            .O(n8658[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4597_7_lut (.I0(GND_net), .I1(n8592[4]), .I2(n442), .I3(n28579), 
            .O(n8568[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_7_i11_2_lut (.I0(duty[5]), .I1(n103[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3488));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4597_7 (.CI(n28579), .I0(n8592[4]), .I1(n442), .CO(n28580));
    SB_LUT4 LessThan_7_i27_2_lut (.I0(duty[13]), .I1(n103[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3489));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i35_2_lut (.I0(duty[17]), .I1(n103[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3490));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4597_6_lut (.I0(GND_net), .I1(n8592[3]), .I2(n369), .I3(n28578), 
            .O(n8568[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n27622), .I0(motor_state[10]), 
            .I1(n1_adj_3559[10]), .CO(n27623));
    SB_CARRY add_4597_6 (.CI(n28578), .I0(n8592[3]), .I1(n369), .CO(n28579));
    SB_LUT4 add_4597_5_lut (.I0(GND_net), .I1(n8592[2]), .I2(n296), .I3(n28577), 
            .O(n8568[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_5 (.CI(n28577), .I0(n8592[2]), .I1(n296), .CO(n28578));
    SB_LUT4 add_4597_4_lut (.I0(GND_net), .I1(n8592[1]), .I2(n223), .I3(n28576), 
            .O(n8568[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_3 (.CI(n29043), .I0(n8678[0]), .I1(n162), .CO(n29044));
    SB_CARRY add_4597_4 (.CI(n28576), .I0(n8592[1]), .I1(n223), .CO(n28577));
    SB_LUT4 add_4601_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n8658[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4601_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4601_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n29043));
    SB_LUT4 add_4597_3_lut (.I0(GND_net), .I1(n8592[0]), .I2(n150), .I3(n28575), 
            .O(n8568[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4600_20_lut (.I0(GND_net), .I1(n8658[17]), .I2(GND_net), 
            .I3(n29042), .O(n8637[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_3 (.CI(n28575), .I0(n8592[0]), .I1(n150), .CO(n28576));
    SB_LUT4 add_4600_19_lut (.I0(GND_net), .I1(n8658[16]), .I2(GND_net), 
            .I3(n29041), .O(n8637[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_19 (.CI(n29041), .I0(n8658[16]), .I1(GND_net), .CO(n29042));
    SB_LUT4 add_4597_2_lut (.I0(GND_net), .I1(n8_adj_3491), .I2(n77), 
            .I3(GND_net), .O(n8568[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4597_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4597_2 (.CI(GND_net), .I0(n8_adj_3491), .I1(n77), .CO(n28575));
    SB_LUT4 add_4600_18_lut (.I0(GND_net), .I1(n8658[15]), .I2(GND_net), 
            .I3(n29040), .O(n8637[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_18 (.CI(n29040), .I0(n8658[15]), .I1(GND_net), .CO(n29041));
    SB_LUT4 add_4600_17_lut (.I0(GND_net), .I1(n8658[14]), .I2(GND_net), 
            .I3(n29039), .O(n8637[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_3559[9]), .I3(n27621), .O(\PID_CONTROLLER.err_23__N_3354 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_17 (.CI(n29039), .I0(n8658[14]), .I1(GND_net), .CO(n29040));
    SB_LUT4 add_4600_16_lut (.I0(GND_net), .I1(n8658[13]), .I2(GND_net), 
            .I3(n29038), .O(n8637[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_16 (.CI(n29038), .I0(n8658[13]), .I1(GND_net), .CO(n29039));
    SB_LUT4 add_4600_15_lut (.I0(GND_net), .I1(n8658[12]), .I2(GND_net), 
            .I3(n29037), .O(n8637[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_15 (.CI(n29037), .I0(n8658[12]), .I1(GND_net), .CO(n29038));
    SB_LUT4 add_4600_14_lut (.I0(GND_net), .I1(n8658[11]), .I2(GND_net), 
            .I3(n29036), .O(n8637[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_14 (.CI(n29036), .I0(n8658[11]), .I1(GND_net), .CO(n29037));
    SB_LUT4 add_4600_13_lut (.I0(GND_net), .I1(n8658[10]), .I2(GND_net), 
            .I3(n29035), .O(n8637[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_13 (.CI(n29035), .I0(n8658[10]), .I1(GND_net), .CO(n29036));
    SB_LUT4 add_4600_12_lut (.I0(GND_net), .I1(n8658[9]), .I2(GND_net), 
            .I3(n29034), .O(n8637[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_12 (.CI(n29034), .I0(n8658[9]), .I1(GND_net), .CO(n29035));
    SB_LUT4 add_4600_11_lut (.I0(GND_net), .I1(n8658[8]), .I2(GND_net), 
            .I3(n29033), .O(n8637[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_11 (.CI(n29033), .I0(n8658[8]), .I1(GND_net), .CO(n29034));
    SB_LUT4 add_4600_10_lut (.I0(GND_net), .I1(n8658[7]), .I2(GND_net), 
            .I3(n29032), .O(n8637[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_10 (.CI(n29032), .I0(n8658[7]), .I1(GND_net), .CO(n29033));
    SB_LUT4 LessThan_7_i13_2_lut (.I0(duty[6]), .I1(n103[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3493));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4600_9_lut (.I0(GND_net), .I1(n8658[6]), .I2(GND_net), 
            .I3(n29031), .O(n8637[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n27621), .I0(motor_state[9]), .I1(n1_adj_3559[9]), 
            .CO(n27622));
    SB_CARRY add_4600_9 (.CI(n29031), .I0(n8658[6]), .I1(GND_net), .CO(n29032));
    SB_LUT4 LessThan_7_i15_2_lut (.I0(duty[7]), .I1(n103[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3494));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4600_8_lut (.I0(GND_net), .I1(n8658[5]), .I2(n524), .I3(n29030), 
            .O(n8637[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_8 (.CI(n29030), .I0(n8658[5]), .I1(n524), .CO(n29031));
    SB_LUT4 add_4600_7_lut (.I0(GND_net), .I1(n8658[4]), .I2(n451), .I3(n29029), 
            .O(n8637[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_7 (.CI(n29029), .I0(n8658[4]), .I1(n451), .CO(n29030));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_3559[8]), .I3(n27620), .O(\PID_CONTROLLER.err_23__N_3354 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4600_6_lut (.I0(GND_net), .I1(n8658[3]), .I2(n378), .I3(n29028), 
            .O(n8637[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_6 (.CI(n29028), .I0(n8658[3]), .I1(n378), .CO(n29029));
    SB_LUT4 LessThan_7_i33_2_lut (.I0(duty[16]), .I1(n103[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3496));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4600_5_lut (.I0(GND_net), .I1(n8658[2]), .I2(n305), .I3(n29027), 
            .O(n8637[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_5 (.CI(n29027), .I0(n8658[2]), .I1(n305), .CO(n29028));
    SB_LUT4 add_4600_4_lut (.I0(GND_net), .I1(n8658[1]), .I2(n232), .I3(n29026), 
            .O(n8637[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_4 (.CI(n29026), .I0(n8658[1]), .I1(n232), .CO(n29027));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n27620), .I0(motor_state[8]), .I1(n1_adj_3559[8]), 
            .CO(n27621));
    SB_LUT4 mult_4_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3497));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_7_i9_2_lut (.I0(duty[4]), .I1(n103[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3498));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i17_2_lut (.I0(duty[8]), .I1(n103[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3499));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_7_i19_2_lut (.I0(duty[9]), .I1(n103[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3500));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4600_3_lut (.I0(GND_net), .I1(n8658[0]), .I2(n159), .I3(n29025), 
            .O(n8637[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4600_3 (.CI(n29025), .I0(n8658[0]), .I1(n159), .CO(n29026));
    SB_LUT4 add_4600_2_lut (.I0(GND_net), .I1(n17_adj_3497), .I2(n86), 
            .I3(GND_net), .O(n8637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4600_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4600_2 (.CI(GND_net), .I0(n17_adj_3497), .I1(n86), .CO(n29025));
    SB_LUT4 LessThan_7_i21_2_lut (.I0(duty[10]), .I1(n103[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3501));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4599_21_lut (.I0(GND_net), .I1(n8637[18]), .I2(GND_net), 
            .I3(n29024), .O(n8615[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4599_20_lut (.I0(GND_net), .I1(n8637[17]), .I2(GND_net), 
            .I3(n29023), .O(n8615[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33353_4_lut (.I0(n21_adj_3501), .I1(n19_adj_3500), .I2(n17_adj_3499), 
            .I3(n9_adj_3498), .O(n39675));
    defparam i33353_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_4_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33339_4_lut (.I0(n27_adj_3489), .I1(n15_adj_3494), .I2(n13_adj_3493), 
            .I3(n11_adj_3488), .O(n39661));
    defparam i33339_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_3559[7]), .I3(n27619), .O(\PID_CONTROLLER.err_23__N_3354 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_7_i12_3_lut (.I0(n103[7]), .I1(n103[16]), .I2(n33_adj_3496), 
            .I3(GND_net), .O(n12_adj_3502));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_7_i10_3_lut (.I0(n103[5]), .I1(n103[6]), .I2(n13_adj_3493), 
            .I3(GND_net), .O(n10_adj_3503));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i30_3_lut (.I0(n12_adj_3502), .I1(n103[17]), .I2(n35_adj_3490), 
            .I3(GND_net), .O(n30_adj_3504));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33880_4_lut (.I0(n13_adj_3493), .I1(n11_adj_3488), .I2(n9_adj_3498), 
            .I3(n39701), .O(n40202));
    defparam i33880_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33874_4_lut (.I0(n19_adj_3500), .I1(n17_adj_3499), .I2(n15_adj_3494), 
            .I3(n40202), .O(n40196));
    defparam i33874_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34472_4_lut (.I0(n25_adj_3487), .I1(n23_adj_3486), .I2(n21_adj_3501), 
            .I3(n40196), .O(n40794));
    defparam i34472_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34103_4_lut (.I0(n31_adj_3485), .I1(n29_adj_3483), .I2(n27_adj_3489), 
            .I3(n40794), .O(n40425));
    defparam i34103_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_4_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4599_20 (.CI(n29023), .I0(n8637[17]), .I1(GND_net), .CO(n29024));
    SB_LUT4 add_4599_19_lut (.I0(GND_net), .I1(n8637[16]), .I2(GND_net), 
            .I3(n29022), .O(n8615[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_19 (.CI(n29022), .I0(n8637[16]), .I1(GND_net), .CO(n29023));
    SB_LUT4 i34545_4_lut (.I0(n37_adj_3482), .I1(n35_adj_3490), .I2(n33_adj_3496), 
            .I3(n40425), .O(n40867));
    defparam i34545_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_7_i16_3_lut (.I0(n103[9]), .I1(n103[21]), .I2(n43_adj_3481), 
            .I3(GND_net), .O(n16_adj_3505));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4599_18_lut (.I0(GND_net), .I1(n8637[15]), .I2(GND_net), 
            .I3(n29021), .O(n8615[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_18 (.CI(n29021), .I0(n8637[15]), .I1(GND_net), .CO(n29022));
    SB_LUT4 add_4599_17_lut (.I0(GND_net), .I1(n8637[14]), .I2(GND_net), 
            .I3(n29020), .O(n8615[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_17 (.CI(n29020), .I0(n8637[14]), .I1(GND_net), .CO(n29021));
    SB_LUT4 add_4599_16_lut (.I0(GND_net), .I1(n8637[13]), .I2(GND_net), 
            .I3(n29019), .O(n8615[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_16 (.CI(n29019), .I0(n8637[13]), .I1(GND_net), .CO(n29020));
    SB_LUT4 add_4599_15_lut (.I0(GND_net), .I1(n8637[12]), .I2(GND_net), 
            .I3(n29018), .O(n8615[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_15 (.CI(n29018), .I0(n8637[12]), .I1(GND_net), .CO(n29019));
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[8]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4599_14_lut (.I0(GND_net), .I1(n8637[11]), .I2(GND_net), 
            .I3(n29017), .O(n8615[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_14 (.CI(n29017), .I0(n8637[11]), .I1(GND_net), .CO(n29018));
    SB_LUT4 add_4599_13_lut (.I0(GND_net), .I1(n8637[10]), .I2(GND_net), 
            .I3(n29016), .O(n8615[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_13 (.CI(n29016), .I0(n8637[10]), .I1(GND_net), .CO(n29017));
    SB_LUT4 add_4599_12_lut (.I0(GND_net), .I1(n8637[9]), .I2(GND_net), 
            .I3(n29015), .O(n8615[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34215_3_lut (.I0(n6), .I1(n103[10]), .I2(n21_adj_3501), .I3(GND_net), 
            .O(n40537));   // verilog/motorControl.v(45[19:35])
    defparam i34215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4599_12 (.CI(n29015), .I0(n8637[9]), .I1(GND_net), .CO(n29016));
    SB_LUT4 add_4599_11_lut (.I0(GND_net), .I1(n8637[8]), .I2(GND_net), 
            .I3(n29014), .O(n8615[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34216_3_lut (.I0(n40537), .I1(n103[11]), .I2(n23_adj_3486), 
            .I3(GND_net), .O(n40538));   // verilog/motorControl.v(45[19:35])
    defparam i34216_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4599_11 (.CI(n29014), .I0(n8637[8]), .I1(GND_net), .CO(n29015));
    SB_LUT4 add_4599_10_lut (.I0(GND_net), .I1(n8637[7]), .I2(GND_net), 
            .I3(n29013), .O(n8615[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4599_10 (.CI(n29013), .I0(n8637[7]), .I1(GND_net), .CO(n29014));
    SB_LUT4 add_4599_9_lut (.I0(GND_net), .I1(n8637[6]), .I2(GND_net), 
            .I3(n29012), .O(n8615[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_9 (.CI(n29012), .I0(n8637[6]), .I1(GND_net), .CO(n29013));
    SB_LUT4 mult_4_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4599_8_lut (.I0(GND_net), .I1(n8637[5]), .I2(n521), .I3(n29011), 
            .O(n8615[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_8 (.CI(n29011), .I0(n8637[5]), .I1(n521), .CO(n29012));
    SB_LUT4 add_4599_7_lut (.I0(GND_net), .I1(n8637[4]), .I2(n448), .I3(n29010), 
            .O(n8615[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_7 (.CI(n29010), .I0(n8637[4]), .I1(n448), .CO(n29011));
    SB_LUT4 add_4599_6_lut (.I0(GND_net), .I1(n8637[3]), .I2(n375), .I3(n29009), 
            .O(n8615[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_6 (.CI(n29009), .I0(n8637[3]), .I1(n375), .CO(n29010));
    SB_LUT4 add_4599_5_lut (.I0(GND_net), .I1(n8637[2]), .I2(n302), .I3(n29008), 
            .O(n8615[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_5 (.CI(n29008), .I0(n8637[2]), .I1(n302), .CO(n29009));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n27619), .I0(motor_state[7]), .I1(n1_adj_3559[7]), 
            .CO(n27620));
    SB_LUT4 unary_minus_8_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4599_4_lut (.I0(GND_net), .I1(n8637[1]), .I2(n229), .I3(n29007), 
            .O(n8615[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4599_4 (.CI(n29007), .I0(n8637[1]), .I1(n229), .CO(n29008));
    SB_LUT4 add_4599_3_lut (.I0(GND_net), .I1(n8637[0]), .I2(n156), .I3(n29006), 
            .O(n8615[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[9]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[22]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4599_3 (.CI(n29006), .I0(n8637[0]), .I1(n156), .CO(n29007));
    SB_LUT4 add_4599_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n8615[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4599_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[23]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4599_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n29006));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_3559[6]), .I3(n27618), .O(\PID_CONTROLLER.err_23__N_3354 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n27618), .I0(motor_state[6]), .I1(n1_adj_3559[6]), 
            .CO(n27619));
    SB_LUT4 add_4598_22_lut (.I0(GND_net), .I1(n8615[19]), .I2(GND_net), 
            .I3(n29005), .O(n8592[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4598_21_lut (.I0(GND_net), .I1(n8615[18]), .I2(GND_net), 
            .I3(n29004), .O(n8592[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_21 (.CI(n29004), .I0(n8615[18]), .I1(GND_net), .CO(n29005));
    SB_LUT4 mult_4_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3491));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4598_20_lut (.I0(GND_net), .I1(n8615[17]), .I2(GND_net), 
            .I3(n29003), .O(n8592[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_3559[5]), .I3(n27617), .O(\PID_CONTROLLER.err_23__N_3354 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_20 (.CI(n29003), .I0(n8615[17]), .I1(GND_net), .CO(n29004));
    SB_LUT4 mult_4_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4598_19_lut (.I0(GND_net), .I1(n8615[16]), .I2(GND_net), 
            .I3(n29002), .O(n8592[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4598_19 (.CI(n29002), .I0(n8615[16]), .I1(GND_net), .CO(n29003));
    SB_LUT4 add_4598_18_lut (.I0(GND_net), .I1(n8615[15]), .I2(GND_net), 
            .I3(n29001), .O(n8592[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_18 (.CI(n29001), .I0(n8615[15]), .I1(GND_net), .CO(n29002));
    SB_LUT4 add_4598_17_lut (.I0(GND_net), .I1(n8615[14]), .I2(GND_net), 
            .I3(n29000), .O(n8592[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_17 (.CI(n29000), .I0(n8615[14]), .I1(GND_net), .CO(n29001));
    SB_LUT4 mult_4_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[10]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[11]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n27617), .I0(motor_state[5]), .I1(n1_adj_3559[5]), 
            .CO(n27618));
    SB_LUT4 mult_4_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3475));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_7_i8_3_lut (.I0(n103[4]), .I1(n103[8]), .I2(n17_adj_3499), 
            .I3(GND_net), .O(n8_adj_3507));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i24_3_lut (.I0(n16_adj_3505), .I1(n103[22]), .I2(n45_adj_3480), 
            .I3(GND_net), .O(n24_adj_3508));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33299_4_lut (.I0(n43_adj_3481), .I1(n25_adj_3487), .I2(n23_adj_3486), 
            .I3(n39675), .O(n39621));
    defparam i33299_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34004_4_lut (.I0(n24_adj_3508), .I1(n8_adj_3507), .I2(n45_adj_3480), 
            .I3(n39593), .O(n40326));   // verilog/motorControl.v(45[19:35])
    defparam i34004_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33597_3_lut (.I0(n40538), .I1(n103[12]), .I2(n25_adj_3487), 
            .I3(GND_net), .O(n39919));   // verilog/motorControl.v(45[19:35])
    defparam i33597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_7_i4_4_lut (.I0(n103[0]), .I1(n103[1]), .I2(duty[1]), 
            .I3(duty[0]), .O(n4_adj_3509));   // verilog/motorControl.v(45[19:35])
    defparam LessThan_7_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_4_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34211_3_lut (.I0(n4_adj_3509), .I1(n103[13]), .I2(n27_adj_3489), 
            .I3(GND_net), .O(n40533));   // verilog/motorControl.v(45[19:35])
    defparam i34211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34212_3_lut (.I0(n40533), .I1(n103[14]), .I2(n29_adj_3483), 
            .I3(GND_net), .O(n40534));   // verilog/motorControl.v(45[19:35])
    defparam i34212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33327_4_lut (.I0(n33_adj_3496), .I1(n31_adj_3485), .I2(n29_adj_3483), 
            .I3(n39661), .O(n39649));
    defparam i33327_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34500_4_lut (.I0(n30_adj_3504), .I1(n10_adj_3503), .I2(n35_adj_3490), 
            .I3(n39641), .O(n40822));   // verilog/motorControl.v(45[19:35])
    defparam i34500_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33599_3_lut (.I0(n40534), .I1(n103[15]), .I2(n31_adj_3485), 
            .I3(GND_net), .O(n39921));   // verilog/motorControl.v(45[19:35])
    defparam i33599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34611_4_lut (.I0(n39921), .I1(n40822), .I2(n35_adj_3490), 
            .I3(n39649), .O(n40933));   // verilog/motorControl.v(45[19:35])
    defparam i34611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_4_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34612_3_lut (.I0(n40933), .I1(n103[18]), .I2(n37_adj_3482), 
            .I3(GND_net), .O(n40934));   // verilog/motorControl.v(45[19:35])
    defparam i34612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34582_3_lut (.I0(n40934), .I1(n103[19]), .I2(n39_adj_3479), 
            .I3(GND_net), .O(n40904));   // verilog/motorControl.v(45[19:35])
    defparam i34582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_4_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33301_4_lut (.I0(n43_adj_3481), .I1(n41_adj_3478), .I2(n39_adj_3479), 
            .I3(n40867), .O(n39623));
    defparam i33301_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[12]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34410_4_lut (.I0(n39919), .I1(n40326), .I2(n45_adj_3480), 
            .I3(n39621), .O(n40732));   // verilog/motorControl.v(45[19:35])
    defparam i34410_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4598_16_lut (.I0(GND_net), .I1(n8615[13]), .I2(GND_net), 
            .I3(n28999), .O(n8592[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_16 (.CI(n28999), .I0(n8615[13]), .I1(GND_net), .CO(n29000));
    SB_LUT4 add_4598_15_lut (.I0(GND_net), .I1(n8615[12]), .I2(GND_net), 
            .I3(n28998), .O(n8592[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_15 (.CI(n28998), .I0(n8615[12]), .I1(GND_net), .CO(n28999));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_3559[4]), .I3(n27616), .O(\PID_CONTROLLER.err_23__N_3354 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4598_14_lut (.I0(GND_net), .I1(n8615[11]), .I2(GND_net), 
            .I3(n28997), .O(n8592[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_14 (.CI(n28997), .I0(n8615[11]), .I1(GND_net), .CO(n28998));
    SB_LUT4 add_4598_13_lut (.I0(GND_net), .I1(n8615[10]), .I2(GND_net), 
            .I3(n28996), .O(n8592[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_13 (.CI(n28996), .I0(n8615[10]), .I1(GND_net), .CO(n28997));
    SB_LUT4 add_4598_12_lut (.I0(GND_net), .I1(n8615[9]), .I2(GND_net), 
            .I3(n28995), .O(n8592[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_12 (.CI(n28995), .I0(n8615[9]), .I1(GND_net), .CO(n28996));
    SB_LUT4 i33605_3_lut (.I0(n40904), .I1(n103[20]), .I2(n41_adj_3478), 
            .I3(GND_net), .O(n39927));   // verilog/motorControl.v(45[19:35])
    defparam i33605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4598_11_lut (.I0(GND_net), .I1(n8615[8]), .I2(GND_net), 
            .I3(n28994), .O(n8592[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n27616), .I0(motor_state[4]), .I1(n1_adj_3559[4]), 
            .CO(n27617));
    SB_CARRY add_4598_11 (.CI(n28994), .I0(n8615[8]), .I1(GND_net), .CO(n28995));
    SB_LUT4 add_4598_10_lut (.I0(GND_net), .I1(n8615[7]), .I2(GND_net), 
            .I3(n28993), .O(n8592[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_10 (.CI(n28993), .I0(n8615[7]), .I1(GND_net), .CO(n28994));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_3559[3]), .I3(n27615), .O(\PID_CONTROLLER.err_23__N_3354 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n27615), .I0(motor_state[3]), .I1(n1_adj_3559[3]), 
            .CO(n27616));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_3559[2]), .I3(n27614), .O(\PID_CONTROLLER.err_23__N_3354 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4598_9_lut (.I0(GND_net), .I1(n8615[6]), .I2(GND_net), 
            .I3(n28992), .O(n8592[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_9 (.CI(n28992), .I0(n8615[6]), .I1(GND_net), .CO(n28993));
    SB_LUT4 add_4598_8_lut (.I0(GND_net), .I1(n8615[5]), .I2(n518), .I3(n28991), 
            .O(n8592[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_8 (.CI(n28991), .I0(n8615[5]), .I1(n518), .CO(n28992));
    SB_LUT4 add_4598_7_lut (.I0(GND_net), .I1(n8615[4]), .I2(n445), .I3(n28990), 
            .O(n8592[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_7 (.CI(n28990), .I0(n8615[4]), .I1(n445), .CO(n28991));
    SB_LUT4 add_4598_6_lut (.I0(GND_net), .I1(n8615[3]), .I2(n372), .I3(n28989), 
            .O(n8592[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_6 (.CI(n28989), .I0(n8615[3]), .I1(n372), .CO(n28990));
    SB_LUT4 add_4598_5_lut (.I0(GND_net), .I1(n8615[2]), .I2(n299), .I3(n28988), 
            .O(n8592[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n27614), .I0(motor_state[2]), .I1(n1_adj_3559[2]), 
            .CO(n27615));
    SB_CARRY add_4598_5 (.CI(n28988), .I0(n8615[2]), .I1(n299), .CO(n28989));
    SB_LUT4 add_4598_4_lut (.I0(GND_net), .I1(n8615[1]), .I2(n226), .I3(n28987), 
            .O(n8592[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_4 (.CI(n28987), .I0(n8615[1]), .I1(n226), .CO(n28988));
    SB_LUT4 add_4598_3_lut (.I0(GND_net), .I1(n8615[0]), .I2(n153), .I3(n28986), 
            .O(n8592[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_3 (.CI(n28986), .I0(n8615[0]), .I1(n153), .CO(n28987));
    SB_LUT4 add_4598_2_lut (.I0(GND_net), .I1(n11_adj_3513), .I2(n80), 
            .I3(GND_net), .O(n8592[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4598_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4598_2 (.CI(GND_net), .I0(n11_adj_3513), .I1(n80), .CO(n28986));
    SB_LUT4 mult_4_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n8568[21]), 
            .I2(GND_net), .I3(n28985), .O(n39021)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_4_add_1225_23_lut (.I0(GND_net), .I1(n8568[20]), .I2(GND_net), 
            .I3(n28984), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_23 (.CI(n28984), .I0(n8568[20]), .I1(GND_net), 
            .CO(n28985));
    SB_LUT4 mult_4_add_1225_22_lut (.I0(GND_net), .I1(n8568[19]), .I2(GND_net), 
            .I3(n28983), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_22 (.CI(n28983), .I0(n8568[19]), .I1(GND_net), 
            .CO(n28984));
    SB_LUT4 mult_4_add_1225_21_lut (.I0(GND_net), .I1(n8568[18]), .I2(GND_net), 
            .I3(n28982), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_21 (.CI(n28982), .I0(n8568[18]), .I1(GND_net), 
            .CO(n28983));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_3559[1]), .I3(n27613), .O(\PID_CONTROLLER.err_23__N_3354 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3330[1]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 mult_4_add_1225_20_lut (.I0(GND_net), .I1(n8568[17]), .I2(GND_net), 
            .I3(n28981), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_20 (.CI(n28981), .I0(n8568[17]), .I1(GND_net), 
            .CO(n28982));
    SB_LUT4 mult_4_add_1225_19_lut (.I0(GND_net), .I1(n8568[16]), .I2(GND_net), 
            .I3(n28980), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34532_4_lut (.I0(n39927), .I1(n40732), .I2(n45_adj_3480), 
            .I3(n39623), .O(n40854));   // verilog/motorControl.v(45[19:35])
    defparam i34532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[13]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[14]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[15]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n27613), .I0(motor_state[1]), .I1(n1_adj_3559[1]), 
            .CO(n27614));
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[16]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_4_add_1225_19 (.CI(n28980), .I0(n8568[16]), .I1(GND_net), 
            .CO(n28981));
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3330[2]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 mult_4_add_1225_18_lut (.I0(GND_net), .I1(n8568[15]), .I2(GND_net), 
            .I3(n28979), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3330[3]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3330[4]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3330[5]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3330[6]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3330[7]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3330[8]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3330[9]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3330[10]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3330[11]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3330[12]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3330[13]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3330[14]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3330[15]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3330[16]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3330[17]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3330[18]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3330[19]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3330[20]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3330[21]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3330[22]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3330[23]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [1]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [2]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [3]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [4]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [5]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [6]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [7]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [8]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [9]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [10]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [11]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [12]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [13]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [14]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [15]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [16]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [17]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [18]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [19]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [20]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [21]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [22]));   // verilog/motorControl.v(36[14] 55[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3354 [23]));   // verilog/motorControl.v(36[14] 55[8])
    SB_LUT4 i34533_3_lut (.I0(n40854), .I1(duty[23]), .I2(n103[23]), .I3(GND_net), 
            .O(n102));   // verilog/motorControl.v(45[19:35])
    defparam i34533_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[17]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_4_add_1225_18 (.CI(n28979), .I0(n8568[15]), .I1(GND_net), 
            .CO(n28980));
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[18]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_add_1225_17_lut (.I0(GND_net), .I1(n8568[14]), .I2(GND_net), 
            .I3(n28978), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_17 (.CI(n28978), .I0(n8568[14]), .I1(GND_net), 
            .CO(n28979));
    SB_LUT4 mult_4_add_1225_16_lut (.I0(GND_net), .I1(n8568[13]), .I2(GND_net), 
            .I3(n28977), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_16 (.CI(n28977), .I0(n8568[13]), .I1(GND_net), 
            .CO(n28978));
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[19]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_add_1225_15_lut (.I0(GND_net), .I1(n8568[12]), .I2(GND_net), 
            .I3(n28976), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_9_i1_4_lut (.I0(\PID_CONTROLLER.err [0]), .I1(n103[0]), 
            .I2(n102), .I3(\Kp[0] ), .O(duty_23__N_3378[0]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i1_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 duty_23__I_0_18_i1_3_lut (.I0(duty_23__N_3378[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[0]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[20]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[21]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_4_add_1225_15 (.CI(n28976), .I0(n8568[12]), .I1(GND_net), 
            .CO(n28977));
    SB_LUT4 mult_4_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35388_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n41708));   // verilog/motorControl.v(36[14] 55[8])
    defparam i35388_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_add_1225_14_lut (.I0(GND_net), .I1(n8568[11]), .I2(GND_net), 
            .I3(n28975), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_14 (.CI(n28975), .I0(n8568[11]), .I1(GND_net), 
            .CO(n28976));
    SB_LUT4 mult_4_add_1225_13_lut (.I0(GND_net), .I1(n8568[10]), .I2(GND_net), 
            .I3(n28974), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_13 (.CI(n28974), .I0(n8568[10]), .I1(GND_net), 
            .CO(n28975));
    SB_LUT4 mult_4_add_1225_12_lut (.I0(GND_net), .I1(n8568[9]), .I2(GND_net), 
            .I3(n28973), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_12 (.CI(n28973), .I0(n8568[9]), .I1(GND_net), 
            .CO(n28974));
    SB_LUT4 mult_4_add_1225_11_lut (.I0(GND_net), .I1(n8568[8]), .I2(GND_net), 
            .I3(n28972), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_11 (.CI(n28972), .I0(n8568[8]), .I1(GND_net), 
            .CO(n28973));
    SB_LUT4 mult_4_add_1225_10_lut (.I0(GND_net), .I1(n8568[7]), .I2(GND_net), 
            .I3(n28971), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_10 (.CI(n28971), .I0(n8568[7]), .I1(GND_net), 
            .CO(n28972));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_3559[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3354 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_add_1225_9_lut (.I0(GND_net), .I1(n8568[6]), .I2(GND_net), 
            .I3(n28970), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_9 (.CI(n28970), .I0(n8568[6]), .I1(GND_net), 
            .CO(n28971));
    SB_LUT4 add_4613_7_lut (.I0(GND_net), .I1(n35928), .I2(n490), .I3(n29185), 
            .O(n8832[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_6_lut (.I0(GND_net), .I1(n8840[3]), .I2(n417), .I3(n29184), 
            .O(n8832[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_6 (.CI(n29184), .I0(n8840[3]), .I1(n417), .CO(n29185));
    SB_LUT4 mult_4_add_1225_8_lut (.I0(GND_net), .I1(n8568[5]), .I2(n512), 
            .I3(n28969), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_5_lut (.I0(GND_net), .I1(n8840[2]), .I2(n344), .I3(n29183), 
            .O(n8832[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_8 (.CI(n28969), .I0(n8568[5]), .I1(n512), 
            .CO(n28970));
    SB_CARRY add_4613_5 (.CI(n29183), .I0(n8840[2]), .I1(n344), .CO(n29184));
    SB_LUT4 mult_4_add_1225_7_lut (.I0(GND_net), .I1(n8568[4]), .I2(n439), 
            .I3(n28968), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_7 (.CI(n28968), .I0(n8568[4]), .I1(n439), 
            .CO(n28969));
    SB_LUT4 mult_4_add_1225_6_lut (.I0(GND_net), .I1(n8568[3]), .I2(n366), 
            .I3(n28967), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_4_lut (.I0(GND_net), .I1(n8840[1]), .I2(n271), .I3(n29182), 
            .O(n8832[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_4 (.CI(n29182), .I0(n8840[1]), .I1(n271), .CO(n29183));
    SB_CARRY mult_4_add_1225_6 (.CI(n28967), .I0(n8568[3]), .I1(n366), 
            .CO(n28968));
    SB_LUT4 add_4613_3_lut (.I0(GND_net), .I1(n8840[0]), .I2(n198), .I3(n29181), 
            .O(n8832[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_add_1225_5_lut (.I0(GND_net), .I1(n8568[2]), .I2(n293), 
            .I3(n28966), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_3559[0]), 
            .CO(n27613));
    SB_CARRY mult_4_add_1225_5 (.CI(n28966), .I0(n8568[2]), .I1(n293), 
            .CO(n28967));
    SB_LUT4 mult_4_add_1225_4_lut (.I0(GND_net), .I1(n8568[1]), .I2(n220), 
            .I3(n28965), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n27612), .O(n103[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_4 (.CI(n28965), .I0(n8568[1]), .I1(n220), 
            .CO(n28966));
    SB_CARRY add_4613_3 (.CI(n29181), .I0(n8840[0]), .I1(n198), .CO(n29182));
    SB_LUT4 mult_4_add_1225_3_lut (.I0(GND_net), .I1(n8568[0]), .I2(n147), 
            .I3(n28964), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_2_lut (.I0(GND_net), .I1(n56_adj_3517), .I2(n125_adj_3518), 
            .I3(GND_net), .O(n8832[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_3 (.CI(n28964), .I0(n8568[0]), .I1(n147), 
            .CO(n28965));
    SB_CARRY add_4613_2 (.CI(GND_net), .I0(n56_adj_3517), .I1(n125_adj_3518), 
            .CO(n29181));
    SB_LUT4 mult_4_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3519), .I2(n74_adj_3520), 
            .I3(GND_net), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_4_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_8_lut (.I0(GND_net), .I1(n8832[5]), .I2(n560), .I3(n29180), 
            .O(n8823[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_7_lut (.I0(GND_net), .I1(n8832[4]), .I2(n487), .I3(n29179), 
            .O(n8823[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_4_add_1225_2 (.CI(GND_net), .I0(n5_adj_3519), .I1(n74_adj_3520), 
            .CO(n28964));
    SB_CARRY add_4612_7 (.CI(n29179), .I0(n8832[4]), .I1(n487), .CO(n29180));
    SB_LUT4 add_4612_6_lut (.I0(GND_net), .I1(n8832[3]), .I2(n414), .I3(n29178), 
            .O(n8823[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_6 (.CI(n29178), .I0(n8832[3]), .I1(n414), .CO(n29179));
    SB_LUT4 add_4612_5_lut (.I0(GND_net), .I1(n8832[2]), .I2(n341), .I3(n29177), 
            .O(n8823[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_5 (.CI(n29177), .I0(n8832[2]), .I1(n341), .CO(n29178));
    SB_LUT4 add_4612_4_lut (.I0(GND_net), .I1(n8832[1]), .I2(n268), .I3(n29176), 
            .O(n8823[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_4 (.CI(n29176), .I0(n8832[1]), .I1(n268), .CO(n29177));
    SB_LUT4 add_4612_3_lut (.I0(GND_net), .I1(n8832[0]), .I2(n195), .I3(n29175), 
            .O(n8823[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_3 (.CI(n29175), .I0(n8832[0]), .I1(n195), .CO(n29176));
    SB_LUT4 add_4612_2_lut (.I0(GND_net), .I1(n53_adj_3521), .I2(n122_adj_3522), 
            .I3(GND_net), .O(n8823[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_2 (.CI(GND_net), .I0(n53_adj_3521), .I1(n122_adj_3522), 
            .CO(n29175));
    SB_LUT4 add_4611_9_lut (.I0(GND_net), .I1(n8823[6]), .I2(GND_net), 
            .I3(n29174), .O(n8813[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_8_lut (.I0(GND_net), .I1(n8823[5]), .I2(n557), .I3(n29173), 
            .O(n8813[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_8 (.CI(n29173), .I0(n8823[5]), .I1(n557), .CO(n29174));
    SB_LUT4 add_4611_7_lut (.I0(GND_net), .I1(n8823[4]), .I2(n484), .I3(n29172), 
            .O(n8813[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_7 (.CI(n29172), .I0(n8823[4]), .I1(n484), .CO(n29173));
    SB_LUT4 add_4611_6_lut (.I0(GND_net), .I1(n8823[3]), .I2(n411), .I3(n29171), 
            .O(n8813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_6 (.CI(n29171), .I0(n8823[3]), .I1(n411), .CO(n29172));
    SB_LUT4 add_4611_5_lut (.I0(GND_net), .I1(n8823[2]), .I2(n338), .I3(n29170), 
            .O(n8813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n27611), .O(n103[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_5 (.CI(n29170), .I0(n8823[2]), .I1(n338), .CO(n29171));
    SB_LUT4 add_4611_4_lut (.I0(GND_net), .I1(n8823[1]), .I2(n265), .I3(n29169), 
            .O(n8813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_4 (.CI(n29169), .I0(n8823[1]), .I1(n265), .CO(n29170));
    SB_LUT4 add_4611_3_lut (.I0(GND_net), .I1(n8823[0]), .I2(n192), .I3(n29168), 
            .O(n8813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_3 (.CI(n29168), .I0(n8823[0]), .I1(n192), .CO(n29169));
    SB_LUT4 add_4611_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_3524), 
            .I3(GND_net), .O(n8813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_3524), .CO(n29168));
    SB_LUT4 add_4610_10_lut (.I0(GND_net), .I1(n8813[7]), .I2(GND_net), 
            .I3(n29167), .O(n8802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_9_lut (.I0(GND_net), .I1(n8813[6]), .I2(GND_net), 
            .I3(n29166), .O(n8802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_9 (.CI(n29166), .I0(n8813[6]), .I1(GND_net), .CO(n29167));
    SB_LUT4 add_4610_8_lut (.I0(GND_net), .I1(n8813[5]), .I2(n554), .I3(n29165), 
            .O(n8802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_24 (.CI(n27611), .I0(GND_net), .I1(n1[22]), 
            .CO(n27612));
    SB_CARRY add_4610_8 (.CI(n29165), .I0(n8813[5]), .I1(n554), .CO(n29166));
    SB_LUT4 add_4610_7_lut (.I0(GND_net), .I1(n8813[4]), .I2(n481), .I3(n29164), 
            .O(n8802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n27610), .O(n103[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_7 (.CI(n29164), .I0(n8813[4]), .I1(n481), .CO(n29165));
    SB_LUT4 add_4610_6_lut (.I0(GND_net), .I1(n8813[3]), .I2(n408), .I3(n29163), 
            .O(n8802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_6 (.CI(n29163), .I0(n8813[3]), .I1(n408), .CO(n29164));
    SB_LUT4 add_4610_5_lut (.I0(GND_net), .I1(n8813[2]), .I2(n335), .I3(n29162), 
            .O(n8802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_5 (.CI(n29162), .I0(n8813[2]), .I1(n335), .CO(n29163));
    SB_LUT4 add_4610_4_lut (.I0(GND_net), .I1(n8813[1]), .I2(n262), .I3(n29161), 
            .O(n8802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_23 (.CI(n27610), .I0(GND_net), .I1(n1[21]), 
            .CO(n27611));
    SB_CARRY add_4610_4 (.CI(n29161), .I0(n8813[1]), .I1(n262), .CO(n29162));
    SB_LUT4 unary_minus_8_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n27609), .O(n103[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_3_lut (.I0(GND_net), .I1(n8813[0]), .I2(n189), .I3(n29160), 
            .O(n8802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_3 (.CI(n29160), .I0(n8813[0]), .I1(n189), .CO(n29161));
    SB_LUT4 add_4610_2_lut (.I0(GND_net), .I1(n47), .I2(n116_adj_3527), 
            .I3(GND_net), .O(n8802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_2 (.CI(GND_net), .I0(n47), .I1(n116_adj_3527), .CO(n29160));
    SB_LUT4 add_4609_11_lut (.I0(GND_net), .I1(n8802[8]), .I2(GND_net), 
            .I3(n29159), .O(n8790[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4609_10_lut (.I0(GND_net), .I1(n8802[7]), .I2(GND_net), 
            .I3(n29158), .O(n8790[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_10 (.CI(n29158), .I0(n8802[7]), .I1(GND_net), .CO(n29159));
    SB_CARRY unary_minus_8_add_3_22 (.CI(n27609), .I0(GND_net), .I1(n1[20]), 
            .CO(n27610));
    SB_LUT4 unary_minus_8_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n27608), .O(n103[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4609_9_lut (.I0(GND_net), .I1(n8802[6]), .I2(GND_net), 
            .I3(n29157), .O(n8790[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_9 (.CI(n29157), .I0(n8802[6]), .I1(GND_net), .CO(n29158));
    SB_CARRY unary_minus_8_add_3_21 (.CI(n27608), .I0(GND_net), .I1(n1[19]), 
            .CO(n27609));
    SB_LUT4 add_4609_8_lut (.I0(GND_net), .I1(n8802[5]), .I2(n551), .I3(n29156), 
            .O(n8790[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_8 (.CI(n29156), .I0(n8802[5]), .I1(n551), .CO(n29157));
    SB_LUT4 add_4609_7_lut (.I0(GND_net), .I1(n8802[4]), .I2(n478), .I3(n29155), 
            .O(n8790[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_7 (.CI(n29155), .I0(n8802[4]), .I1(n478), .CO(n29156));
    SB_LUT4 add_4609_6_lut (.I0(GND_net), .I1(n8802[3]), .I2(n405), .I3(n29154), 
            .O(n8790[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n27607), .O(n103[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_6 (.CI(n29154), .I0(n8802[3]), .I1(n405), .CO(n29155));
    SB_CARRY unary_minus_8_add_3_20 (.CI(n27607), .I0(GND_net), .I1(n1[18]), 
            .CO(n27608));
    SB_LUT4 add_4609_5_lut (.I0(GND_net), .I1(n8802[2]), .I2(n332), .I3(n29153), 
            .O(n8790[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_5 (.CI(n29153), .I0(n8802[2]), .I1(n332), .CO(n29154));
    SB_LUT4 unary_minus_8_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n27606), .O(n103[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4609_4_lut (.I0(GND_net), .I1(n8802[1]), .I2(n259), .I3(n29152), 
            .O(n8790[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_4 (.CI(n29152), .I0(n8802[1]), .I1(n259), .CO(n29153));
    SB_LUT4 add_4609_3_lut (.I0(GND_net), .I1(n8802[0]), .I2(n186), .I3(n29151), 
            .O(n8790[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_3 (.CI(n29151), .I0(n8802[0]), .I1(n186), .CO(n29152));
    SB_LUT4 add_4609_2_lut (.I0(GND_net), .I1(n44), .I2(n113_adj_3531), 
            .I3(GND_net), .O(n8790[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_2 (.CI(GND_net), .I0(n44), .I1(n113_adj_3531), .CO(n29151));
    SB_LUT4 add_4608_12_lut (.I0(GND_net), .I1(n8790[9]), .I2(GND_net), 
            .I3(n29150), .O(n8777[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_11_lut (.I0(GND_net), .I1(n8790[8]), .I2(GND_net), 
            .I3(n29149), .O(n8777[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_11 (.CI(n29149), .I0(n8790[8]), .I1(GND_net), .CO(n29150));
    SB_LUT4 add_4608_10_lut (.I0(GND_net), .I1(n8790[7]), .I2(GND_net), 
            .I3(n29148), .O(n8777[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_10 (.CI(n29148), .I0(n8790[7]), .I1(GND_net), .CO(n29149));
    SB_LUT4 add_4608_9_lut (.I0(GND_net), .I1(n8790[6]), .I2(GND_net), 
            .I3(n29147), .O(n8777[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_9 (.CI(n29147), .I0(n8790[6]), .I1(GND_net), .CO(n29148));
    SB_CARRY unary_minus_8_add_3_19 (.CI(n27606), .I0(GND_net), .I1(n1[17]), 
            .CO(n27607));
    SB_LUT4 add_4608_8_lut (.I0(GND_net), .I1(n8790[5]), .I2(n548), .I3(n29146), 
            .O(n8777[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_8 (.CI(n29146), .I0(n8790[5]), .I1(n548), .CO(n29147));
    SB_LUT4 unary_minus_8_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n27605), .O(n103[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4608_7_lut (.I0(GND_net), .I1(n8790[4]), .I2(n475), .I3(n29145), 
            .O(n8777[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4608_7 (.CI(n29145), .I0(n8790[4]), .I1(n475), .CO(n29146));
    SB_LUT4 add_4608_6_lut (.I0(GND_net), .I1(n8790[3]), .I2(n402), .I3(n29144), 
            .O(n8777[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_6 (.CI(n29144), .I0(n8790[3]), .I1(n402), .CO(n29145));
    SB_LUT4 add_4608_5_lut (.I0(GND_net), .I1(n8790[2]), .I2(n329), .I3(n29143), 
            .O(n8777[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_5 (.CI(n29143), .I0(n8790[2]), .I1(n329), .CO(n29144));
    SB_LUT4 add_4608_4_lut (.I0(GND_net), .I1(n8790[1]), .I2(n256), .I3(n29142), 
            .O(n8777[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4608_4 (.CI(n29142), .I0(n8790[1]), .I1(n256), .CO(n29143));
    SB_LUT4 mult_4_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4608_3_lut (.I0(GND_net), .I1(n8790[0]), .I2(n183), .I3(n29141), 
            .O(n8777[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_3 (.CI(n29141), .I0(n8790[0]), .I1(n183), .CO(n29142));
    SB_LUT4 unary_minus_8_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4608_2_lut (.I0(GND_net), .I1(n41_adj_3535), .I2(n110_adj_3536), 
            .I3(GND_net), .O(n8777[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_2 (.CI(GND_net), .I0(n41_adj_3535), .I1(n110_adj_3536), 
            .CO(n29141));
    SB_LUT4 add_4607_13_lut (.I0(GND_net), .I1(n8777[10]), .I2(GND_net), 
            .I3(n29140), .O(n8763[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_12_lut (.I0(GND_net), .I1(n8777[9]), .I2(GND_net), 
            .I3(n29139), .O(n8763[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4607_12 (.CI(n29139), .I0(n8777[9]), .I1(GND_net), .CO(n29140));
    SB_LUT4 add_4607_11_lut (.I0(GND_net), .I1(n8777[8]), .I2(GND_net), 
            .I3(n29138), .O(n8763[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_8_add_3_18 (.CI(n27605), .I0(GND_net), .I1(n1[16]), 
            .CO(n27606));
    SB_CARRY add_4607_11 (.CI(n29138), .I0(n8777[8]), .I1(GND_net), .CO(n29139));
    SB_LUT4 unary_minus_8_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n27604), .O(n103[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_10_lut (.I0(GND_net), .I1(n8777[7]), .I2(GND_net), 
            .I3(n29137), .O(n8763[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4607_10 (.CI(n29137), .I0(n8777[7]), .I1(GND_net), .CO(n29138));
    SB_LUT4 add_4607_9_lut (.I0(GND_net), .I1(n8777[6]), .I2(GND_net), 
            .I3(n29136), .O(n8763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_9 (.CI(n29136), .I0(n8777[6]), .I1(GND_net), .CO(n29137));
    SB_LUT4 unary_minus_8_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4607_8_lut (.I0(GND_net), .I1(n8777[5]), .I2(n545), .I3(n29135), 
            .O(n8763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_8 (.CI(n29135), .I0(n8777[5]), .I1(n545), .CO(n29136));
    SB_LUT4 mult_4_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_8_add_3_17 (.CI(n27604), .I0(GND_net), .I1(n1[15]), 
            .CO(n27605));
    SB_LUT4 add_4607_7_lut (.I0(GND_net), .I1(n8777[4]), .I2(n472), .I3(n29134), 
            .O(n8763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n27603), .O(n103[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_16 (.CI(n27603), .I0(GND_net), .I1(n1[14]), 
            .CO(n27604));
    SB_CARRY add_4607_7 (.CI(n29134), .I0(n8777[4]), .I1(n472), .CO(n29135));
    SB_LUT4 add_4607_6_lut (.I0(GND_net), .I1(n8777[3]), .I2(n399), .I3(n29133), 
            .O(n8763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n27602), .O(n103[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_6 (.CI(n29133), .I0(n8777[3]), .I1(n399), .CO(n29134));
    SB_CARRY unary_minus_8_add_3_15 (.CI(n27602), .I0(GND_net), .I1(n1[13]), 
            .CO(n27603));
    SB_LUT4 unary_minus_8_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n27601), .O(n103[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_14 (.CI(n27601), .I0(GND_net), .I1(n1[12]), 
            .CO(n27602));
    SB_LUT4 unary_minus_8_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n27600), .O(n103[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3543));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3544));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4607_5_lut (.I0(GND_net), .I1(n8777[2]), .I2(n326), .I3(n29132), 
            .O(n8763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_5 (.CI(n29132), .I0(n8777[2]), .I1(n326), .CO(n29133));
    SB_LUT4 add_4607_4_lut (.I0(GND_net), .I1(n8777[1]), .I2(n253), .I3(n29131), 
            .O(n8763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_4 (.CI(n29131), .I0(n8777[1]), .I1(n253), .CO(n29132));
    SB_LUT4 add_4607_3_lut (.I0(GND_net), .I1(n8777[0]), .I2(n180), .I3(n29130), 
            .O(n8763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_3 (.CI(n29130), .I0(n8777[0]), .I1(n180), .CO(n29131));
    SB_LUT4 mult_4_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4607_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_3545), 
            .I3(GND_net), .O(n8763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_8_add_3_13 (.CI(n27600), .I0(GND_net), .I1(n1[11]), 
            .CO(n27601));
    SB_CARRY add_4607_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_3545), .CO(n29130));
    SB_LUT4 mult_4_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4606_14_lut (.I0(GND_net), .I1(n8763[11]), .I2(GND_net), 
            .I3(n29129), .O(n8748[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_13_lut (.I0(GND_net), .I1(n8763[10]), .I2(GND_net), 
            .I3(n29128), .O(n8748[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_13 (.CI(n29128), .I0(n8763[10]), .I1(GND_net), .CO(n29129));
    SB_LUT4 unary_minus_8_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n27599), .O(n103[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_12_lut (.I0(GND_net), .I1(n8763[9]), .I2(GND_net), 
            .I3(n29127), .O(n8748[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4606_12 (.CI(n29127), .I0(n8763[9]), .I1(GND_net), .CO(n29128));
    SB_LUT4 add_4606_11_lut (.I0(GND_net), .I1(n8763[8]), .I2(GND_net), 
            .I3(n29126), .O(n8748[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_12 (.CI(n27599), .I0(GND_net), .I1(n1[10]), 
            .CO(n27600));
    SB_CARRY add_4606_11 (.CI(n29126), .I0(n8763[8]), .I1(GND_net), .CO(n29127));
    SB_LUT4 unary_minus_8_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n27598), .O(n103[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_10_lut (.I0(GND_net), .I1(n8763[7]), .I2(GND_net), 
            .I3(n29125), .O(n8748[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_10 (.CI(n29125), .I0(n8763[7]), .I1(GND_net), .CO(n29126));
    SB_CARRY unary_minus_8_add_3_11 (.CI(n27598), .I0(GND_net), .I1(n1[9]), 
            .CO(n27599));
    SB_LUT4 add_4606_9_lut (.I0(GND_net), .I1(n8763[6]), .I2(GND_net), 
            .I3(n29124), .O(n8748[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_9 (.CI(n29124), .I0(n8763[6]), .I1(GND_net), .CO(n29125));
    SB_LUT4 add_4606_8_lut (.I0(GND_net), .I1(n8763[5]), .I2(n542), .I3(n29123), 
            .O(n8748[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_8 (.CI(n29123), .I0(n8763[5]), .I1(n542), .CO(n29124));
    SB_LUT4 add_4606_7_lut (.I0(GND_net), .I1(n8763[4]), .I2(n469), .I3(n29122), 
            .O(n8748[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_7 (.CI(n29122), .I0(n8763[4]), .I1(n469), .CO(n29123));
    SB_LUT4 unary_minus_8_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n27597), .O(n103[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_6_lut (.I0(GND_net), .I1(n8763[3]), .I2(n396), .I3(n29121), 
            .O(n8748[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_4_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i365_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4606_6 (.CI(n29121), .I0(n8763[3]), .I1(n396), .CO(n29122));
    SB_LUT4 add_4606_5_lut (.I0(GND_net), .I1(n8763[2]), .I2(n323), .I3(n29120), 
            .O(n8748[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_5 (.CI(n29120), .I0(n8763[2]), .I1(n323), .CO(n29121));
    SB_LUT4 add_4606_4_lut (.I0(GND_net), .I1(n8763[1]), .I2(n250), .I3(n29119), 
            .O(n8748[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_4 (.CI(n29119), .I0(n8763[1]), .I1(n250), .CO(n29120));
    SB_LUT4 add_4606_3_lut (.I0(GND_net), .I1(n8763[0]), .I2(n177), .I3(n29118), 
            .O(n8748[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_3 (.CI(n29118), .I0(n8763[0]), .I1(n177), .CO(n29119));
    SB_LUT4 add_4606_2_lut (.I0(GND_net), .I1(n35_adj_3544), .I2(n104_adj_3543), 
            .I3(GND_net), .O(n8748[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_2 (.CI(GND_net), .I0(n35_adj_3544), .I1(n104_adj_3543), 
            .CO(n29118));
    SB_LUT4 add_4605_15_lut (.I0(GND_net), .I1(n8748[12]), .I2(GND_net), 
            .I3(n29117), .O(n8732[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4605_14_lut (.I0(GND_net), .I1(n8748[11]), .I2(GND_net), 
            .I3(n29116), .O(n8732[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_14 (.CI(n29116), .I0(n8748[11]), .I1(GND_net), .CO(n29117));
    SB_LUT4 add_4605_13_lut (.I0(GND_net), .I1(n8748[10]), .I2(GND_net), 
            .I3(n29115), .O(n8732[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_13 (.CI(n29115), .I0(n8748[10]), .I1(GND_net), .CO(n29116));
    SB_LUT4 add_4605_12_lut (.I0(GND_net), .I1(n8748[9]), .I2(GND_net), 
            .I3(n29114), .O(n8732[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_12 (.CI(n29114), .I0(n8748[9]), .I1(GND_net), .CO(n29115));
    SB_LUT4 add_4605_11_lut (.I0(GND_net), .I1(n8748[8]), .I2(GND_net), 
            .I3(n29113), .O(n8732[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_11 (.CI(n29113), .I0(n8748[8]), .I1(GND_net), .CO(n29114));
    SB_LUT4 add_4605_10_lut (.I0(GND_net), .I1(n8748[7]), .I2(GND_net), 
            .I3(n29112), .O(n8732[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_10 (.CI(n29112), .I0(n8748[7]), .I1(GND_net), .CO(n29113));
    SB_LUT4 add_4605_9_lut (.I0(GND_net), .I1(n8748[6]), .I2(GND_net), 
            .I3(n29111), .O(n8732[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_9 (.CI(n29111), .I0(n8748[6]), .I1(GND_net), .CO(n29112));
    SB_LUT4 add_4605_8_lut (.I0(GND_net), .I1(n8748[5]), .I2(n539), .I3(n29110), 
            .O(n8732[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_10 (.CI(n27597), .I0(GND_net), .I1(n1[8]), 
            .CO(n27598));
    SB_LUT4 unary_minus_8_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n27596), .O(n103[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_8 (.CI(n29110), .I0(n8748[5]), .I1(n539), .CO(n29111));
    SB_LUT4 add_4605_7_lut (.I0(GND_net), .I1(n8748[4]), .I2(n466), .I3(n29109), 
            .O(n8732[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4605_7 (.CI(n29109), .I0(n8748[4]), .I1(n466), .CO(n29110));
    SB_LUT4 mult_4_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3545));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4605_6_lut (.I0(GND_net), .I1(n8748[3]), .I2(n393), .I3(n29108), 
            .O(n8732[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_9 (.CI(n27596), .I0(GND_net), .I1(n1[7]), 
            .CO(n27597));
    SB_LUT4 mult_4_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4605_6 (.CI(n29108), .I0(n8748[3]), .I1(n393), .CO(n29109));
    SB_LUT4 add_4605_5_lut (.I0(GND_net), .I1(n8748[2]), .I2(n320), .I3(n29107), 
            .O(n8732[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_5 (.CI(n29107), .I0(n8748[2]), .I1(n320), .CO(n29108));
    SB_LUT4 unary_minus_8_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n27595), .O(n103[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_8_add_3_8 (.CI(n27595), .I0(GND_net), .I1(n1[6]), 
            .CO(n27596));
    SB_LUT4 add_4605_4_lut (.I0(GND_net), .I1(n8748[1]), .I2(n247), .I3(n29106), 
            .O(n8732[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_8_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n27594), .O(n103[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_8_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_4 (.CI(n29106), .I0(n8748[1]), .I1(n247), .CO(n29107));
    SB_CARRY unary_minus_8_add_3_7 (.CI(n27594), .I0(GND_net), .I1(n1[5]), 
            .CO(n27595));
    SB_LUT4 add_4605_3_lut (.I0(GND_net), .I1(n8748[0]), .I2(n174), .I3(n29105), 
            .O(n8732[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_3 (.CI(n29105), .I0(n8748[0]), .I1(n174), .CO(n29106));
    SB_LUT4 unary_minus_8_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4605_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8732[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29105));
    SB_LUT4 mult_4_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3536));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3535));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3531));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_8_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3527));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3524));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3522));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3521));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3520));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3519));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3518));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3517));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_8_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(46[19:28])
    defparam unary_minus_8_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_4_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_3549), .I1(\Kp[4] ), .I2(n8847[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8840[3]));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 i2_4_lut_adj_841 (.I0(n4_adj_3550), .I1(\Kp[3] ), .I2(n8853[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8847[2]));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut_adj_841.LUT_INIT = 16'h965a;
    SB_LUT4 mult_4_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(GND_net), .I3(GND_net), .O(n207));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22962_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8858[0]));   // verilog/motorControl.v(41[17:23])
    defparam i22962_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_3_lut (.I0(n27395), .I1(n207), .I2(n8858[0]), .I3(GND_net), 
            .O(n8853[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_4_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22929_4_lut (.I0(n8853[1]), .I1(\Kp[3] ), .I2(n4_adj_3550), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_3551));   // verilog/motorControl.v(41[17:23])
    defparam i22929_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22964_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n27420));   // verilog/motorControl.v(41[17:23])
    defparam i22964_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_3_lut (.I0(n6_adj_3551), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [20]), 
            .I3(GND_net), .O(n14_adj_3552));   // verilog/motorControl.v(41[17:23])
    defparam i4_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22898_4_lut (.I0(n8847[2]), .I1(\Kp[4] ), .I2(n6_adj_3549), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_3553));   // verilog/motorControl.v(41[17:23])
    defparam i22898_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i2_4_lut_adj_842 (.I0(\Kp[0] ), .I1(\Kp[5] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [18]), .O(n12_adj_3554));   // verilog/motorControl.v(41[17:23])
    defparam i2_4_lut_adj_842.LUT_INIT = 16'h9c50;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_3555));   // verilog/motorControl.v(41[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i5_4_lut (.I0(n8858[0]), .I1(n27420), .I2(n207), .I3(n27395), 
            .O(n15_adj_3556));   // verilog/motorControl.v(41[17:23])
    defparam i5_4_lut.LUT_INIT = 16'h366c;
    SB_LUT4 i7_4_lut (.I0(n8_adj_3553), .I1(n14_adj_3552), .I2(\Kp[1] ), 
            .I3(\PID_CONTROLLER.err [22]), .O(n17_adj_3557));   // verilog/motorControl.v(41[17:23])
    defparam i7_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 i9_4_lut (.I0(n17_adj_3557), .I1(n15_adj_3556), .I2(n11_adj_3555), 
            .I3(n12_adj_3554), .O(n35928));   // verilog/motorControl.v(41[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[0]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33037_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n39357));   // verilog/motorControl.v(43[10:25])
    defparam i33037_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3470));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i22921_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n27361), .I3(n8853[0]), .O(n4_adj_3550));   // verilog/motorControl.v(41[17:23])
    defparam i22921_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n8853[0]), .I3(n27361), .O(n8847[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i22908_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n8847[0]));   // verilog/motorControl.v(41[17:23])
    defparam i22908_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22910_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n27361));   // verilog/motorControl.v(41[17:23])
    defparam i22910_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22941_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n27395));   // verilog/motorControl.v(41[17:23])
    defparam i22941_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22939_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8853[0]));   // verilog/motorControl.v(41[17:23])
    defparam i22939_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22890_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_3558), .I3(n8847[1]), .O(n6_adj_3549));   // verilog/motorControl.v(41[17:23])
    defparam i22890_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_843 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8847[1]), .I3(n4_adj_3558), .O(n8840[2]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut_adj_843.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_844 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8847[0]), .I3(n27318), .O(n8840[1]));   // verilog/motorControl.v(41[17:23])
    defparam i2_3_lut_4_lut_adj_844.LUT_INIT = 16'h8778;
    SB_LUT4 i22882_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n27318), .I3(n8847[0]), .O(n4_adj_3558));   // verilog/motorControl.v(41[17:23])
    defparam i22882_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i22871_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n27318));   // verilog/motorControl.v(41[17:23])
    defparam i22871_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22869_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8840[0]));   // verilog/motorControl.v(41[17:23])
    defparam i22869_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_9_i24_3_lut (.I0(n39021), .I1(n103[23]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[23]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i24_3_lut (.I0(duty_23__N_3378[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[23]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i23_3_lut (.I0(n28[22]), .I1(n103[22]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[22]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i23_3_lut (.I0(duty_23__N_3378[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[22]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i22_3_lut (.I0(n28[21]), .I1(n103[21]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[21]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i22_3_lut (.I0(duty_23__N_3378[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[21]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i21_3_lut (.I0(n28[20]), .I1(n103[20]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[20]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i21_3_lut (.I0(duty_23__N_3378[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[20]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i20_3_lut (.I0(n28[19]), .I1(n103[19]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[19]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i20_3_lut (.I0(duty_23__N_3378[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[19]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i19_3_lut (.I0(n28[18]), .I1(n103[18]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[18]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i19_3_lut (.I0(duty_23__N_3378[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[18]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i18_3_lut (.I0(n28[17]), .I1(n103[17]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[17]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i18_3_lut (.I0(duty_23__N_3378[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[17]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i17_3_lut (.I0(n28[16]), .I1(n103[16]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[16]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i17_3_lut (.I0(duty_23__N_3378[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[16]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i16_3_lut (.I0(n28[15]), .I1(n103[15]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[15]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i16_3_lut (.I0(duty_23__N_3378[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[15]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i15_3_lut (.I0(n28[14]), .I1(n103[14]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[14]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i15_3_lut (.I0(duty_23__N_3378[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[14]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i14_3_lut (.I0(n28[13]), .I1(n103[13]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[13]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i14_3_lut (.I0(duty_23__N_3378[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[13]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i13_3_lut (.I0(n28[12]), .I1(n103[12]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[12]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i13_3_lut (.I0(duty_23__N_3378[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[12]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i12_3_lut (.I0(n28[11]), .I1(n103[11]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[11]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i12_3_lut (.I0(duty_23__N_3378[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[11]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i11_3_lut (.I0(n28[10]), .I1(n103[10]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[10]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i11_3_lut (.I0(duty_23__N_3378[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[10]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i10_3_lut (.I0(n28[9]), .I1(n103[9]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[9]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i10_3_lut (.I0(duty_23__N_3378[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[9]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i9_3_lut (.I0(n28[8]), .I1(n103[8]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[8]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i9_3_lut (.I0(duty_23__N_3378[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[8]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i8_3_lut (.I0(n28[7]), .I1(n103[7]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[7]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i8_3_lut (.I0(duty_23__N_3378[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[7]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i7_3_lut (.I0(n28[6]), .I1(n103[6]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[6]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i7_3_lut (.I0(duty_23__N_3378[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[6]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i6_3_lut (.I0(n28[5]), .I1(n103[5]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[5]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i6_3_lut (.I0(duty_23__N_3378[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[5]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i5_3_lut (.I0(n28[4]), .I1(n103[4]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[4]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i5_3_lut (.I0(duty_23__N_3378[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[4]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i4_3_lut (.I0(n28[3]), .I1(n103[3]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[3]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i4_3_lut (.I0(duty_23__N_3378[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[3]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i3_3_lut (.I0(n28[2]), .I1(n103[2]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[2]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i3_3_lut (.I0(duty_23__N_3378[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[2]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_9_i2_3_lut (.I0(n28[1]), .I1(n103[1]), .I2(n102), .I3(GND_net), 
            .O(duty_23__N_3378[1]));   // verilog/motorControl.v(45[16] 47[10])
    defparam mux_9_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_18_i2_3_lut (.I0(duty_23__N_3378[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3402), .I3(GND_net), .O(duty_23__N_3330[1]));   // verilog/motorControl.v(45[16] 47[10])
    defparam duty_23__I_0_18_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[1]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33271_2_lut_4_lut (.I0(duty[21]), .I1(n103[21]), .I2(duty[9]), 
            .I3(n103[9]), .O(n39593));
    defparam i33271_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i33319_2_lut_4_lut (.I0(duty[16]), .I1(n103[16]), .I2(duty[7]), 
            .I3(n103[7]), .O(n39641));
    defparam i33319_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i4_4_lut_4_lut (.I0(PWMLimit[0]), .I1(duty[1]), 
            .I2(PWMLimit[1]), .I3(duty[0]), .O(n4_adj_3474));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i4_4_lut_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3473));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33383_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n39705));
    defparam i33383_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_3476));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33419_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n39741));
    defparam i33419_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(43[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_4_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3513));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_4_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(41[17:23])
    defparam mult_4_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[2]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[3]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[4]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3559[5]));   // verilog/motorControl.v(37[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n18494, encoder1_position, clk32MHz, 
            n18495, n18475, n18476, n18477, n18478, n18479, n18480, 
            n18496, n18497, n18492, n18493, n18490, n18491, n18488, 
            n18489, n18486, n18487, n18484, n18485, n18481, n18482, 
            n18483, data_o, count_enable, n17899, n2681, GND_net, 
            n18510, PIN_6_c_0, reg_B, PIN_7_c_1, n34961, n17911) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18494;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n18495;
    input n18475;
    input n18476;
    input n18477;
    input n18478;
    input n18479;
    input n18480;
    input n18496;
    input n18497;
    input n18492;
    input n18493;
    input n18490;
    input n18491;
    input n18488;
    input n18489;
    input n18486;
    input n18487;
    input n18484;
    input n18485;
    input n18481;
    input n18482;
    input n18483;
    output [1:0]data_o;
    output count_enable;
    input n17899;
    output [23:0]n2681;
    input GND_net;
    input n18510;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    output n34961;
    input n17911;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2671, n27690, n27689, n27688, n27687, 
        n27686, n27685, n27684, n27683, n27682, n27681, n27680, 
        n27679, n27678, n27677, n27676, n27675, n27674, n27673, 
        n27672, n27671, n27670, n27669, n27668, count_direction, 
        n27667;
    
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18494));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18495));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n18475));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n18476));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n18477));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n18478));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n18479));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n18480));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18496));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18497));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18492));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18493));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18490));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18491));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18488));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18489));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18486));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18487));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n18484));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18485));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n18481));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n18482));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n18483));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17899));   // quad.v(35[10] 41[6])
    SB_LUT4 add_593_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2671), 
            .I3(n27690), .O(n2681[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_593_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2671), 
            .I3(n27689), .O(n2681[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_24 (.CI(n27689), .I0(encoder1_position[22]), .I1(n2671), 
            .CO(n27690));
    SB_LUT4 add_593_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2671), 
            .I3(n27688), .O(n2681[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_23 (.CI(n27688), .I0(encoder1_position[21]), .I1(n2671), 
            .CO(n27689));
    SB_LUT4 add_593_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2671), 
            .I3(n27687), .O(n2681[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_22 (.CI(n27687), .I0(encoder1_position[20]), .I1(n2671), 
            .CO(n27688));
    SB_LUT4 add_593_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2671), 
            .I3(n27686), .O(n2681[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_21 (.CI(n27686), .I0(encoder1_position[19]), .I1(n2671), 
            .CO(n27687));
    SB_LUT4 add_593_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2671), 
            .I3(n27685), .O(n2681[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_20 (.CI(n27685), .I0(encoder1_position[18]), .I1(n2671), 
            .CO(n27686));
    SB_LUT4 add_593_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2671), 
            .I3(n27684), .O(n2681[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_19 (.CI(n27684), .I0(encoder1_position[17]), .I1(n2671), 
            .CO(n27685));
    SB_LUT4 add_593_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2671), 
            .I3(n27683), .O(n2681[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_18 (.CI(n27683), .I0(encoder1_position[16]), .I1(n2671), 
            .CO(n27684));
    SB_LUT4 add_593_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2671), 
            .I3(n27682), .O(n2681[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_17 (.CI(n27682), .I0(encoder1_position[15]), .I1(n2671), 
            .CO(n27683));
    SB_LUT4 add_593_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2671), 
            .I3(n27681), .O(n2681[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_16 (.CI(n27681), .I0(encoder1_position[14]), .I1(n2671), 
            .CO(n27682));
    SB_LUT4 add_593_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2671), 
            .I3(n27680), .O(n2681[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_15 (.CI(n27680), .I0(encoder1_position[13]), .I1(n2671), 
            .CO(n27681));
    SB_LUT4 add_593_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2671), 
            .I3(n27679), .O(n2681[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_14 (.CI(n27679), .I0(encoder1_position[12]), .I1(n2671), 
            .CO(n27680));
    SB_LUT4 add_593_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2671), 
            .I3(n27678), .O(n2681[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_13 (.CI(n27678), .I0(encoder1_position[11]), .I1(n2671), 
            .CO(n27679));
    SB_LUT4 add_593_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2671), 
            .I3(n27677), .O(n2681[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_12 (.CI(n27677), .I0(encoder1_position[10]), .I1(n2671), 
            .CO(n27678));
    SB_LUT4 add_593_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2671), 
            .I3(n27676), .O(n2681[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_11 (.CI(n27676), .I0(encoder1_position[9]), .I1(n2671), 
            .CO(n27677));
    SB_LUT4 add_593_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2671), 
            .I3(n27675), .O(n2681[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_10 (.CI(n27675), .I0(encoder1_position[8]), .I1(n2671), 
            .CO(n27676));
    SB_LUT4 add_593_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2671), 
            .I3(n27674), .O(n2681[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_9 (.CI(n27674), .I0(encoder1_position[7]), .I1(n2671), 
            .CO(n27675));
    SB_LUT4 add_593_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2671), 
            .I3(n27673), .O(n2681[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_8 (.CI(n27673), .I0(encoder1_position[6]), .I1(n2671), 
            .CO(n27674));
    SB_LUT4 add_593_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2671), 
            .I3(n27672), .O(n2681[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_7 (.CI(n27672), .I0(encoder1_position[5]), .I1(n2671), 
            .CO(n27673));
    SB_LUT4 add_593_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2671), 
            .I3(n27671), .O(n2681[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_6 (.CI(n27671), .I0(encoder1_position[4]), .I1(n2671), 
            .CO(n27672));
    SB_LUT4 add_593_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2671), 
            .I3(n27670), .O(n2681[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_5 (.CI(n27670), .I0(encoder1_position[3]), .I1(n2671), 
            .CO(n27671));
    SB_LUT4 add_593_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2671), 
            .I3(n27669), .O(n2681[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_4 (.CI(n27669), .I0(encoder1_position[2]), .I1(n2671), 
            .CO(n27670));
    SB_LUT4 add_593_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2671), 
            .I3(n27668), .O(n2681[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_3 (.CI(n27668), .I0(encoder1_position[1]), .I1(n2671), 
            .CO(n27669));
    SB_LUT4 add_593_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n27667), .O(n2681[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_593_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_593_2 (.CI(n27667), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n27668));
    SB_CARRY add_593_1 (.CI(GND_net), .I0(n2671), .I1(n2671), .CO(n27667));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i895_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2671));   // quad.v(37[5] 40[8])
    defparam i895_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n18510(n18510), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B}), .PIN_7_c_1(PIN_7_c_1), 
            .n34961(n34961), .GND_net(GND_net), .n17911(n17911)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n18510, data_o, clk32MHz, PIN_6_c_0, reg_B, 
            PIN_7_c_1, n34961, GND_net, n17911) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18510;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    output n34961;
    input GND_net;
    input n17911;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n2, cnt_next_2__N_3459;
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18510));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_6_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_7_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n34961));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34961), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22839_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22839_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1141__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17911));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1141__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1141__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3459));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22848_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22848_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22841_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22841_2_lut.LUT_INIT = 16'h6666;
    
endmodule
