// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jan 29 23:28:20 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(122[22:39])
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(123[21:45])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n17980, n6;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire sda_enable, scl, scl_enable;
    wire [22:0]pwm_setpoint_22__N_3;
    
    wire RX_N_2;
    wire [31:0]motor_state_23__N_74;
    wire [25:0]encoder0_position_scaled_23__N_26;
    wire [23:0]displacement_23__N_50;
    
    wire n26017;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n25899, n25898, n25897, n25896, n26016, n25895;
    wire [3:0]state_3__N_319;
    
    wire n5, n11, n7, n8, n13810, n21, n23, n25894, n2696, 
        n26015, n26014, n25592, n22903, n18102, n18101, n18100, 
        n18099, n18098, n18097, n18096, n18095, n18091, n18090, 
        n18089, n18088, n18087, n35036;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n25893, n25892, n20, n19, n16, n11_adj_4785, n9, n6_adj_4786, 
        n5_adj_4787, n4, n3, n4_adj_4788, n5_adj_4789, n6_adj_4790, 
        n7_adj_4791, n8_adj_4792, n9_adj_4793, n10, n11_adj_4794, 
        n12, n13, n14, n15, n16_adj_4795, n17, n18, n19_adj_4796, 
        n20_adj_4797, n21_adj_4798, n22, n23_adj_4799, n24, n25, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    
    wire n34768;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    
    wire n25891, n26013, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n519, n518, n517, n516, n515, n514, n513, n511, n510, 
        n509, n26012, n25591, n122, n123, n9711, n34, n31, n30, 
        n28, n22_adj_4800, n21_adj_4801, n25890, n17_adj_4802, n16_adj_4803, 
        n31208, n771, n31159, n31157, n31155, n16_adj_4804, n12_adj_4805, 
        n10_adj_4806, n8_adj_4807, n22885, n26011, n5_adj_4808, n26010, 
        n25889, n25888, n22925, n25590, n26009, n26008, n26007, 
        n25589, n22937, n26006, n25887, n25886, n25885, n26005, 
        n25588, n26160, n26159, n25884, n21943, n25883, n25882, 
        n26004, n26158, n25587, n26003, n26157, n26156, n26155, 
        n26002, n26001, n26000, n26154, n25586, n25999, n25998, 
        n25997, n26153, n25585, n25996, n22927, n25995, n26152, 
        n25994, n26151, n25993, n26150, n25992, n26149, n25991, 
        n26148, n25990, n26147, n25989, n25988, n25987, n26146, 
        n25986, n26145, n25985, n25984, n26144, n26143, n26142, 
        n25983, n25982, n25981, n25980, n25979, n26141, n25978, 
        n25977, n26140, n26139, n26138, n26137, n26136, n25976, 
        n25975, n25974, n26135, n26134, n25973, n25972, n25606, 
        n25605, n26133, n25971, n26132, n25654, n26131, n26130, 
        n25970, n25969, n25968, n25604, n26129, n26128, n22757, 
        n26127, n25653, n26126, n26125, n25603, n25652, n26124, 
        n25651, n26123, n25855, n26122, n8_adj_4809, n26121, n26120, 
        n26119, n25854, n26118, n26117, n26116, n25602, n25650, 
        n25853, n16621, n21898, n26115, n26114, n26113, n26112, 
        n35882, n25649, n25601, n22743, n25852, n26111, n25851, 
        n25600, n25648, n25850, n26110, n26109, n26108, n26107, 
        n25849, n23001, n26106, n26105, n25848, n25593, n25647, 
        n26104, n25599, n26103, n25597, n25598, n25958, n25847, 
        n25957, n25646, n25645, n25956, n25596, n25846, n6_adj_4810, 
        n25595, n25845, n35879, n25644, n25643, n25844, n26102, 
        n21828, n21826, n26101, n25955, n25954, n25843, n16614, 
        n26100, n26099, n25842, n25953, n16613, n26098, n3303;
    wire [31:0]\FRAME_MATCHER.state_31__N_2579 ;
    
    wire n25841, n25840, n26097, n25839, n25952, n26096, n26095, 
        n26094, n25594, n25951, n26093, n26092, n26091, n25838, 
        n26090, n26089, n25837, n26088, n26087, n26086, n25836, 
        n25950, n26085, n25835, n25834, n25833, n25949, n26084, 
        n26083, n26082, n32929, n32812, n25948, n25947, n32337, 
        n25946, n25945, n25944, n26081, n26080, n23011, n23007, 
        n25943, n22919, n22893, n26079, n26078, n25942, n25941, 
        n25940, n22989, n26077, n25939, n4452, n25938, n26076, 
        n25937, n25936, n26075, n25935, n25934, n26074, n26073, 
        n25933, n26072, n26071, n26070, n25553, n25932, n26069, 
        n25931, n25930, n26068, n26067, n26066, n25929, n25552, 
        n26065, n26064, n18086, n26063, n26062, n26061, n26060, 
        n26059, n26058, n26057, n14_adj_4811, n9_adj_4812, n25928, 
        n26056, n26055, n25927, n26054, n25926, n25925, n25924, 
        n26053, n26052, n26051, n25923, n25922, n26050, n26049, 
        n25921, n26048, n26047, n25551, n26046, n25920, n25550, 
        n26045, n25549, n30_adj_4813, n29, n26044, n28_adj_4814, 
        n27, n26043, n25548, n26042, n25919, n26041, n26040, n25918, 
        n26039, n26038, n22895, n22965, n26037, n18_adj_4815, n26036, 
        n22997, n26035, n25917, n26034, n25916, n26033, n25915, 
        n22209, n22915, n25914, n26032, n25913, n25912, n25911, 
        n3_adj_4816, n22_adj_4817, n20_adj_4818, n18_adj_4819, n14_adj_4820, 
        n13_adj_4821, n7_adj_4822, n4_adj_4823, n22632, n18575, n18574, 
        n18573, n18572, n18571, n18570, n18569, n18568, n18567, 
        n18566, n18565, n18564, n18563, n18562, n18561, n18560, 
        n18559, n18558, n18557, n18556, n18555, n18554, n18553, 
        n18552, n18551, n18550, n18549, n18548, n18547, n18546, 
        n18545, n18544, n18541, n18540, n18536, n18535, n18534, 
        n18533, n18532, n18531, n18530, n18529, n18528, n18527, 
        n18526, n18525, n18524, n18523, n18522, n18521, n18520, 
        n18519, n18518, n18517, n18516, n18515, n18514, n18513, 
        n18512, n18511, n18510, n18509, n18508, n18507, n18506, 
        n18505, n18504, n18503, n18502, n18501, n18500, n18499, 
        n18498, n18497, n18496, n18495, n18494, n18493, n18492, 
        n18491, n18490, n18489, n435, n434, n433, n425, n26, 
        n24_adj_4824, n22_adj_4825, n18_adj_4826, n18488, n18485, 
        n18484, n18483, n18482, n18481, n18480, n18479, n18478, 
        n18477, n18476, n18475, n18474, n18473, n18472, n18471, 
        n18470, n18469, n18468, n18467, n18466, n18465, n18464, 
        n18463, n18462, n18461, n18460, n18459, n18458, n18457, 
        n18456, n18455, n18454, n18453, n18452, n18451, n18450, 
        n18447, n18446, n18445, n18444, n18443, n18442, n18441, 
        n18440, n18439, n18438, n18437, n18436, n18435, n18434, 
        n18433, n18085, n18432, n18431, n10_adj_4827, n18430, n18429, 
        n18428, n18427, n18426, n18425, n18424, n2, n18423, n15_adj_4828, 
        n18422, n31225, n18421, n18420, n18419, n18418, n18417, 
        n18416, n18415, n18414, n18413, n18412, n18411, n18410, 
        n18409, n18408, n18407, n18406, n3_adj_4829, n18405, n18404, 
        n18403, n18402, n18401, n18400, n18399, n18398, n18397, 
        n18396, n18395, n18394, n18393, n18392, n18391, n18390, 
        n18389, n18388, n18387, n18386, n18385, n18384, n18383, 
        n5_adj_4830, n18382, n18381, n18380, n18379, n18378, n18377, 
        n18376, n18375, n18374, n18373, n18372, n18371, n18370, 
        n18369, n18368, n63, n18367, n18366, n18365, n18364, n18363, 
        n18362, n18361, n18360, n4_adj_4831, n18359, n18358, quadA_debounced, 
        quadB_debounced, n18357, n18356, n18355, n18354, n18353, 
        n18352, n18351, n18350, n18349, n18348, n10_adj_4832, quadA_debounced_adj_4833, 
        quadB_debounced_adj_4834, n18347, n18346, n18345, n18344, 
        n18343, n18342, n18341, n18340, n34773, n18339, n18338, 
        n18337, n18336, n15_adj_4835, n18335, n18334, n18333, n18332, 
        n18331, n18330, n18329, n18328, n18327, n18326, n18325, 
        n18324, n18323, n18322, n18317, n18316, n18315, n18314, 
        n18313, n18312, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n18311, n18_adj_4836, n18310, n18309, n18084, n7_adj_4837, 
        n18308, n18307, n18306, n18305, n18304, n18303, n18302, 
        n18083, n18301, n18300, n18299, n18298, n18297, n18296, 
        n18295, n18294, n18293, n18292, n18291, n18290;
    wire [2:0]r_SM_Main_adj_5007;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5009;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3404;
    
    wire n24_adj_4839, n18289, n18288, n18287, n18286, n18285, n18284, 
        n18283, n4_adj_4840, n18282, n18281, n18280, n18279, n18278, 
        n18277, n18276, n18275, n18274, n18273, n18272, n18271, 
        n18270;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17_adj_4841, n25_adj_4842, n22_adj_4843, n5019;
    wire [1:0]reg_B_adj_5018;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n4_adj_4846, n15_adj_4847, n34918;
    wire [7:0]state_adj_5030;   // verilog/i2c_controller.v(32[12:17])
    
    wire n13_adj_4848, n12_adj_4849;
    wire [7:0]state_7__N_3815;
    
    wire n18082, n34852, n34922, n18081, n4604, n34871;
    wire [7:0]state_7__N_3831;
    
    wire n7_adj_4850, n34851, n4922, n34775, n18080, n18079, n18078, 
        n18077, n18076, n18075, n18074, n18073, n34753, n34747, 
        n34745, n18230, n18229, n18228, n18227, n18226, n18225, 
        n18224, n18223, n5276, n5273, n32360, n7_adj_4851, n8_adj_4852, 
        n9_adj_4853, n10_adj_4854, n11_adj_4855, n12_adj_4856, n13_adj_4857, 
        n14_adj_4858, n15_adj_4859, n16_adj_4860, n17_adj_4861, n18_adj_4862, 
        n19_adj_4863, n20_adj_4864, n21_adj_4865, n22_adj_4866, n23_adj_4867, 
        n24_adj_4868, n25_adj_4869, n619, n33043, n12_adj_4870, n674, 
        n675, n676, n677, n678, n679, n700, n728, n729, n730, 
        n731, n732, n733, n752, n753, n754, n755, n756, n757, 
        n758, n35048, n778, n5277, n5275, n806, n807, n808, 
        n809, n810, n811, n812, n8_adj_4871, n830, n831, n832, 
        n833, n834, n835, n836, n837, n856, n7_adj_4872, n883, 
        n884, n885, n886, n887, n888, n889, n890, n891, n908, 
        n909, n910, n911, n912, n913, n914, n915, n916, n922, 
        n923, n924, n925, n926, n927, n928, n929, n930, n931, 
        n25910, n934, n961, n962, n963, n964, n965, n966, n967, 
        n968, n969, n970, n986, n987, n988, n989, n990, n991, 
        n992, n993, n994, n995, n1012, n1039, n1040, n1041, 
        n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
        n1072, n1073, n1074, n1090, n1117, n1118, n1119, n1120, 
        n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
        n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
        n1150, n1151, n1152, n1153, n1168, n31767, n1195, n1196, 
        n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
        n1205, n1206, n1207, n1220, n1221, n1222, n1223, n1224, 
        n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
        n1246, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1298, 
        n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
        n1307, n1308, n1309, n1310, n1311, n1324, n1351, n1352, 
        n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
        n1361, n1362, n1363, n1364, n1365, n1376, n1377, n1378, 
        n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
        n1387, n1388, n1389, n1390, n1402, n1429, n1430, n1431, 
        n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
        n1440, n1441, n1442, n1443, n1444, n1454, n1455, n1456, 
        n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
        n1465, n1466, n1467, n1468, n1469, n1480, n1507, n1508, 
        n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
        n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1532, 
        n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
        n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
        n1558, n1585, n1586, n1587, n1588, n1589, n1590, n1591, 
        n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
        n1600, n1601, n1602, n1610, n1611, n1612, n1613, n1614, 
        n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n28827, n1636, n1663, 
        n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, 
        n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
        n1680, n1681, n1688, n1689, n1690, n1691, n1692, n1693, 
        n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, 
        n1702, n1703, n1704, n1705, n1706, n1714, n1741, n1742, 
        n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
        n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
        n1759, n1760, n1766, n1767, n1768, n1769, n1770, n1771, 
        n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
        n1780, n1781, n1782, n1783, n1784, n1785, n1792, n1819, 
        n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, 
        n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
        n1836, n1837, n1838, n1839, n1844, n1845, n1846, n1847, 
        n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
        n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
        n1864, n1870, n1897, n1898, n1899, n1900, n1901, n1902, 
        n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
        n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
        n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
        n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
        n1938, n1939, n1940, n1941, n1942, n1943, n1948, n30475, 
        n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
        n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
        n1991, n1992, n1993, n1994, n1995, n1996, n1997, n2000, 
        n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
        n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
        n2017, n2018, n2019, n2020, n2021, n2022, n2026, n2053, 
        n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, 
        n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
        n2070, n2071, n2073, n2076, n5522, n5521, n5520, n5519, 
        n5518, n5517, n5516, n5515, n5514, n5513, n5512, n5511, 
        n5510, n5509, n5508, n5507, n5506, n5505, n5504, n5502, 
        n5501, n16458, n17982, n17831, n17825, n17813, n33025, 
        n63_adj_4873, n29331, n18072, n18071, n18070, n26031, n18069, 
        n18068, n18067, n16606, n18066, n18065, n18064, n32040, 
        n34666, n4_adj_4874, n6_adj_4875, n7_adj_4876, n8_adj_4877, 
        n9_adj_4878, n10_adj_4879, n11_adj_4880, n12_adj_4881, n13_adj_4882, 
        n15_adj_4883, n17_adj_4884, n19_adj_4885, n21_adj_4886, n34774, 
        n23_adj_4887, n25_adj_4888, n27_adj_4889, n34772, n29_adj_4890, 
        n30_adj_4891, n31_adj_4892, n33, n35, n29947, n30466, n19_adj_4893, 
        n28_adj_4894, n34434, n34424, n27_adj_4895, n26_adj_4896, 
        n25_adj_4897, n5_adj_4898, n30471, n18166, n18165, n18164, 
        n18163, n18162, n18161, n18160, n18159, n18060, n18059, 
        n18058, n18057, n18055, n18052, n18051, n18050, n18049, 
        n18048, n18047, n26460, n16544, n26459, n26458, n26457, 
        n26456, n26455, n5278, n2_adj_4899, n3_adj_4900, n4_adj_4901, 
        n5_adj_4902, n6_adj_4903, n7_adj_4904, n8_adj_4905, n9_adj_4906, 
        n10_adj_4907, n11_adj_4908, n12_adj_4909, n13_adj_4910, n14_adj_4911, 
        n15_adj_4912, n16_adj_4913, n17_adj_4914, n18_adj_4915, n19_adj_4916, 
        n20_adj_4917, n21_adj_4918, n22_adj_4919, n23_adj_4920, n24_adj_4921, 
        n25_adj_4922, n26454, n26453, n26452, n26451, n26450, n26449, 
        n26448, n26447, n26446, n26445, n26444, n26443, n26442, 
        n26441, n26440, n26439, n26438, n34142, n26437, n34136, 
        n34134, n34130, n34127, n34710, n36350, n35944, n13_adj_4923, 
        n23_adj_4924, n27_adj_4925, n29_adj_4926, n37, n39, n43, 
        n45, n34622, n49, n9799, n34624, n4_adj_4927, n6_adj_4928, 
        n24_adj_4929, n21_adj_4930, n20_adj_4931, n5_adj_4932, n17_adj_4933, 
        n26030, n25909, n31153, n14_adj_4934, n10_adj_4935, n22933, 
        n34061, n18046, n18045, n34058, n20_adj_4936, n18_adj_4937, 
        n16_adj_4938, n18044, n34923, n30480, n34037, n34036, n26029, 
        n26028, n34_adj_4939, n33_adj_4940, n32, n31_adj_4941, n30_adj_4942, 
        n28_adj_4943, n26_adj_4944, n24_adj_4945, n19_adj_4946, n16_adj_4947, 
        n18043, n18042, n18040, n37_adj_4948, n36, n30_adj_4949, 
        n32962, n29_adj_4950, n28_adj_4951, n27_adj_4952, n26_adj_4953, 
        n25_adj_4954, n24_adj_4955, n23_adj_4956, n22_adj_4957, n21_adj_4958, 
        n26027, n4_adj_4959, n35425, n32355, n34921, n16549, n16456, 
        n31986, n33075, n13933, n32238, n26026, n25908, n25907, 
        n26025, n33995, n26024, n25906, n25905, n26023, n25904, 
        n25903, n26022, n25902, n25901, n26021, n26020, n26019, 
        n26018, n33988, n6_adj_4960, n25900, n32029;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced, 
            quadB_debounced}), .VCC_net(VCC_net), .reg_B({reg_B}), .n32962(n32962), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n18541(n18541), .n18057(n18057), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_LUT4 i13911_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18491));   // verilog/coms.v(127[12] 300[6])
    defparam i13911_3_lut.LUT_INIT = 16'hcaca;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13912_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18492));   // verilog/coms.v(127[12] 300[6])
    defparam i13912_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h3_38 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_50[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF h2_37 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(state_7__N_3831[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.GND_net(GND_net), .clk32MHz(clk32MHz), .\state[1] (state[1]), 
            .n29331(n29331), .n17813(n17813), .n31208(n31208), .VCC_net(VCC_net), 
            .timer({timer}), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .neopxl_color({neopxl_color}), .LED_c(LED_c), .\state_3__N_319[1] (state_3__N_319[1]), 
            .n18064(n18064), .n18060(n18060), .n18575(n18575), .n18574(n18574), 
            .n18573(n18573), .n18572(n18572), .n18571(n18571), .n18570(n18570), 
            .n18569(n18569), .n18568(n18568), .n18567(n18567), .n18566(n18566), 
            .n18565(n18565), .n18564(n18564), .n18563(n18563), .n18562(n18562), 
            .n18561(n18561), .n18560(n18560), .n18559(n18559), .n18558(n18558), 
            .n18557(n18557), .n18556(n18556), .n18555(n18555), .n18554(n18554), 
            .n18553(n18553), .n18552(n18552), .n18551(n18551), .n18550(n18550), 
            .n18549(n18549), .n18548(n18548), .n18547(n18547), .n18546(n18546), 
            .n18545(n18545), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[10] 49[2])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13913_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18493));   // verilog/coms.v(127[12] 300[6])
    defparam i13913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13914_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18494));   // verilog/coms.v(127[12] 300[6])
    defparam i13914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13915_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18495));   // verilog/coms.v(127[12] 300[6])
    defparam i13915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13916_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18496));   // verilog/coms.v(127[12] 300[6])
    defparam i13916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13917_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18497));   // verilog/coms.v(127[12] 300[6])
    defparam i13917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13918_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18498));   // verilog/coms.v(127[12] 300[6])
    defparam i13918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13919_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18499));   // verilog/coms.v(127[12] 300[6])
    defparam i13919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13920_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18500));   // verilog/coms.v(127[12] 300[6])
    defparam i13920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13921_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18501));   // verilog/coms.v(127[12] 300[6])
    defparam i13921_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dir_42 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i13922_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18502));   // verilog/coms.v(127[12] 300[6])
    defparam i13922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13923_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18503));   // verilog/coms.v(127[12] 300[6])
    defparam i13923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13924_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18504));   // verilog/coms.v(127[12] 300[6])
    defparam i13924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13925_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18505));   // verilog/coms.v(127[12] 300[6])
    defparam i13925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13926_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18506));   // verilog/coms.v(127[12] 300[6])
    defparam i13926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13927_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18507));   // verilog/coms.v(127[12] 300[6])
    defparam i13927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13928_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18508));   // verilog/coms.v(127[12] 300[6])
    defparam i13928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13929_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18509));   // verilog/coms.v(127[12] 300[6])
    defparam i13929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13930_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18510));   // verilog/coms.v(127[12] 300[6])
    defparam i13930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13931_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18511));   // verilog/coms.v(127[12] 300[6])
    defparam i13931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13932_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18512));   // verilog/coms.v(127[12] 300[6])
    defparam i13932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13933_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18513));   // verilog/coms.v(127[12] 300[6])
    defparam i13933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13934_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18514));   // verilog/coms.v(127[12] 300[6])
    defparam i13934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13935_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18515));   // verilog/coms.v(127[12] 300[6])
    defparam i13935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13936_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18516));   // verilog/coms.v(127[12] 300[6])
    defparam i13936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13937_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18517));   // verilog/coms.v(127[12] 300[6])
    defparam i13937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13938_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18518));   // verilog/coms.v(127[12] 300[6])
    defparam i13938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13939_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18519));   // verilog/coms.v(127[12] 300[6])
    defparam i13939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13940_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18520));   // verilog/coms.v(127[12] 300[6])
    defparam i13940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13941_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18521));   // verilog/coms.v(127[12] 300[6])
    defparam i13941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13942_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18522));   // verilog/coms.v(127[12] 300[6])
    defparam i13942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13943_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18523));   // verilog/coms.v(127[12] 300[6])
    defparam i13943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13944_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18524));   // verilog/coms.v(127[12] 300[6])
    defparam i13944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13945_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18525));   // verilog/coms.v(127[12] 300[6])
    defparam i13945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13946_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18526));   // verilog/coms.v(127[12] 300[6])
    defparam i13946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13947_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18527));   // verilog/coms.v(127[12] 300[6])
    defparam i13947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13948_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18528));   // verilog/coms.v(127[12] 300[6])
    defparam i13948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13949_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18529));   // verilog/coms.v(127[12] 300[6])
    defparam i13949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13950_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18530));   // verilog/coms.v(127[12] 300[6])
    defparam i13950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13951_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18531));   // verilog/coms.v(127[12] 300[6])
    defparam i13951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13952_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18532));   // verilog/coms.v(127[12] 300[6])
    defparam i13952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13953_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18533));   // verilog/coms.v(127[12] 300[6])
    defparam i13953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13954_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18534));   // verilog/coms.v(127[12] 300[6])
    defparam i13954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13955_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18535));   // verilog/coms.v(127[12] 300[6])
    defparam i13955_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13956_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18536));   // verilog/coms.v(127[12] 300[6])
    defparam i13956_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13960_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4), .I3(n16549), 
            .O(n18540));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13960_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13961_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n32962), 
            .I3(GND_net), .O(n18541));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut (.I0(n34058), .I1(state_adj_5030[2]), .I2(n4604), 
            .I3(n11), .O(n5_adj_4808));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13_4_lut.LUT_INIT = 16'h5cfc;
    SB_LUT4 i13964_3_lut (.I0(quadA_debounced_adj_4833), .I1(reg_B_adj_5018[1]), 
            .I2(n33025), .I3(GND_net), .O(n18544));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13965_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n29331), .I3(GND_net), .O(n18545));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13966_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n29331), .I3(GND_net), .O(n18546));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13967_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n29331), .I3(GND_net), .O(n18547));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13968_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n29331), .I3(GND_net), .O(n18548));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13969_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n29331), .I3(GND_net), .O(n18549));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13970_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n29331), .I3(GND_net), .O(n18550));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13971_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n29331), .I3(GND_net), .O(n18551));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13972_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n29331), .I3(GND_net), .O(n18552));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13973_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n29331), .I3(GND_net), .O(n18553));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13974_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n29331), .I3(GND_net), .O(n18554));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13975_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n29331), .I3(GND_net), .O(n18555));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13976_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n29331), .I3(GND_net), .O(n18556));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13977_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n29331), .I3(GND_net), .O(n18557));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13978_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n29331), .I3(GND_net), .O(n18558));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i409_3_lut_4_lut (.I0(n2), .I1(encoder0_position[23]), 
            .I2(n619), .I3(n5273), .O(n674));
    defparam encoder0_position_23__I_0_i409_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 i13979_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n29331), .I3(GND_net), .O(n18559));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13980_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n29331), .I3(GND_net), .O(n18560));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13981_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n29331), .I3(GND_net), .O(n18561));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13982_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n29331), .I3(GND_net), .O(n18562));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13983_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n29331), .I3(GND_net), .O(n18563));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13984_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n29331), .I3(GND_net), .O(n18564));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13985_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n29331), .I3(GND_net), .O(n18565));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13986_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n29331), .I3(GND_net), .O(n18566));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13987_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n29331), .I3(GND_net), .O(n18567));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13988_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n29331), .I3(GND_net), .O(n18568));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13989_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n29331), .I3(GND_net), .O(n18569));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13990_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n29331), .I3(GND_net), .O(n18570));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13991_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n29331), .I3(GND_net), .O(n18571));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13992_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n29331), .I3(GND_net), .O(n18572));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13993_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n29331), .I3(GND_net), .O(n18573));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13994_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n29331), .I3(GND_net), .O(n18574));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13995_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n29331), .I3(GND_net), .O(n18575));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_3_lut (.I0(duty[1]), .I1(n35425), .I2(n24), .I3(n25585), 
            .O(pwm_setpoint_22__N_3[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13908_3_lut (.I0(n17980), .I1(r_Bit_Index[0]), .I2(n17825), 
            .I3(GND_net), .O(n18488));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13908_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 mux_59_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4799));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25007_3_lut_4_lut (.I0(n3_adj_4829), .I1(n4_adj_4927), .I2(n5275), 
            .I3(n4_adj_4831), .O(n31159));
    defparam i25007_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13742_3_lut (.I0(n17982), .I1(r_Bit_Index_adj_5009[0]), .I2(n17831), 
            .I3(GND_net), .O(n18322));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13742_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4798));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13479_3_lut (.I0(quadB_debounced_adj_4834), .I1(reg_B_adj_5018[0]), 
            .I2(n33025), .I3(GND_net), .O(n18059));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i25001_3_lut_4_lut (.I0(n3_adj_4829), .I1(n4_adj_4927), .I2(n5278), 
            .I3(n7), .O(n31153));
    defparam i25001_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13480_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n29331), .I3(GND_net), .O(n18060));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13480_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n5_adj_4898), .I1(n122), .I2(n2696), .I3(n63_adj_4873), 
            .O(n6_adj_4928));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i3_4_lut (.I0(n36350), .I1(n6_adj_4928), .I2(n16621), .I3(n4452), 
            .O(n8_adj_4809));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hcfce;
    SB_LUT4 i4_4_lut (.I0(n122), .I1(n8_adj_4809), .I2(n63), .I3(n5_adj_4932), 
            .O(n35882));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 i25003_3_lut_4_lut (.I0(n3_adj_4829), .I1(n4_adj_4927), .I2(n5277), 
            .I3(n6), .O(n31155));
    defparam i25003_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1628 (.I0(n19_adj_4893), .I1(n2696), .I2(n16621), 
            .I3(n4452), .O(n30480));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1628.LUT_INIT = 16'heeef;
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n30480), .I2(n63_adj_4873), .I3(GND_net), 
            .O(n7_adj_4822));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_LUT4 i2_4_lut (.I0(n7_adj_4822), .I1(n123), .I2(n16613), .I3(n9711), 
            .O(n6_adj_4810));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'haeaf;
    SB_LUT4 i3_4_lut_adj_1629 (.I0(n63), .I1(n6_adj_4810), .I2(n16606), 
            .I3(\FRAME_MATCHER.state_31__N_2579 [1]), .O(n35879));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1629.LUT_INIT = 16'hdfdd;
    SB_LUT4 i25005_3_lut_4_lut (.I0(n3_adj_4829), .I1(n4_adj_4927), .I2(n5276), 
            .I3(n5), .O(n31157));
    defparam i25005_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i28890_2_lut_3_lut (.I0(n3_adj_4829), .I1(n4_adj_4927), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n619));
    defparam i28890_2_lut_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 i13484_4_lut (.I0(n31208), .I1(state[1]), .I2(state_3__N_319[1]), 
            .I3(n17813), .O(n18064));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13484_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i13485_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18065));   // verilog/coms.v(127[12] 300[6])
    defparam i13485_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13486_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18066));   // verilog/coms.v(127[12] 300[6])
    defparam i13486_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13487_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18067));   // verilog/coms.v(127[12] 300[6])
    defparam i13487_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13488_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18068));   // verilog/coms.v(127[12] 300[6])
    defparam i13488_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13489_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18069));   // verilog/coms.v(127[12] 300[6])
    defparam i13489_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13490_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18070));   // verilog/coms.v(127[12] 300[6])
    defparam i13490_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13491_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18071));   // verilog/coms.v(127[12] 300[6])
    defparam i13491_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13492_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18072));   // verilog/coms.v(127[12] 300[6])
    defparam i13492_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13493_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18073));   // verilog/coms.v(127[12] 300[6])
    defparam i13493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13494_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18074));   // verilog/coms.v(127[12] 300[6])
    defparam i13494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13495_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18075));   // verilog/coms.v(127[12] 300[6])
    defparam i13495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13496_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18076));   // verilog/coms.v(127[12] 300[6])
    defparam i13496_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13497_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18077));   // verilog/coms.v(127[12] 300[6])
    defparam i13497_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13498_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18078));   // verilog/coms.v(127[12] 300[6])
    defparam i13498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13499_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18079));   // verilog/coms.v(127[12] 300[6])
    defparam i13499_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13500_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18080));   // verilog/coms.v(127[12] 300[6])
    defparam i13500_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13501_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18081));   // verilog/coms.v(127[12] 300[6])
    defparam i13501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13502_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18082));   // verilog/coms.v(127[12] 300[6])
    defparam i13502_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13503_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18083));   // verilog/coms.v(127[12] 300[6])
    defparam i13503_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13504_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18084));   // verilog/coms.v(127[12] 300[6])
    defparam i13504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13505_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n32040), .I3(GND_net), .O(n18085));   // verilog/coms.v(127[12] 300[6])
    defparam i13505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13506_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n32040), .I3(GND_net), .O(n18086));   // verilog/coms.v(127[12] 300[6])
    defparam i13506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13507_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n32040), .I3(GND_net), .O(n18087));   // verilog/coms.v(127[12] 300[6])
    defparam i13507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13508_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n32040), .I3(GND_net), .O(n18088));   // verilog/coms.v(127[12] 300[6])
    defparam i13508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13509_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n32040), .I3(GND_net), .O(n18089));   // verilog/coms.v(127[12] 300[6])
    defparam i13509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13510_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n32040), .I3(GND_net), .O(n18090));   // verilog/coms.v(127[12] 300[6])
    defparam i13510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13511_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n32040), .I3(GND_net), .O(n18091));   // verilog/coms.v(127[12] 300[6])
    defparam i13511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13515_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n30475), .I3(GND_net), .O(n18095));   // verilog/coms.v(127[12] 300[6])
    defparam i13515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13516_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n30475), .I3(GND_net), .O(n18096));   // verilog/coms.v(127[12] 300[6])
    defparam i13516_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1733_2 (.CI(VCC_net), .I0(n514), .I1(GND_net), .CO(n25650));
    SB_LUT4 encoder0_position_23__I_0_add_460_8_lut (.I0(n35048), .I1(n674), 
            .I2(VCC_net), .I3(n25553), .O(n752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_513_9_lut (.I0(n35036), .I1(n752), 
            .I2(VCC_net), .I3(n25649), .O(n830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_460_7_lut (.I0(GND_net), .I1(n675), 
            .I2(GND_net), .I3(n25552), .O(n728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_513_8_lut (.I0(GND_net), .I1(n753), 
            .I2(VCC_net), .I3(n25648), .O(n806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_3 (.CI(n25585), .I0(n35425), .I1(n24), .CO(n25586));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i13517_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n30475), .I3(GND_net), .O(n18097));   // verilog/coms.v(127[12] 300[6])
    defparam i13517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_2_lut (.I0(duty[0]), .I1(n35425), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_3[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4797));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF h1_36 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_CARRY encoder0_position_23__I_0_add_513_8 (.CI(n25648), .I0(n753), 
            .I1(VCC_net), .CO(n25649));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 LessThan_687_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4878));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4796));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_513_7_lut (.I0(GND_net), .I1(n754), 
            .I2(GND_net), .I3(n25647), .O(n807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_7 (.CI(n25647), .I0(n754), 
            .I1(GND_net), .CO(n25648));
    SB_CARRY add_615_2 (.CI(VCC_net), .I0(n35425), .I1(n25), .CO(n25585));
    SB_LUT4 mux_59_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_687_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4880));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4884));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4889));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4883));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_23__I_0_add_513_6_lut (.I0(GND_net), .I1(n755), 
            .I2(GND_net), .I3(n25646), .O(n808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_6 (.CI(n25646), .I0(n755), 
            .I1(GND_net), .CO(n25647));
    SB_LUT4 encoder0_position_23__I_0_add_513_5_lut (.I0(GND_net), .I1(n756), 
            .I2(VCC_net), .I3(n25645), .O(n809)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_687_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4882));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4876));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_59_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_687_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4886));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4887));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4885));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4890));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4892));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_59_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_687_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4888));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_687_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_59_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_513_5 (.CI(n25645), .I0(n756), 
            .I1(VCC_net), .CO(n25646));
    SB_CARRY encoder0_position_23__I_0_add_460_7 (.CI(n25552), .I0(n675), 
            .I1(GND_net), .CO(n25553));
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_460_6_lut (.I0(GND_net), .I1(n676), 
            .I2(GND_net), .I3(n25551), .O(n729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_59_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_513_4_lut (.I0(GND_net), .I1(n757), 
            .I2(GND_net), .I3(n25644), .O(n810)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4869));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4868));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4867));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_460_6 (.CI(n25551), .I0(n676), 
            .I1(GND_net), .CO(n25552));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4866));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4865));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_513_4 (.CI(n25644), .I0(n757), 
            .I1(GND_net), .CO(n25645));
    SB_LUT4 encoder0_position_23__I_0_add_460_5_lut (.I0(GND_net), .I1(n677), 
            .I2(VCC_net), .I3(n25550), .O(n730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4864));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4863));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4862));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_513_3_lut (.I0(GND_net), .I1(n758), 
            .I2(VCC_net), .I3(n25643), .O(n811)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_5 (.CI(n25550), .I0(n677), 
            .I1(VCC_net), .CO(n25551));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4861));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4860));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4859));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_513_3 (.CI(n25643), .I0(n758), 
            .I1(VCC_net), .CO(n25644));
    SB_LUT4 mux_59_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_460_4_lut (.I0(GND_net), .I1(n678), 
            .I2(GND_net), .I3(n25549), .O(n731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_513_2_lut (.I0(GND_net), .I1(n516), 
            .I2(GND_net), .I3(VCC_net), .O(n812)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_2_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_23__I_0_add_460_4 (.CI(n25549), .I0(n678), 
            .I1(GND_net), .CO(n25550));
    SB_CARRY encoder0_position_23__I_0_add_513_2 (.CI(VCC_net), .I0(n516), 
            .I1(GND_net), .CO(n25643));
    SB_LUT4 encoder0_position_23__I_0_add_460_3_lut (.I0(GND_net), .I1(n679), 
            .I2(VCC_net), .I3(n25548), .O(n732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_460_3 (.CI(n25548), .I0(n679), 
            .I1(VCC_net), .CO(n25549));
    SB_LUT4 encoder0_position_23__I_0_add_460_2_lut (.I0(GND_net), .I1(n515), 
            .I2(GND_net), .I3(VCC_net), .O(n733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_2 (.CI(VCC_net), .I0(n515), 
            .I1(GND_net), .CO(n25548));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4858));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4857));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4856));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4795));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_59_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_59_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4855));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4854));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4853));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_615_24_lut (.I0(duty[22]), .I1(n35425), .I2(n3), .I3(n25606), 
            .O(pwm_setpoint_22__N_3[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_24_lut.LUT_INIT = 16'h8BB8;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4852));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4851));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_615_23_lut (.I0(duty[21]), .I1(n35425), .I2(n4_adj_4788), 
            .I3(n25605), .O(pwm_setpoint_22__N_3[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_59_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_615_23 (.CI(n25605), .I0(n35425), .I1(n4_adj_4788), .CO(n25606));
    SB_LUT4 add_615_22_lut (.I0(duty[20]), .I1(n35425), .I2(n5_adj_4789), 
            .I3(n25604), .O(pwm_setpoint_22__N_3[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_615_22 (.CI(n25604), .I0(n35425), .I1(n5_adj_4789), .CO(n25605));
    SB_LUT4 add_615_21_lut (.I0(duty[19]), .I1(n35425), .I2(n6_adj_4790), 
            .I3(n25603), .O(pwm_setpoint_22__N_3[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_615_21 (.CI(n25603), .I0(n35425), .I1(n6_adj_4790), .CO(n25604));
    SB_LUT4 encoder0_position_23__I_0_add_1361_26_lut (.I0(GND_net), .I1(n2000), 
            .I2(VCC_net), .I3(n26160), .O(n2053)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_25_lut (.I0(GND_net), .I1(n2001), 
            .I2(VCC_net), .I3(n26159), .O(n2054)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_25 (.CI(n26159), .I0(n2001), 
            .I1(VCC_net), .CO(n26160));
    SB_LUT4 encoder0_position_23__I_0_add_1361_24_lut (.I0(GND_net), .I1(n2002), 
            .I2(VCC_net), .I3(n26158), .O(n2055)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_24 (.CI(n26158), .I0(n2002), 
            .I1(VCC_net), .CO(n26159));
    SB_LUT4 encoder0_position_23__I_0_add_1361_23_lut (.I0(GND_net), .I1(n2003), 
            .I2(VCC_net), .I3(n26157), .O(n2056)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_50[23]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_50[22]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_CARRY encoder0_position_23__I_0_add_1361_23 (.CI(n26157), .I0(n2003), 
            .I1(VCC_net), .CO(n26158));
    SB_LUT4 encoder0_position_23__I_0_add_1361_22_lut (.I0(GND_net), .I1(n2004), 
            .I2(VCC_net), .I3(n26156), .O(n2057)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_22 (.CI(n26156), .I0(n2004), 
            .I1(VCC_net), .CO(n26157));
    SB_LUT4 encoder0_position_23__I_0_add_1361_21_lut (.I0(GND_net), .I1(n2005), 
            .I2(VCC_net), .I3(n26155), .O(n2058)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_21 (.CI(n26155), .I0(n2005), 
            .I1(VCC_net), .CO(n26156));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1361_20_lut (.I0(GND_net), .I1(n2006), 
            .I2(VCC_net), .I3(n26154), .O(n2059)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_20 (.CI(n26154), .I0(n2006), 
            .I1(VCC_net), .CO(n26155));
    SB_LUT4 encoder0_position_23__I_0_add_1361_19_lut (.I0(GND_net), .I1(n2007), 
            .I2(VCC_net), .I3(n26153), .O(n2060)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_19 (.CI(n26153), .I0(n2007), 
            .I1(VCC_net), .CO(n26154));
    SB_LUT4 encoder0_position_23__I_0_add_1361_18_lut (.I0(GND_net), .I1(n2008), 
            .I2(VCC_net), .I3(n26152), .O(n2061)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_18 (.CI(n26152), .I0(n2008), 
            .I1(VCC_net), .CO(n26153));
    SB_LUT4 encoder0_position_23__I_0_add_1361_17_lut (.I0(GND_net), .I1(n2009), 
            .I2(VCC_net), .I3(n26151), .O(n2062)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4921));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4920));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4919));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_17 (.CI(n26151), .I0(n2009), 
            .I1(VCC_net), .CO(n26152));
    SB_LUT4 add_615_20_lut (.I0(duty[18]), .I1(n35425), .I2(n7_adj_4791), 
            .I3(n25602), .O(pwm_setpoint_22__N_3[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4918));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1361_16_lut (.I0(GND_net), .I1(n2010), 
            .I2(VCC_net), .I3(n26150), .O(n2063)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_16 (.CI(n26150), .I0(n2010), 
            .I1(VCC_net), .CO(n26151));
    SB_LUT4 encoder0_position_23__I_0_add_1361_15_lut (.I0(GND_net), .I1(n2011), 
            .I2(VCC_net), .I3(n26149), .O(n2064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_15 (.CI(n26149), .I0(n2011), 
            .I1(VCC_net), .CO(n26150));
    SB_LUT4 encoder0_position_23__I_0_add_1361_14_lut (.I0(GND_net), .I1(n2012), 
            .I2(VCC_net), .I3(n26148), .O(n2065)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4917));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_14 (.CI(n26148), .I0(n2012), 
            .I1(VCC_net), .CO(n26149));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4916));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1361_13_lut (.I0(GND_net), .I1(n2013), 
            .I2(VCC_net), .I3(n26147), .O(n2066)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4915));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_13 (.CI(n26147), .I0(n2013), 
            .I1(VCC_net), .CO(n26148));
    SB_LUT4 encoder0_position_23__I_0_add_1361_12_lut (.I0(GND_net), .I1(n2014), 
            .I2(VCC_net), .I3(n26146), .O(n2067)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4914));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_12 (.CI(n26146), .I0(n2014), 
            .I1(VCC_net), .CO(n26147));
    SB_LUT4 encoder0_position_23__I_0_add_1361_11_lut (.I0(GND_net), .I1(n2015), 
            .I2(VCC_net), .I3(n26145), .O(n2068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_11 (.CI(n26145), .I0(n2015), 
            .I1(VCC_net), .CO(n26146));
    SB_LUT4 encoder0_position_23__I_0_add_1361_10_lut (.I0(GND_net), .I1(n2016), 
            .I2(VCC_net), .I3(n26144), .O(n2069)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_10 (.CI(n26144), .I0(n2016), 
            .I1(VCC_net), .CO(n26145));
    SB_LUT4 encoder0_position_23__I_0_add_1361_9_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n26143), .O(n2070)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_9 (.CI(n26143), .I0(n2017), 
            .I1(VCC_net), .CO(n26144));
    SB_LUT4 encoder0_position_23__I_0_add_1361_8_lut (.I0(GND_net), .I1(n2018), 
            .I2(GND_net), .I3(n26142), .O(n2071)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_8 (.CI(n26142), .I0(n2018), 
            .I1(GND_net), .CO(n26143));
    SB_LUT4 i13518_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n30475), .I3(GND_net), .O(n18098));   // verilog/coms.v(127[12] 300[6])
    defparam i13518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_7_lut (.I0(n2073), .I1(n2019), 
            .I2(GND_net), .I3(n26141), .O(n33995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_615_20 (.CI(n25602), .I0(n35425), .I1(n7_adj_4791), .CO(n25603));
    SB_CARRY encoder0_position_23__I_0_add_1361_7 (.CI(n26141), .I0(n2019), 
            .I1(GND_net), .CO(n26142));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4913));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1361_6_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n26140), .O(n2073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_19_lut (.I0(duty[17]), .I1(n35425), .I2(n8_adj_4792), 
            .I3(n25601), .O(pwm_setpoint_22__N_3[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_615_19 (.CI(n25601), .I0(n35425), .I1(n8_adj_4792), .CO(n25602));
    SB_CARRY encoder0_position_23__I_0_add_1361_6 (.CI(n26140), .I0(n2020), 
            .I1(VCC_net), .CO(n26141));
    SB_LUT4 encoder0_position_23__I_0_add_1361_5_lut (.I0(n6_adj_4960), .I1(n2021), 
            .I2(GND_net), .I3(n26139), .O(n34037)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_23__I_0_add_1361_5 (.CI(n26139), .I0(n2021), 
            .I1(GND_net), .CO(n26140));
    SB_LUT4 encoder0_position_23__I_0_add_1361_4_lut (.I0(n2076), .I1(n2022), 
            .I2(VCC_net), .I3(n26138), .O(n6_adj_4960)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_4 (.CI(n26138), .I0(n2022), 
            .I1(VCC_net), .CO(n26139));
    SB_LUT4 encoder0_position_23__I_0_add_1361_3_lut (.I0(GND_net), .I1(n931), 
            .I2(GND_net), .I3(n26137), .O(n2076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_3 (.CI(n26137), .I0(n931), 
            .I1(GND_net), .CO(n26138));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4912));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n26137));
    SB_LUT4 add_1777_23_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n26136), .O(n5501)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1777_22_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n26135), .O(n5502)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_22 (.CI(n26135), .I0(GND_net), .I1(VCC_net), .CO(n26136));
    SB_LUT4 add_615_18_lut (.I0(duty[16]), .I1(n35425), .I2(n9_adj_4793), 
            .I3(n25600), .O(pwm_setpoint_22__N_3[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1777_21_lut (.I0(encoder0_position[23]), .I1(GND_net), .I2(n619), 
            .I3(n26134), .O(encoder0_position_scaled_23__N_26[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1777_21 (.CI(n26134), .I0(GND_net), .I1(n619), .CO(n26135));
    SB_CARRY add_615_18 (.CI(n25600), .I0(n35425), .I1(n9_adj_4793), .CO(n25601));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4786));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1777_20_lut (.I0(GND_net), .I1(GND_net), .I2(n700), .I3(n26133), 
            .O(n5504)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4911));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1777_20 (.CI(n26133), .I0(GND_net), .I1(n700), .CO(n26134));
    SB_LUT4 add_1777_19_lut (.I0(GND_net), .I1(GND_net), .I2(n778), .I3(n26132), 
            .O(n5505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_17_lut (.I0(duty[15]), .I1(n35425), .I2(n10), .I3(n25599), 
            .O(pwm_setpoint_22__N_3[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1777_19 (.CI(n26132), .I0(GND_net), .I1(n778), .CO(n26133));
    SB_LUT4 i13519_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n30475), .I3(GND_net), .O(n18099));   // verilog/coms.v(127[12] 300[6])
    defparam i13519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4910));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4909));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4908));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4907));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_59_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_1777_18_lut (.I0(GND_net), .I1(GND_net), .I2(n856), .I3(n26131), 
            .O(n5506)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_18 (.CI(n26131), .I0(GND_net), .I1(n856), .CO(n26132));
    SB_LUT4 add_1777_17_lut (.I0(GND_net), .I1(GND_net), .I2(n934), .I3(n26130), 
            .O(n5507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_17 (.CI(n25599), .I0(n35425), .I1(n10), .CO(n25600));
    SB_CARRY add_1777_17 (.CI(n26130), .I0(GND_net), .I1(n934), .CO(n26131));
    SB_LUT4 add_1777_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1012), .I3(n26129), 
            .O(n5508)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_16 (.CI(n26129), .I0(GND_net), .I1(n1012), .CO(n26130));
    SB_LUT4 add_1777_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1090), .I3(n26128), 
            .O(n5509)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_16_lut (.I0(duty[14]), .I1(n35425), .I2(n11_adj_4794), 
            .I3(n25598), .O(pwm_setpoint_22__N_3[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_615_16 (.CI(n25598), .I0(n35425), .I1(n11_adj_4794), 
            .CO(n25599));
    SB_CARRY add_1777_15 (.CI(n26128), .I0(GND_net), .I1(n1090), .CO(n26129));
    SB_LUT4 add_1777_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1168), .I3(n26127), 
            .O(n5510)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4906));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4905));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4935));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4904));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4903));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[29]), .I2(pwm_counter[25]), 
            .I3(pwm_counter[26]), .O(n14_adj_4934));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[30]), .I1(n14_adj_4934), .I2(n10_adj_4935), 
            .I3(pwm_counter[24]), .O(n16456));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_1777_14 (.CI(n26127), .I0(GND_net), .I1(n1168), .CO(n26128));
    SB_LUT4 add_1777_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1246), .I3(n26126), 
            .O(n5511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_13 (.CI(n26126), .I0(GND_net), .I1(n1246), .CO(n26127));
    SB_LUT4 add_1777_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1324), .I3(n26125), 
            .O(n5512)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_15_lut (.I0(duty[13]), .I1(n35425), .I2(n12), .I3(n25597), 
            .O(pwm_setpoint_22__N_3[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1777_12 (.CI(n26125), .I0(GND_net), .I1(n1324), .CO(n26126));
    SB_LUT4 add_1777_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1402), .I3(n26124), 
            .O(n5513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_11 (.CI(n26124), .I0(GND_net), .I1(n1402), .CO(n26125));
    SB_CARRY add_615_15 (.CI(n25597), .I0(n35425), .I1(n12), .CO(n25598));
    SB_LUT4 add_1777_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1480), .I3(n26123), 
            .O(n5514)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3158_i20_3_lut (.I0(encoder0_position[19]), .I1(n6), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4902));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1777_10 (.CI(n26123), .I0(GND_net), .I1(n1480), .CO(n26124));
    SB_LUT4 add_1777_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1558), .I3(n26122), 
            .O(n5515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_9 (.CI(n26122), .I0(GND_net), .I1(n1558), .CO(n26123));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4901));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1777_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1636), .I3(n26121), 
            .O(n5516)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1494_3_lut (.I0(n2026), .I1(n5521), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[1]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1494_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4900));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3158_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n425));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1777_8 (.CI(n26121), .I0(GND_net), .I1(n1636), .CO(n26122));
    SB_LUT4 add_1777_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1714), .I3(n26120), 
            .O(n5517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_7 (.CI(n26120), .I0(GND_net), .I1(n1714), .CO(n26121));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4787));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1493_3_lut (.I0(n1948), .I1(n5520), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[2]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1493_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1492_3_lut (.I0(n1870), .I1(n5519), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[3]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1492_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1491_3_lut (.I0(n1792), .I1(n5518), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[4]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1491_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1490_3_lut (.I0(n1714), .I1(n5517), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[5]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1490_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1489_3_lut (.I0(n1636), .I1(n5516), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[6]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1489_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1488_3_lut (.I0(n1558), .I1(n5515), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[7]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1488_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1487_3_lut (.I0(n1480), .I1(n5514), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[8]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1487_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1486_3_lut (.I0(n1402), .I1(n5513), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[9]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1486_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1485_3_lut (.I0(n1324), .I1(n5512), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[10]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1485_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_1777_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1792), .I3(n26119), 
            .O(n5518)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1484_3_lut (.I0(n1246), .I1(n5511), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[11]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1484_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1483_3_lut (.I0(n1168), .I1(n5510), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[12]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1483_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1482_3_lut (.I0(n1090), .I1(n5509), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[13]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1482_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1481_3_lut (.I0(n1012), .I1(n5508), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[14]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1481_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1480_3_lut (.I0(n934), .I1(n5507), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[15]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1480_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1479_3_lut (.I0(n856), .I1(n5506), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[16]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1479_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1478_3_lut (.I0(n778), .I1(n5505), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[17]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1478_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1477_3_lut (.I0(n700), .I1(n5504), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[18]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1477_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY add_1777_6 (.CI(n26119), .I0(GND_net), .I1(n1792), .CO(n26120));
    SB_LUT4 mux_59_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_59_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13579_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n30471), .I3(GND_net), .O(n18159));   // verilog/coms.v(127[12] 300[6])
    defparam i13579_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_50[21]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_50[20]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_50[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_50[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_50[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_50[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_50[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_50[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_50[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_50[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_50[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_50[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_50[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_50[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_50[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_50[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_50[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_50[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_50[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_50[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_50[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i13580_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n30471), .I3(GND_net), .O(n18160));   // verilog/coms.v(127[12] 300[6])
    defparam i13580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13581_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n30471), .I3(GND_net), .O(n18161));   // verilog/coms.v(127[12] 300[6])
    defparam i13581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_59_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_1777_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1870), .I3(n26118), 
            .O(n5519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13582_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n30471), .I3(GND_net), .O(n18162));   // verilog/coms.v(127[12] 300[6])
    defparam i13582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13583_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n30471), .I3(GND_net), .O(n18163));   // verilog/coms.v(127[12] 300[6])
    defparam i13583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13520_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n30475), .I3(GND_net), .O(n18100));   // verilog/coms.v(127[12] 300[6])
    defparam i13520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13584_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n30471), .I3(GND_net), .O(n18164));   // verilog/coms.v(127[12] 300[6])
    defparam i13584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13521_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n30475), .I3(GND_net), .O(n18101));   // verilog/coms.v(127[12] 300[6])
    defparam i13521_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1777_5 (.CI(n26118), .I0(GND_net), .I1(n1870), .CO(n26119));
    SB_LUT4 i13522_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n30475), .I3(GND_net), .O(n18102));   // verilog/coms.v(127[12] 300[6])
    defparam i13522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1777_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1948), .I3(n26117), 
            .O(n5520)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_4 (.CI(n26117), .I0(GND_net), .I1(n1948), .CO(n26118));
    SB_LUT4 add_1777_3_lut (.I0(GND_net), .I1(GND_net), .I2(n2026), .I3(n26116), 
            .O(n5521)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13585_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n30471), .I3(GND_net), .O(n18165));   // verilog/coms.v(127[12] 300[6])
    defparam i13585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13586_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n30471), .I3(GND_net), .O(n18166));   // verilog/coms.v(127[12] 300[6])
    defparam i13586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4899));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1373_3_lut (.I0(n2010), .I1(n2063), 
            .I2(n2026), .I3(GND_net), .O(n29_adj_4926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1374_3_lut (.I0(n2011), .I1(n2064), 
            .I2(n2026), .I3(GND_net), .O(n27_adj_4925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1365_3_lut (.I0(n2002), .I1(n2055), 
            .I2(n2026), .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1365_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1777_3 (.CI(n26116), .I0(GND_net), .I1(n2026), .CO(n26117));
    SB_LUT4 add_1777_2_lut (.I0(GND_net), .I1(GND_net), .I2(n22965), .I3(VCC_net), 
            .O(n5522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1777_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1777_2 (.CI(VCC_net), .I0(GND_net), .I1(n22965), .CO(n26116));
    SB_LUT4 encoder0_position_23__I_0_add_1308_24_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n26115), .O(n1975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_23_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n26114), .O(n1976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_23 (.CI(n26114), .I0(n1923), 
            .I1(VCC_net), .CO(n26115));
    SB_LUT4 encoder0_position_23__I_0_add_1308_22_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n26113), .O(n1977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_22 (.CI(n26113), .I0(n1924), 
            .I1(VCC_net), .CO(n26114));
    SB_LUT4 encoder0_position_23__I_0_add_1308_21_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n26112), .O(n1978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_21 (.CI(n26112), .I0(n1925), 
            .I1(VCC_net), .CO(n26113));
    SB_LUT4 encoder0_position_23__I_0_add_1308_20_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n26111), .O(n1979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_20 (.CI(n26111), .I0(n1926), 
            .I1(VCC_net), .CO(n26112));
    SB_LUT4 encoder0_position_23__I_0_add_1308_19_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n26110), .O(n1980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1381_3_lut (.I0(n2018), .I1(n2071), 
            .I2(n2026), .I3(GND_net), .O(n13_adj_4923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_19 (.CI(n26110), .I0(n1927), 
            .I1(VCC_net), .CO(n26111));
    SB_LUT4 encoder0_position_23__I_0_i1368_3_lut (.I0(n2005), .I1(n2058), 
            .I2(n2026), .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n2020), .I1(n33995), .I2(n2026), .I3(n2019), 
            .O(n5_adj_4830));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i27932_3_lut (.I0(n931), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n34036));
    defparam i27932_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 encoder0_position_23__I_0_i1363_3_lut (.I0(n2000), .I1(n2053), 
            .I2(n2026), .I3(GND_net), .O(n49));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1366_3_lut (.I0(n2003), .I1(n2056), 
            .I2(n2026), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_18_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n26109), .O(n1981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(n34036), .I1(n5_adj_4830), .I2(n34037), 
            .I3(n2026), .O(n28827));
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'h88c0;
    SB_CARRY encoder0_position_23__I_0_add_1308_18 (.CI(n26109), .I0(n1928), 
            .I1(VCC_net), .CO(n26110));
    SB_LUT4 encoder0_position_23__I_0_add_1308_17_lut (.I0(GND_net), .I1(n1929), 
            .I2(VCC_net), .I3(n26108), .O(n1982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1631 (.I0(n2016), .I1(n29_adj_4926), .I2(n2069), 
            .I3(n2026), .O(n24_adj_4955));
    defparam i4_4_lut_adj_1631.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_23__I_0_add_1308_17 (.CI(n26108), .I0(n1929), 
            .I1(VCC_net), .CO(n26109));
    SB_LUT4 encoder0_position_23__I_0_add_1308_16_lut (.I0(GND_net), .I1(n1930), 
            .I2(VCC_net), .I3(n26107), .O(n1983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1632 (.I0(n28827), .I1(n2001), .I2(n2054), .I3(n2026), 
            .O(n22_adj_4957));
    defparam i2_4_lut_adj_1632.LUT_INIT = 16'heefa;
    SB_DFFSR encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
            .C(clk32MHz), .D(n5501), .R(n2_adj_4899));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_CARRY encoder0_position_23__I_0_add_1308_16 (.CI(n26107), .I0(n1930), 
            .I1(VCC_net), .CO(n26108));
    SB_LUT4 encoder0_position_23__I_0_add_1308_15_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n26106), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1633 (.I0(n2007), .I1(n49), .I2(n2060), .I3(n2026), 
            .O(n23_adj_4956));
    defparam i3_4_lut_adj_1633.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_23__I_0_add_1308_15 (.CI(n26106), .I0(n1931), 
            .I1(VCC_net), .CO(n26107));
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n2014), .I1(n43), .I2(n2067), .I3(n2026), 
            .O(n21_adj_4958));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_23__I_0_add_1308_14_lut (.I0(GND_net), .I1(n1932), 
            .I2(VCC_net), .I3(n26105), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_14 (.CI(n26105), .I0(n1932), 
            .I1(VCC_net), .CO(n26106));
    SB_LUT4 encoder0_position_23__I_0_i1369_3_lut (.I0(n2006), .I1(n2059), 
            .I2(n2026), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1376_3_lut (.I0(n2013), .I1(n2066), 
            .I2(n2026), .I3(GND_net), .O(n23_adj_4924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_13_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n26104), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut (.I0(n2008), .I1(n27_adj_4925), .I2(n2061), .I3(n2026), 
            .O(n28_adj_4951));
    defparam i8_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i6_4_lut_adj_1635 (.I0(n2004), .I1(n45), .I2(n2057), .I3(n2026), 
            .O(n26_adj_4953));
    defparam i6_4_lut_adj_1635.LUT_INIT = 16'heefc;
    SB_DFFSR encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
            .C(clk32MHz), .D(n5502), .R(n2_adj_4899));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i7_4_lut_adj_1636 (.I0(n2012), .I1(n13_adj_4923), .I2(n2065), 
            .I3(n2026), .O(n27_adj_4952));
    defparam i7_4_lut_adj_1636.LUT_INIT = 16'heefc;
    SB_LUT4 i5_4_lut (.I0(n2017), .I1(n23_adj_4924), .I2(n2070), .I3(n2026), 
            .O(n25_adj_4954));
    defparam i5_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 i10_4_lut (.I0(n2009), .I1(n39), .I2(n2062), .I3(n2026), 
            .O(n30_adj_4949));
    defparam i10_4_lut.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_23__I_0_add_1308_13 (.CI(n26104), .I0(n1933), 
            .I1(VCC_net), .CO(n26105));
    SB_LUT4 i16_4_lut_adj_1637 (.I0(n21_adj_4958), .I1(n23_adj_4956), .I2(n22_adj_4957), 
            .I3(n24_adj_4955), .O(n36));
    defparam i16_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n2015), .I1(n37), .I2(n2068), .I3(n2026), 
            .O(n29_adj_4950));
    defparam i9_4_lut.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_23__I_0_add_1308_12_lut (.I0(GND_net), .I1(n1934), 
            .I2(VCC_net), .I3(n26103), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(n25_adj_4954), .I1(n27_adj_4952), .I2(n26_adj_4953), 
            .I3(n28_adj_4951), .O(n37_adj_4948));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_23__I_0_add_1308_12 (.CI(n26103), .I0(n1934), 
            .I1(VCC_net), .CO(n26104));
    SB_LUT4 i29240_4_lut (.I0(n37_adj_4948), .I1(n29_adj_4950), .I2(n36), 
            .I3(n30_adj_4949), .O(n22965));
    defparam i29240_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i11_4_lut (.I0(n2002), .I1(n2011), .I2(n2008), .I3(n2001), 
            .O(n30_adj_4942));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i463_3_lut (.I0(n675), .I1(n728), 
            .I2(n700), .I3(GND_net), .O(n753));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18306_3_lut (.I0(n931), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n22885));
    defparam i18306_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_615_14_lut (.I0(duty[12]), .I1(n35425), .I2(n13), .I3(n25596), 
            .O(pwm_setpoint_22__N_3[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut_adj_1638 (.I0(n2019), .I1(n2018), .I2(n22885), .I3(n2020), 
            .O(n31986));
    defparam i2_4_lut_adj_1638.LUT_INIT = 16'h8880;
    SB_LUT4 i15_4_lut (.I0(n2003), .I1(n30_adj_4942), .I2(n2015), .I3(n2014), 
            .O(n34_adj_4939));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1639 (.I0(n2000), .I1(n2016), .I2(n2010), .I3(n2006), 
            .O(n32));
    defparam i13_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_1308_11_lut (.I0(GND_net), .I1(n1935), 
            .I2(VCC_net), .I3(n26102), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut (.I0(n2009), .I1(n2004), .I2(n2013), .I3(n2007), 
            .O(n33_adj_4940));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2017), .I1(n2005), .I2(n2012), .I3(n31986), 
            .O(n31_adj_4941));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29236_4_lut (.I0(n31_adj_4941), .I1(n33_adj_4940), .I2(n32), 
            .I3(n34_adj_4939), .O(n2026));
    defparam i29236_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_23__I_0_add_1308_11 (.CI(n26102), .I0(n1935), 
            .I1(VCC_net), .CO(n26103));
    SB_LUT4 encoder0_position_23__I_0_add_1308_10_lut (.I0(GND_net), .I1(n1936), 
            .I2(VCC_net), .I3(n26101), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_10 (.CI(n26101), .I0(n1936), 
            .I1(VCC_net), .CO(n26102));
    SB_LUT4 encoder0_position_23__I_0_add_1308_9_lut (.I0(GND_net), .I1(n1937), 
            .I2(VCC_net), .I3(n26100), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_9 (.CI(n26100), .I0(n1937), 
            .I1(VCC_net), .CO(n26101));
    SB_LUT4 encoder0_position_23__I_0_add_1308_8_lut (.I0(GND_net), .I1(n1938), 
            .I2(VCC_net), .I3(n26099), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_8 (.CI(n26099), .I0(n1938), 
            .I1(VCC_net), .CO(n26100));
    SB_LUT4 encoder0_position_23__I_0_add_1308_7_lut (.I0(GND_net), .I1(n1939), 
            .I2(GND_net), .I3(n26098), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_7 (.CI(n26098), .I0(n1939), 
            .I1(GND_net), .CO(n26099));
    SB_LUT4 encoder0_position_23__I_0_add_1308_6_lut (.I0(GND_net), .I1(n1940), 
            .I2(GND_net), .I3(n26097), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_6 (.CI(n26097), .I0(n1940), 
            .I1(GND_net), .CO(n26098));
    SB_LUT4 encoder0_position_23__I_0_add_1308_5_lut (.I0(GND_net), .I1(n1941), 
            .I2(VCC_net), .I3(n26096), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_5 (.CI(n26096), .I0(n1941), 
            .I1(VCC_net), .CO(n26097));
    SB_LUT4 encoder0_position_23__I_0_add_1308_4_lut (.I0(GND_net), .I1(n1942), 
            .I2(GND_net), .I3(n26095), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_4 (.CI(n26095), .I0(n1942), 
            .I1(GND_net), .CO(n26096));
    SB_LUT4 encoder0_position_23__I_0_add_1308_3_lut (.I0(GND_net), .I1(n1943), 
            .I2(VCC_net), .I3(n26094), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_3 (.CI(n26094), .I0(n1943), 
            .I1(VCC_net), .CO(n26095));
    SB_LUT4 encoder0_position_23__I_0_add_1308_2_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(VCC_net), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_2 (.CI(VCC_net), .I0(n930), 
            .I1(GND_net), .CO(n26094));
    SB_LUT4 encoder0_position_23__I_0_add_1255_23_lut (.I0(GND_net), .I1(n1844), 
            .I2(VCC_net), .I3(n26093), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_22_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n26092), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_22 (.CI(n26092), .I0(n1845), 
            .I1(VCC_net), .CO(n26093));
    SB_LUT4 encoder0_position_23__I_0_add_1255_21_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n26091), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_21 (.CI(n26091), .I0(n1846), 
            .I1(VCC_net), .CO(n26092));
    SB_LUT4 encoder0_position_23__I_0_add_1255_20_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n26090), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_14 (.CI(n25596), .I0(n35425), .I1(n13), .CO(n25597));
    SB_CARRY encoder0_position_23__I_0_add_1255_20 (.CI(n26090), .I0(n1847), 
            .I1(VCC_net), .CO(n26091));
    SB_LUT4 encoder0_position_23__I_0_add_1255_19_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n26089), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_19 (.CI(n26089), .I0(n1848), 
            .I1(VCC_net), .CO(n26090));
    SB_LUT4 encoder0_position_23__I_0_add_1255_18_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n26088), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_18 (.CI(n26088), .I0(n1849), 
            .I1(VCC_net), .CO(n26089));
    SB_LUT4 encoder0_position_23__I_0_add_1255_17_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n26087), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_17 (.CI(n26087), .I0(n1850), 
            .I1(VCC_net), .CO(n26088));
    SB_LUT4 encoder0_position_23__I_0_add_1255_16_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n26086), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_16 (.CI(n26086), .I0(n1851), 
            .I1(VCC_net), .CO(n26087));
    SB_LUT4 encoder0_position_23__I_0_add_1255_15_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n26085), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_15 (.CI(n26085), .I0(n1852), 
            .I1(VCC_net), .CO(n26086));
    SB_LUT4 encoder0_position_23__I_0_add_1255_14_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n26084), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_14 (.CI(n26084), .I0(n1853), 
            .I1(VCC_net), .CO(n26085));
    SB_LUT4 encoder0_position_23__I_0_add_1255_13_lut (.I0(GND_net), .I1(n1854), 
            .I2(VCC_net), .I3(n26083), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_13_lut (.I0(duty[11]), .I1(n35425), .I2(n14), .I3(n25595), 
            .O(pwm_setpoint_22__N_3[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1255_13 (.CI(n26083), .I0(n1854), 
            .I1(VCC_net), .CO(n26084));
    SB_LUT4 encoder0_position_23__I_0_i465_3_lut (.I0(n677), .I1(n730), 
            .I2(n700), .I3(GND_net), .O(n755));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i467_3_lut (.I0(n679), .I1(n732), 
            .I2(n700), .I3(GND_net), .O(n757));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i466_3_lut (.I0(n678), .I1(n731), 
            .I2(n700), .I3(GND_net), .O(n756));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i464_3_lut (.I0(n676), .I1(n729), 
            .I2(n700), .I3(GND_net), .O(n754));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i468_3_lut (.I0(n515), .I1(n733), 
            .I2(n700), .I3(GND_net), .O(n758));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3158_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17636_2_lut (.I0(n516), .I1(n758), .I2(GND_net), .I3(GND_net), 
            .O(n22209));
    defparam i17636_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n754), .I1(n22209), .I2(n756), .I3(n757), 
            .O(n4_adj_4959));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'ha8a0;
    SB_LUT4 encoder0_position_23__I_0_add_1255_12_lut (.I0(GND_net), .I1(n1855), 
            .I2(VCC_net), .I3(n26082), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_12 (.CI(n26082), .I0(n1855), 
            .I1(VCC_net), .CO(n26083));
    SB_LUT4 encoder0_position_23__I_0_add_1255_11_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n26081), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_11 (.CI(n26081), .I0(n1856), 
            .I1(VCC_net), .CO(n26082));
    SB_LUT4 encoder0_position_23__I_0_add_1255_10_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n26080), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_10 (.CI(n26080), .I0(n1857), 
            .I1(VCC_net), .CO(n26081));
    SB_LUT4 encoder0_position_23__I_0_add_1255_9_lut (.I0(GND_net), .I1(n1858), 
            .I2(VCC_net), .I3(n26079), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_9 (.CI(n26079), .I0(n1858), 
            .I1(VCC_net), .CO(n26080));
    SB_LUT4 i28873_4_lut (.I0(n752), .I1(n755), .I2(n753), .I3(n4_adj_4959), 
            .O(n778));
    defparam i28873_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 i28862_1_lut (.I0(n778), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35036));
    defparam i28862_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25010_4_lut (.I0(encoder0_position[22]), .I1(n33988), .I2(encoder0_position[23]), 
            .I3(n3_adj_4829), .O(n675));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i25010_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i25008_3_lut (.I0(encoder0_position[21]), .I1(n31159), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n676));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i25008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25002_3_lut (.I0(encoder0_position[18]), .I1(n31153), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n679));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i25002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25004_3_lut (.I0(encoder0_position[19]), .I1(n31155), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n678));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i25004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25006_3_lut (.I0(encoder0_position[20]), .I1(n31157), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n677));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i25006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3158_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18416_4_lut (.I0(n515), .I1(n677), .I2(n678), .I3(n679), 
            .O(n22997));
    defparam i18416_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i28884_4_lut (.I0(n676), .I1(n674), .I2(n675), .I3(n22997), 
            .O(n700));
    defparam i28884_4_lut.LUT_INIT = 16'h1333;
    SB_LUT4 i1_2_lut (.I0(n514), .I1(n6), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4837));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1641 (.I0(n4_adj_4831), .I1(n2), .I2(n5), .I3(n7_adj_4837), 
            .O(n4_adj_4927));
    defparam i1_4_lut_adj_1641.LUT_INIT = 16'hc888;
    SB_LUT4 i3483_2_lut (.I0(n2), .I1(encoder0_position[23]), .I2(GND_net), 
            .I3(GND_net), .O(n509));
    defparam i3483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28874_1_lut (.I0(n700), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35048));
    defparam i28874_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1255_8_lut (.I0(GND_net), .I1(n1859), 
            .I2(VCC_net), .I3(n26078), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_8 (.CI(n26078), .I0(n1859), 
            .I1(VCC_net), .CO(n26079));
    SB_LUT4 encoder0_position_23__I_0_add_1255_7_lut (.I0(GND_net), .I1(n1860), 
            .I2(GND_net), .I3(n26077), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_7 (.CI(n26077), .I0(n1860), 
            .I1(GND_net), .CO(n26078));
    SB_LUT4 encoder0_position_23__I_0_add_1255_6_lut (.I0(GND_net), .I1(n1861), 
            .I2(GND_net), .I3(n26076), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_6 (.CI(n26076), .I0(n1861), 
            .I1(GND_net), .CO(n26077));
    SB_LUT4 encoder0_position_23__I_0_add_1255_5_lut (.I0(GND_net), .I1(n1862), 
            .I2(VCC_net), .I3(n26075), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_59_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_23__I_0_add_1255_5 (.CI(n26075), .I0(n1862), 
            .I1(VCC_net), .CO(n26076));
    SB_LUT4 encoder0_position_23__I_0_add_1255_4_lut (.I0(GND_net), .I1(n1863), 
            .I2(GND_net), .I3(n26074), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_26[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_3[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 mux_3158_i19_3_lut (.I0(encoder0_position[18]), .I1(n7), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n514));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1255_4 (.CI(n26074), .I0(n1863), 
            .I1(GND_net), .CO(n26075));
    SB_LUT4 encoder0_position_23__I_0_add_1255_3_lut (.I0(GND_net), .I1(n1864), 
            .I2(VCC_net), .I3(n26073), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_3 (.CI(n26073), .I0(n1864), 
            .I1(VCC_net), .CO(n26074));
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1255_2_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(VCC_net), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_2 (.CI(VCC_net), .I0(n929), 
            .I1(GND_net), .CO(n26073));
    SB_LUT4 encoder0_position_23__I_0_add_1202_22_lut (.I0(GND_net), .I1(n1766), 
            .I2(VCC_net), .I3(n26072), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1202_21_lut (.I0(GND_net), .I1(n1767), 
            .I2(VCC_net), .I3(n26071), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_21 (.CI(n26071), .I0(n1767), 
            .I1(VCC_net), .CO(n26072));
    SB_LUT4 encoder0_position_23__I_0_add_1202_20_lut (.I0(GND_net), .I1(n1768), 
            .I2(VCC_net), .I3(n26070), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_20 (.CI(n26070), .I0(n1768), 
            .I1(VCC_net), .CO(n26071));
    SB_LUT4 encoder0_position_23__I_0_add_1202_19_lut (.I0(GND_net), .I1(n1769), 
            .I2(VCC_net), .I3(n26069), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_19 (.CI(n26069), .I0(n1769), 
            .I1(VCC_net), .CO(n26070));
    SB_LUT4 encoder0_position_23__I_0_add_1202_18_lut (.I0(GND_net), .I1(n1770), 
            .I2(VCC_net), .I3(n26068), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_18 (.CI(n26068), .I0(n1770), 
            .I1(VCC_net), .CO(n26069));
    SB_CARRY add_615_13 (.CI(n25595), .I0(n35425), .I1(n14), .CO(n25596));
    SB_LUT4 encoder0_position_23__I_0_add_1202_17_lut (.I0(GND_net), .I1(n1771), 
            .I2(VCC_net), .I3(n26067), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_17 (.CI(n26067), .I0(n1771), 
            .I1(VCC_net), .CO(n26068));
    SB_LUT4 encoder0_position_23__I_0_add_1202_16_lut (.I0(GND_net), .I1(n1772), 
            .I2(VCC_net), .I3(n26066), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_16 (.CI(n26066), .I0(n1772), 
            .I1(VCC_net), .CO(n26067));
    SB_LUT4 encoder0_position_23__I_0_add_1202_15_lut (.I0(GND_net), .I1(n1773), 
            .I2(VCC_net), .I3(n26065), .O(n1826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_15 (.CI(n26065), .I0(n1773), 
            .I1(VCC_net), .CO(n26066));
    SB_LUT4 encoder0_position_23__I_0_add_1202_14_lut (.I0(GND_net), .I1(n1774), 
            .I2(VCC_net), .I3(n26064), .O(n1827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_14 (.CI(n26064), .I0(n1774), 
            .I1(VCC_net), .CO(n26065));
    SB_LUT4 encoder0_position_23__I_0_add_1202_13_lut (.I0(GND_net), .I1(n1775), 
            .I2(VCC_net), .I3(n26063), .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_13 (.CI(n26063), .I0(n1775), 
            .I1(VCC_net), .CO(n26064));
    SB_LUT4 encoder0_position_23__I_0_add_1202_12_lut (.I0(GND_net), .I1(n1776), 
            .I2(VCC_net), .I3(n26062), .O(n1829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_12 (.CI(n26062), .I0(n1776), 
            .I1(VCC_net), .CO(n26063));
    SB_LUT4 encoder0_position_23__I_0_add_1202_11_lut (.I0(GND_net), .I1(n1777), 
            .I2(VCC_net), .I3(n26061), .O(n1830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_11 (.CI(n26061), .I0(n1777), 
            .I1(VCC_net), .CO(n26062));
    SB_LUT4 encoder0_position_23__I_0_add_1202_10_lut (.I0(GND_net), .I1(n1778), 
            .I2(VCC_net), .I3(n26060), .O(n1831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_10 (.CI(n26060), .I0(n1778), 
            .I1(VCC_net), .CO(n26061));
    SB_LUT4 encoder0_position_23__I_0_add_1202_9_lut (.I0(GND_net), .I1(n1779), 
            .I2(VCC_net), .I3(n26059), .O(n1832)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_9 (.CI(n26059), .I0(n1779), 
            .I1(VCC_net), .CO(n26060));
    SB_LUT4 encoder0_position_23__I_0_add_1202_8_lut (.I0(GND_net), .I1(n1780), 
            .I2(VCC_net), .I3(n26058), .O(n1833)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_8 (.CI(n26058), .I0(n1780), 
            .I1(VCC_net), .CO(n26059));
    SB_LUT4 mux_59_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_1202_7_lut (.I0(GND_net), .I1(n1781), 
            .I2(GND_net), .I3(n26057), .O(n1834)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_7 (.CI(n26057), .I0(n1781), 
            .I1(GND_net), .CO(n26058));
    SB_LUT4 encoder0_position_23__I_0_add_1202_6_lut (.I0(GND_net), .I1(n1782), 
            .I2(GND_net), .I3(n26056), .O(n1835)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_6 (.CI(n26056), .I0(n1782), 
            .I1(GND_net), .CO(n26057));
    SB_LUT4 encoder0_position_23__I_0_add_1202_5_lut (.I0(GND_net), .I1(n1783), 
            .I2(VCC_net), .I3(n26055), .O(n1836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1642 (.I0(n22632), .I1(n16614), .I2(GND_net), 
            .I3(GND_net), .O(n4922));
    defparam i1_2_lut_adj_1642.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_23__I_0_add_1202_5 (.CI(n26055), .I0(n1783), 
            .I1(VCC_net), .CO(n26056));
    SB_LUT4 encoder0_position_23__I_0_add_1202_4_lut (.I0(GND_net), .I1(n1784), 
            .I2(GND_net), .I3(n26054), .O(n1837)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_4 (.CI(n26054), .I0(n1784), 
            .I1(GND_net), .CO(n26055));
    SB_LUT4 encoder0_position_23__I_0_add_1202_3_lut (.I0(GND_net), .I1(n1785), 
            .I2(VCC_net), .I3(n26053), .O(n1838)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_3 (.CI(n26053), .I0(n1785), 
            .I1(VCC_net), .CO(n26054));
    SB_LUT4 encoder0_position_23__I_0_add_1202_2_lut (.I0(GND_net), .I1(n928), 
            .I2(GND_net), .I3(VCC_net), .O(n1839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_2 (.CI(VCC_net), .I0(n928), 
            .I1(GND_net), .CO(n26053));
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4794));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1149_21_lut (.I0(GND_net), .I1(n1688), 
            .I2(VCC_net), .I3(n26052), .O(n1741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_20_lut (.I0(GND_net), .I1(n1689), 
            .I2(VCC_net), .I3(n26051), .O(n1742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_20 (.CI(n26051), .I0(n1689), 
            .I1(VCC_net), .CO(n26052));
    SB_LUT4 encoder0_position_23__I_0_add_1149_19_lut (.I0(GND_net), .I1(n1690), 
            .I2(VCC_net), .I3(n26050), .O(n1743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4816));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1149_19 (.CI(n26050), .I0(n1690), 
            .I1(VCC_net), .CO(n26051));
    SB_LUT4 encoder0_position_23__I_0_add_1149_18_lut (.I0(GND_net), .I1(n1691), 
            .I2(VCC_net), .I3(n26049), .O(n1744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_18 (.CI(n26049), .I0(n1691), 
            .I1(VCC_net), .CO(n26050));
    SB_LUT4 add_615_12_lut (.I0(duty[10]), .I1(n35425), .I2(n15), .I3(n25594), 
            .O(pwm_setpoint_22__N_3[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1149_17_lut (.I0(GND_net), .I1(n1692), 
            .I2(VCC_net), .I3(n26048), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_12 (.CI(n25594), .I0(n35425), .I1(n15), .CO(n25595));
    SB_CARRY encoder0_position_23__I_0_add_1149_17 (.CI(n26048), .I0(n1692), 
            .I1(VCC_net), .CO(n26049));
    SB_LUT4 encoder0_position_23__I_0_add_1149_16_lut (.I0(GND_net), .I1(n1693), 
            .I2(VCC_net), .I3(n26047), .O(n1746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_16 (.CI(n26047), .I0(n1693), 
            .I1(VCC_net), .CO(n26048));
    SB_LUT4 encoder0_position_23__I_0_add_1149_15_lut (.I0(GND_net), .I1(n1694), 
            .I2(VCC_net), .I3(n26046), .O(n1747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_15 (.CI(n26046), .I0(n1694), 
            .I1(VCC_net), .CO(n26047));
    SB_LUT4 encoder0_position_23__I_0_add_1149_14_lut (.I0(GND_net), .I1(n1695), 
            .I2(VCC_net), .I3(n26045), .O(n1748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_14 (.CI(n26045), .I0(n1695), 
            .I1(VCC_net), .CO(n26046));
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1149_13_lut (.I0(GND_net), .I1(n1696), 
            .I2(VCC_net), .I3(n26044), .O(n1749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_13 (.CI(n26044), .I0(n1696), 
            .I1(VCC_net), .CO(n26045));
    SB_LUT4 encoder0_position_23__I_0_add_1149_12_lut (.I0(GND_net), .I1(n1697), 
            .I2(VCC_net), .I3(n26043), .O(n1750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_12 (.CI(n26043), .I0(n1697), 
            .I1(VCC_net), .CO(n26044));
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_add_1149_11_lut (.I0(GND_net), .I1(n1698), 
            .I2(VCC_net), .I3(n26042), .O(n1751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_11 (.CI(n26042), .I0(n1698), 
            .I1(VCC_net), .CO(n26043));
    SB_LUT4 encoder0_position_23__I_0_add_1149_10_lut (.I0(GND_net), .I1(n1699), 
            .I2(VCC_net), .I3(n26041), .O(n1752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4793));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1149_10 (.CI(n26041), .I0(n1699), 
            .I1(VCC_net), .CO(n26042));
    SB_LUT4 encoder0_position_23__I_0_add_1149_9_lut (.I0(GND_net), .I1(n1700), 
            .I2(VCC_net), .I3(n26040), .O(n1753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_9 (.CI(n26040), .I0(n1700), 
            .I1(VCC_net), .CO(n26041));
    SB_LUT4 encoder0_position_23__I_0_add_1149_8_lut (.I0(GND_net), .I1(n1701), 
            .I2(VCC_net), .I3(n26039), .O(n1754)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3158_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4842), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1149_8 (.CI(n26039), .I0(n1701), 
            .I1(VCC_net), .CO(n26040));
    SB_LUT4 encoder0_position_23__I_0_add_1149_7_lut (.I0(GND_net), .I1(n1702), 
            .I2(GND_net), .I3(n26038), .O(n1755)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_7 (.CI(n26038), .I0(n1702), 
            .I1(GND_net), .CO(n26039));
    SB_LUT4 encoder0_position_23__I_0_add_1149_6_lut (.I0(GND_net), .I1(n1703), 
            .I2(GND_net), .I3(n26037), .O(n1756)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1332_3_lut (.I0(n930), .I1(n1997), 
            .I2(n1948), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1149_6 (.CI(n26037), .I0(n1703), 
            .I1(GND_net), .CO(n26038));
    SB_LUT4 encoder0_position_23__I_0_add_1149_5_lut (.I0(GND_net), .I1(n1704), 
            .I2(VCC_net), .I3(n26036), .O(n1757)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_5 (.CI(n26036), .I0(n1704), 
            .I1(VCC_net), .CO(n26037));
    SB_LUT4 encoder0_position_23__I_0_i1331_3_lut (.I0(n1943), .I1(n1996), 
            .I2(n1948), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4792));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1149_4_lut (.I0(GND_net), .I1(n1705), 
            .I2(GND_net), .I3(n26035), .O(n1758)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1330_3_lut (.I0(n1942), .I1(n1995), 
            .I2(n1948), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1149_4 (.CI(n26035), .I0(n1705), 
            .I1(GND_net), .CO(n26036));
    SB_LUT4 encoder0_position_23__I_0_add_1149_3_lut (.I0(GND_net), .I1(n1706), 
            .I2(VCC_net), .I3(n26034), .O(n1759)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_3 (.CI(n26034), .I0(n1706), 
            .I1(VCC_net), .CO(n26035));
    SB_LUT4 encoder0_position_23__I_0_i1329_3_lut (.I0(n1941), .I1(n1994), 
            .I2(n1948), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1149_2_lut (.I0(GND_net), .I1(n927), 
            .I2(GND_net), .I3(VCC_net), .O(n1760)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_2 (.CI(VCC_net), .I0(n927), 
            .I1(GND_net), .CO(n26034));
    SB_LUT4 encoder0_position_23__I_0_add_1096_20_lut (.I0(GND_net), .I1(n1610), 
            .I2(VCC_net), .I3(n26033), .O(n1663)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_19_lut (.I0(GND_net), .I1(n1611), 
            .I2(VCC_net), .I3(n26032), .O(n1664)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_19 (.CI(n26032), .I0(n1611), 
            .I1(VCC_net), .CO(n26033));
    SB_LUT4 encoder0_position_23__I_0_i1328_3_lut (.I0(n1940), .I1(n1993), 
            .I2(n1948), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1096_18_lut (.I0(GND_net), .I1(n1612), 
            .I2(VCC_net), .I3(n26031), .O(n1665)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1327_3_lut (.I0(n1939), .I1(n1992), 
            .I2(n1948), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_18 (.CI(n26031), .I0(n1612), 
            .I1(VCC_net), .CO(n26032));
    SB_LUT4 encoder0_position_23__I_0_add_1096_17_lut (.I0(GND_net), .I1(n1613), 
            .I2(VCC_net), .I3(n26030), .O(n1666)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_17 (.CI(n26030), .I0(n1613), 
            .I1(VCC_net), .CO(n26031));
    SB_LUT4 encoder0_position_23__I_0_add_1096_16_lut (.I0(GND_net), .I1(n1614), 
            .I2(VCC_net), .I3(n26029), .O(n1667)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1326_3_lut (.I0(n1938), .I1(n1991), 
            .I2(n1948), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1326_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_16 (.CI(n26029), .I0(n1614), 
            .I1(VCC_net), .CO(n26030));
    SB_LUT4 encoder0_position_23__I_0_add_1096_15_lut (.I0(GND_net), .I1(n1615), 
            .I2(VCC_net), .I3(n26028), .O(n1668)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1325_3_lut (.I0(n1937), .I1(n1990), 
            .I2(n1948), .I3(GND_net), .O(n2015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1325_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_15 (.CI(n26028), .I0(n1615), 
            .I1(VCC_net), .CO(n26029));
    SB_LUT4 add_615_11_lut (.I0(duty[9]), .I1(n35425), .I2(n16_adj_4795), 
            .I3(n25593), .O(pwm_setpoint_22__N_3[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1096_14_lut (.I0(GND_net), .I1(n1616), 
            .I2(VCC_net), .I3(n26027), .O(n1669)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_14 (.CI(n26027), .I0(n1616), 
            .I1(VCC_net), .CO(n26028));
    SB_LUT4 encoder0_position_23__I_0_add_1096_13_lut (.I0(GND_net), .I1(n1617), 
            .I2(VCC_net), .I3(n26026), .O(n1670)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_13 (.CI(n26026), .I0(n1617), 
            .I1(VCC_net), .CO(n26027));
    SB_LUT4 encoder0_position_23__I_0_add_1096_12_lut (.I0(GND_net), .I1(n1618), 
            .I2(VCC_net), .I3(n26025), .O(n1671)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1324_3_lut (.I0(n1936), .I1(n1989), 
            .I2(n1948), .I3(GND_net), .O(n2014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1323_3_lut (.I0(n1935), .I1(n1988), 
            .I2(n1948), .I3(GND_net), .O(n2013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1322_3_lut (.I0(n1934), .I1(n1987), 
            .I2(n1948), .I3(GND_net), .O(n2012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1322_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_12 (.CI(n26025), .I0(n1618), 
            .I1(VCC_net), .CO(n26026));
    SB_LUT4 encoder0_position_23__I_0_add_1096_11_lut (.I0(GND_net), .I1(n1619), 
            .I2(VCC_net), .I3(n26024), .O(n1672)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1321_3_lut (.I0(n1933), .I1(n1986), 
            .I2(n1948), .I3(GND_net), .O(n2011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_11 (.CI(n26024), .I0(n1619), 
            .I1(VCC_net), .CO(n26025));
    SB_LUT4 encoder0_position_23__I_0_add_1096_10_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n26023), .O(n1673)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_10 (.CI(n26023), .I0(n1620), 
            .I1(VCC_net), .CO(n26024));
    SB_LUT4 encoder0_position_23__I_0_add_1096_9_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n26022), .O(n1674)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1320_3_lut (.I0(n1932), .I1(n1985), 
            .I2(n1948), .I3(GND_net), .O(n2010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4791));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1096_9 (.CI(n26022), .I0(n1621), 
            .I1(VCC_net), .CO(n26023));
    SB_LUT4 encoder0_position_23__I_0_add_1096_8_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n26021), .O(n1675)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1319_3_lut (.I0(n1931), .I1(n1984), 
            .I2(n1948), .I3(GND_net), .O(n2009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_8 (.CI(n26021), .I0(n1622), 
            .I1(VCC_net), .CO(n26022));
    SB_LUT4 encoder0_position_23__I_0_add_1096_7_lut (.I0(GND_net), .I1(n1623), 
            .I2(GND_net), .I3(n26020), .O(n1676)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_7 (.CI(n26020), .I0(n1623), 
            .I1(GND_net), .CO(n26021));
    SB_LUT4 encoder0_position_23__I_0_add_1096_6_lut (.I0(GND_net), .I1(n1624), 
            .I2(GND_net), .I3(n26019), .O(n1677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_6 (.CI(n26019), .I0(n1624), 
            .I1(GND_net), .CO(n26020));
    SB_LUT4 encoder0_position_23__I_0_add_1096_5_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n26018), .O(n1678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_5 (.CI(n26018), .I0(n1625), 
            .I1(VCC_net), .CO(n26019));
    SB_LUT4 encoder0_position_23__I_0_add_1096_4_lut (.I0(GND_net), .I1(n1626), 
            .I2(GND_net), .I3(n26017), .O(n1679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_4 (.CI(n26017), .I0(n1626), 
            .I1(GND_net), .CO(n26018));
    SB_LUT4 encoder0_position_23__I_0_i1318_3_lut (.I0(n1930), .I1(n1983), 
            .I2(n1948), .I3(GND_net), .O(n2008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1096_3_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n26016), .O(n1680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_3 (.CI(n26016), .I0(n1627), 
            .I1(VCC_net), .CO(n26017));
    SB_LUT4 encoder0_position_23__I_0_add_1096_2_lut (.I0(GND_net), .I1(n926), 
            .I2(GND_net), .I3(VCC_net), .O(n1681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1317_3_lut (.I0(n1929), .I1(n1982), 
            .I2(n1948), .I3(GND_net), .O(n2007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_2 (.CI(VCC_net), .I0(n926), 
            .I1(GND_net), .CO(n26016));
    SB_LUT4 encoder0_position_23__I_0_add_1043_19_lut (.I0(GND_net), .I1(n1532), 
            .I2(VCC_net), .I3(n26015), .O(n1585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1043_18_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n26014), .O(n1586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_18 (.CI(n26014), .I0(n1533), 
            .I1(VCC_net), .CO(n26015));
    SB_LUT4 encoder0_position_23__I_0_i1316_3_lut (.I0(n1928), .I1(n1981), 
            .I2(n1948), .I3(GND_net), .O(n2006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_17_lut (.I0(GND_net), .I1(n1534), 
            .I2(VCC_net), .I3(n26013), .O(n1587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_17 (.CI(n26013), .I0(n1534), 
            .I1(VCC_net), .CO(n26014));
    SB_LUT4 encoder0_position_23__I_0_i1315_3_lut (.I0(n1927), .I1(n1980), 
            .I2(n1948), .I3(GND_net), .O(n2005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1314_3_lut (.I0(n1926), .I1(n1979), 
            .I2(n1948), .I3(GND_net), .O(n2004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_16_lut (.I0(GND_net), .I1(n1535), 
            .I2(VCC_net), .I3(n26012), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_16 (.CI(n26012), .I0(n1535), 
            .I1(VCC_net), .CO(n26013));
    SB_LUT4 encoder0_position_23__I_0_add_1043_15_lut (.I0(GND_net), .I1(n1536), 
            .I2(VCC_net), .I3(n26011), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_15 (.CI(n26011), .I0(n1536), 
            .I1(VCC_net), .CO(n26012));
    SB_LUT4 encoder0_position_23__I_0_add_1043_14_lut (.I0(GND_net), .I1(n1537), 
            .I2(VCC_net), .I3(n26010), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1313_3_lut (.I0(n1925), .I1(n1978), 
            .I2(n1948), .I3(GND_net), .O(n2003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1312_3_lut (.I0(n1924), .I1(n1977), 
            .I2(n1948), .I3(GND_net), .O(n2002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1311_3_lut (.I0(n1923), .I1(n1976), 
            .I2(n1948), .I3(GND_net), .O(n2001));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_615_11 (.CI(n25593), .I0(n35425), .I1(n16_adj_4795), 
            .CO(n25594));
    SB_LUT4 encoder0_position_23__I_0_i1264_3_lut (.I0(n1851), .I1(n1904), 
            .I2(n1870), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1261_3_lut (.I0(n1848), .I1(n1901), 
            .I2(n1870), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1268_3_lut (.I0(n1855), .I1(n1908), 
            .I2(n1870), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1259_3_lut (.I0(n1846), .I1(n1899), 
            .I2(n1870), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1043_14 (.CI(n26010), .I0(n1537), 
            .I1(VCC_net), .CO(n26011));
    SB_LUT4 encoder0_position_23__I_0_i1274_3_lut (.I0(n1861), .I1(n1914), 
            .I2(n1870), .I3(GND_net), .O(n1939));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1275_3_lut (.I0(n1862), .I1(n1915), 
            .I2(n1870), .I3(GND_net), .O(n1940));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_13_lut (.I0(GND_net), .I1(n1538), 
            .I2(VCC_net), .I3(n26009), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_13 (.CI(n26009), .I0(n1538), 
            .I1(VCC_net), .CO(n26010));
    SB_LUT4 encoder0_position_23__I_0_i1273_3_lut (.I0(n1860), .I1(n1913), 
            .I2(n1870), .I3(GND_net), .O(n1938));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_12_lut (.I0(GND_net), .I1(n1539), 
            .I2(VCC_net), .I3(n26008), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_12 (.CI(n26008), .I0(n1539), 
            .I1(VCC_net), .CO(n26009));
    SB_LUT4 encoder0_position_23__I_0_i1271_3_lut (.I0(n1858), .I1(n1911), 
            .I2(n1870), .I3(GND_net), .O(n1936));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_11_lut (.I0(GND_net), .I1(n1540), 
            .I2(VCC_net), .I3(n26007), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1269_3_lut (.I0(n1856), .I1(n1909), 
            .I2(n1870), .I3(GND_net), .O(n1934));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1266_3_lut (.I0(n1853), .I1(n1906), 
            .I2(n1870), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1043_11 (.CI(n26007), .I0(n1540), 
            .I1(VCC_net), .CO(n26008));
    SB_LUT4 encoder0_position_23__I_0_add_1043_10_lut (.I0(GND_net), .I1(n1541), 
            .I2(VCC_net), .I3(n26006), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1270_3_lut (.I0(n1857), .I1(n1910), 
            .I2(n1870), .I3(GND_net), .O(n1935));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1262_3_lut (.I0(n1849), .I1(n1902), 
            .I2(n1870), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1265_3_lut (.I0(n1852), .I1(n1905), 
            .I2(n1870), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1043_10 (.CI(n26006), .I0(n1541), 
            .I1(VCC_net), .CO(n26007));
    SB_LUT4 encoder0_position_23__I_0_add_1043_9_lut (.I0(GND_net), .I1(n1542), 
            .I2(VCC_net), .I3(n26005), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_9 (.CI(n26005), .I0(n1542), 
            .I1(VCC_net), .CO(n26006));
    SB_LUT4 encoder0_position_23__I_0_add_1043_8_lut (.I0(GND_net), .I1(n1543), 
            .I2(VCC_net), .I3(n26004), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1258_3_lut (.I0(n1845), .I1(n1898), 
            .I2(n1870), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1278_3_lut (.I0(n929), .I1(n1918), 
            .I2(n1870), .I3(GND_net), .O(n1943));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1277_3_lut (.I0(n1864), .I1(n1917), 
            .I2(n1870), .I3(GND_net), .O(n1942));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1276_3_lut (.I0(n1863), .I1(n1916), 
            .I2(n1870), .I3(GND_net), .O(n1941));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1276_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1043_8 (.CI(n26004), .I0(n1543), 
            .I1(VCC_net), .CO(n26005));
    SB_LUT4 encoder0_position_23__I_0_add_1043_7_lut (.I0(GND_net), .I1(n1544), 
            .I2(GND_net), .I3(n26003), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3158_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4839), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_7 (.CI(n26003), .I0(n1544), 
            .I1(GND_net), .CO(n26004));
    SB_LUT4 encoder0_position_23__I_0_i1217_3_lut (.I0(n1779), .I1(n1832), 
            .I2(n1792), .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_6_lut (.I0(GND_net), .I1(n1545), 
            .I2(GND_net), .I3(n26002), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_6 (.CI(n26002), .I0(n1545), 
            .I1(GND_net), .CO(n26003));
    SB_LUT4 encoder0_position_23__I_0_add_1043_5_lut (.I0(GND_net), .I1(n1546), 
            .I2(VCC_net), .I3(n26001), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1215_3_lut (.I0(n1777), .I1(n1830), 
            .I2(n1792), .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1218_3_lut (.I0(n1780), .I1(n1833), 
            .I2(n1792), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1214_3_lut (.I0(n1776), .I1(n1829), 
            .I2(n1792), .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1213_3_lut (.I0(n1775), .I1(n1828), 
            .I2(n1792), .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1206_3_lut (.I0(n1768), .I1(n1821), 
            .I2(n1792), .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1209_3_lut (.I0(n1771), .I1(n1824), 
            .I2(n1792), .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1216_3_lut (.I0(n1778), .I1(n1831), 
            .I2(n1792), .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1210_3_lut (.I0(n1772), .I1(n1825), 
            .I2(n1792), .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1210_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1043_5 (.CI(n26001), .I0(n1546), 
            .I1(VCC_net), .CO(n26002));
    SB_LUT4 encoder0_position_23__I_0_i1205_3_lut (.I0(n1767), .I1(n1820), 
            .I2(n1792), .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_4_lut (.I0(GND_net), .I1(n1547), 
            .I2(GND_net), .I3(n26000), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_4 (.CI(n26000), .I0(n1547), 
            .I1(GND_net), .CO(n26001));
    SB_LUT4 encoder0_position_23__I_0_add_1043_3_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n25999), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_3 (.CI(n25999), .I0(n1548), 
            .I1(VCC_net), .CO(n26000));
    SB_LUT4 encoder0_position_23__I_0_i1212_3_lut (.I0(n1774), .I1(n1827), 
            .I2(n1792), .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1207_3_lut (.I0(n1769), .I1(n1822), 
            .I2(n1792), .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1204_3_lut (.I0(n1766), .I1(n1819), 
            .I2(n1792), .I3(GND_net), .O(n1844));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_2_lut (.I0(GND_net), .I1(n925), 
            .I2(GND_net), .I3(VCC_net), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_2 (.CI(VCC_net), .I0(n925), 
            .I1(GND_net), .CO(n25999));
    SB_LUT4 encoder0_position_23__I_0_add_990_18_lut (.I0(GND_net), .I1(n1454), 
            .I2(VCC_net), .I3(n25998), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1222_3_lut (.I0(n1784), .I1(n1837), 
            .I2(n1792), .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_17_lut (.I0(GND_net), .I1(n1455), 
            .I2(VCC_net), .I3(n25997), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1220_3_lut (.I0(n1782), .I1(n1835), 
            .I2(n1792), .I3(GND_net), .O(n1860));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1221_3_lut (.I0(n1783), .I1(n1836), 
            .I2(n1792), .I3(GND_net), .O(n1861));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1208_3_lut (.I0(n1770), .I1(n1823), 
            .I2(n1792), .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1211_3_lut (.I0(n1773), .I1(n1826), 
            .I2(n1792), .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1211_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_990_17 (.CI(n25997), .I0(n1455), 
            .I1(VCC_net), .CO(n25998));
    SB_LUT4 encoder0_position_23__I_0_add_990_16_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n25996), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_16 (.CI(n25996), .I0(n1456), 
            .I1(VCC_net), .CO(n25997));
    SB_LUT4 encoder0_position_23__I_0_i1165_3_lut (.I0(n1702), .I1(n1755), 
            .I2(n1714), .I3(GND_net), .O(n1780));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_15_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n25995), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_15 (.CI(n25995), .I0(n1457), 
            .I1(VCC_net), .CO(n25996));
    SB_LUT4 encoder0_position_23__I_0_add_990_14_lut (.I0(GND_net), .I1(n1458), 
            .I2(VCC_net), .I3(n25994), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_14 (.CI(n25994), .I0(n1458), 
            .I1(VCC_net), .CO(n25995));
    SB_LUT4 encoder0_position_23__I_0_add_990_13_lut (.I0(GND_net), .I1(n1459), 
            .I2(VCC_net), .I3(n25993), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_13 (.CI(n25993), .I0(n1459), 
            .I1(VCC_net), .CO(n25994));
    SB_LUT4 encoder0_position_23__I_0_add_990_12_lut (.I0(GND_net), .I1(n1460), 
            .I2(VCC_net), .I3(n25992), .O(n1513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_12 (.CI(n25992), .I0(n1460), 
            .I1(VCC_net), .CO(n25993));
    SB_LUT4 encoder0_position_23__I_0_i1154_3_lut (.I0(n1691), .I1(n1744), 
            .I2(n1714), .I3(GND_net), .O(n1769));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1161_3_lut (.I0(n1698), .I1(n1751), 
            .I2(n1714), .I3(GND_net), .O(n1776));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1153_3_lut (.I0(n1690), .I1(n1743), 
            .I2(n1714), .I3(GND_net), .O(n1768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1159_3_lut (.I0(n1696), .I1(n1749), 
            .I2(n1714), .I3(GND_net), .O(n1774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_11_lut (.I0(GND_net), .I1(n1461), 
            .I2(VCC_net), .I3(n25991), .O(n1514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_11 (.CI(n25991), .I0(n1461), 
            .I1(VCC_net), .CO(n25992));
    SB_LUT4 encoder0_position_23__I_0_i1162_3_lut (.I0(n1699), .I1(n1752), 
            .I2(n1714), .I3(GND_net), .O(n1777));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1163_3_lut (.I0(n1700), .I1(n1753), 
            .I2(n1714), .I3(GND_net), .O(n1778));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_10_lut (.I0(GND_net), .I1(n1462), 
            .I2(VCC_net), .I3(n25990), .O(n1515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_10 (.CI(n25990), .I0(n1462), 
            .I1(VCC_net), .CO(n25991));
    SB_LUT4 encoder0_position_23__I_0_i1156_3_lut (.I0(n1693), .I1(n1746), 
            .I2(n1714), .I3(GND_net), .O(n1771));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_9_lut (.I0(GND_net), .I1(n1463), 
            .I2(VCC_net), .I3(n25989), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1151_3_lut (.I0(n1688), .I1(n1741), 
            .I2(n1714), .I3(GND_net), .O(n1766));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1151_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_990_9 (.CI(n25989), .I0(n1463), 
            .I1(VCC_net), .CO(n25990));
    SB_LUT4 encoder0_position_23__I_0_i1158_3_lut (.I0(n1695), .I1(n1748), 
            .I2(n1714), .I3(GND_net), .O(n1773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_8_lut (.I0(GND_net), .I1(n1464), 
            .I2(VCC_net), .I3(n25988), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_8 (.CI(n25988), .I0(n1464), 
            .I1(VCC_net), .CO(n25989));
    SB_LUT4 encoder0_position_23__I_0_add_990_7_lut (.I0(GND_net), .I1(n1465), 
            .I2(GND_net), .I3(n25987), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_7 (.CI(n25987), .I0(n1465), 
            .I1(GND_net), .CO(n25988));
    SB_LUT4 encoder0_position_23__I_0_add_990_6_lut (.I0(GND_net), .I1(n1466), 
            .I2(GND_net), .I3(n25986), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1155_3_lut (.I0(n1692), .I1(n1745), 
            .I2(n1714), .I3(GND_net), .O(n1770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1164_3_lut (.I0(n1701), .I1(n1754), 
            .I2(n1714), .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1160_3_lut (.I0(n1697), .I1(n1750), 
            .I2(n1714), .I3(GND_net), .O(n1775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1152_3_lut (.I0(n1689), .I1(n1742), 
            .I2(n1714), .I3(GND_net), .O(n1767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1157_3_lut (.I0(n1694), .I1(n1747), 
            .I2(n1714), .I3(GND_net), .O(n1772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1168_3_lut (.I0(n1705), .I1(n1758), 
            .I2(n1714), .I3(GND_net), .O(n1783));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1168_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_990_6 (.CI(n25986), .I0(n1466), 
            .I1(GND_net), .CO(n25987));
    SB_LUT4 encoder0_position_23__I_0_i1166_3_lut (.I0(n1703), .I1(n1756), 
            .I2(n1714), .I3(GND_net), .O(n1781));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1167_3_lut (.I0(n1704), .I1(n1757), 
            .I2(n1714), .I3(GND_net), .O(n1782));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1109_3_lut (.I0(n1621), .I1(n1674), 
            .I2(n1636), .I3(GND_net), .O(n1699));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1106_3_lut (.I0(n1618), .I1(n1671), 
            .I2(n1636), .I3(GND_net), .O(n1696));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_990_5_lut (.I0(GND_net), .I1(n1467), 
            .I2(VCC_net), .I3(n25985), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1100_3_lut (.I0(n1612), .I1(n1665), 
            .I2(n1636), .I3(GND_net), .O(n1690));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1099_3_lut (.I0(n1611), .I1(n1664), 
            .I2(n1636), .I3(GND_net), .O(n1689));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1099_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_990_5 (.CI(n25985), .I0(n1467), 
            .I1(VCC_net), .CO(n25986));
    SB_LUT4 encoder0_position_23__I_0_i1101_3_lut (.I0(n1613), .I1(n1666), 
            .I2(n1636), .I3(GND_net), .O(n1691));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1104_3_lut (.I0(n1616), .I1(n1669), 
            .I2(n1636), .I3(GND_net), .O(n1694));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_10_lut (.I0(duty[8]), .I1(n35425), .I2(n17), .I3(n25592), 
            .O(pwm_setpoint_22__N_3[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_990_4_lut (.I0(GND_net), .I1(n1468), 
            .I2(GND_net), .I3(n25984), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1107_3_lut (.I0(n1619), .I1(n1672), 
            .I2(n1636), .I3(GND_net), .O(n1697));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_990_4 (.CI(n25984), .I0(n1468), 
            .I1(GND_net), .CO(n25985));
    SB_CARRY add_615_10 (.CI(n25592), .I0(n35425), .I1(n17), .CO(n25593));
    SB_LUT4 encoder0_position_23__I_0_add_990_3_lut (.I0(GND_net), .I1(n1469), 
            .I2(VCC_net), .I3(n25983), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_3 (.CI(n25983), .I0(n1469), 
            .I1(VCC_net), .CO(n25984));
    SB_LUT4 encoder0_position_23__I_0_add_990_2_lut (.I0(GND_net), .I1(n924), 
            .I2(GND_net), .I3(VCC_net), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_2 (.CI(VCC_net), .I0(n924), 
            .I1(GND_net), .CO(n25983));
    SB_LUT4 encoder0_position_23__I_0_i1103_3_lut (.I0(n1615), .I1(n1668), 
            .I2(n1636), .I3(GND_net), .O(n1693));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1108_3_lut (.I0(n1620), .I1(n1673), 
            .I2(n1636), .I3(GND_net), .O(n1698));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1111_3_lut (.I0(n1623), .I1(n1676), 
            .I2(n1636), .I3(GND_net), .O(n1701));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1102_3_lut (.I0(n1614), .I1(n1667), 
            .I2(n1636), .I3(GND_net), .O(n1692));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_17_lut (.I0(GND_net), .I1(n1376), 
            .I2(VCC_net), .I3(n25982), .O(n1429)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_16_lut (.I0(GND_net), .I1(n1377), 
            .I2(VCC_net), .I3(n25981), .O(n1430)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_16 (.CI(n25981), .I0(n1377), 
            .I1(VCC_net), .CO(n25982));
    SB_LUT4 encoder0_position_23__I_0_i1105_3_lut (.I0(n1617), .I1(n1670), 
            .I2(n1636), .I3(GND_net), .O(n1695));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_15_lut (.I0(GND_net), .I1(n1378), 
            .I2(VCC_net), .I3(n25980), .O(n1431)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1098_3_lut (.I0(n1610), .I1(n1663), 
            .I2(n1636), .I3(GND_net), .O(n1688));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1116_3_lut (.I0(n926), .I1(n1681), 
            .I2(n1636), .I3(GND_net), .O(n1706));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_15 (.CI(n25980), .I0(n1378), 
            .I1(VCC_net), .CO(n25981));
    SB_LUT4 encoder0_position_23__I_0_i1115_3_lut (.I0(n1627), .I1(n1680), 
            .I2(n1636), .I3(GND_net), .O(n1705));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1114_3_lut (.I0(n1626), .I1(n1679), 
            .I2(n1636), .I3(GND_net), .O(n1704));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1054_3_lut (.I0(n1541), .I1(n1594), 
            .I2(n1558), .I3(GND_net), .O(n1619));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1056_3_lut (.I0(n1543), .I1(n1596), 
            .I2(n1558), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_9_lut (.I0(duty[7]), .I1(n35425), .I2(n18), .I3(n25591), 
            .O(pwm_setpoint_22__N_3[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_937_14_lut (.I0(GND_net), .I1(n1379), 
            .I2(VCC_net), .I3(n25979), .O(n1432)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1046_3_lut (.I0(n1533), .I1(n1586), 
            .I2(n1558), .I3(GND_net), .O(n1611));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1051_3_lut (.I0(n1538), .I1(n1591), 
            .I2(n1558), .I3(GND_net), .O(n1616));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1055_3_lut (.I0(n1542), .I1(n1595), 
            .I2(n1558), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1057_3_lut (.I0(n1544), .I1(n1597), 
            .I2(n1558), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1057_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_14 (.CI(n25979), .I0(n1379), 
            .I1(VCC_net), .CO(n25980));
    SB_LUT4 encoder0_position_23__I_0_i1045_3_lut (.I0(n1532), .I1(n1585), 
            .I2(n1558), .I3(GND_net), .O(n1610));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1052_3_lut (.I0(n1539), .I1(n1592), 
            .I2(n1558), .I3(GND_net), .O(n1617));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13643_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n30466), 
            .I3(GND_net), .O(n18223));   // verilog/coms.v(127[12] 300[6])
    defparam i13643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13644_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n30466), 
            .I3(GND_net), .O(n18224));   // verilog/coms.v(127[12] 300[6])
    defparam i13644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1050_3_lut (.I0(n1537), .I1(n1590), 
            .I2(n1558), .I3(GND_net), .O(n1615));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1047_3_lut (.I0(n1534), .I1(n1587), 
            .I2(n1558), .I3(GND_net), .O(n1612));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1049_3_lut (.I0(n1536), .I1(n1589), 
            .I2(n1558), .I3(GND_net), .O(n1614));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13645_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n30466), 
            .I3(GND_net), .O(n18225));   // verilog/coms.v(127[12] 300[6])
    defparam i13645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1048_3_lut (.I0(n1535), .I1(n1588), 
            .I2(n1558), .I3(GND_net), .O(n1613));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1053_3_lut (.I0(n1540), .I1(n1593), 
            .I2(n1558), .I3(GND_net), .O(n1618));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1060_3_lut (.I0(n1547), .I1(n1600), 
            .I2(n1558), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1058_3_lut (.I0(n1545), .I1(n1598), 
            .I2(n1558), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_13_lut (.I0(GND_net), .I1(n1380), 
            .I2(VCC_net), .I3(n25978), .O(n1433)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1003_3_lut (.I0(n1465), .I1(n1518), 
            .I2(n1480), .I3(GND_net), .O(n1543));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i996_3_lut (.I0(n1458), .I1(n1511), 
            .I2(n1480), .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13646_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n30466), 
            .I3(GND_net), .O(n18226));   // verilog/coms.v(127[12] 300[6])
    defparam i13646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i999_3_lut (.I0(n1461), .I1(n1514), 
            .I2(n1480), .I3(GND_net), .O(n1539));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1001_3_lut (.I0(n1463), .I1(n1516), 
            .I2(n1480), .I3(GND_net), .O(n1541));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i995_3_lut (.I0(n1457), .I1(n1510), 
            .I2(n1480), .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13647_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n30466), 
            .I3(GND_net), .O(n18227));   // verilog/coms.v(127[12] 300[6])
    defparam i13647_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_13 (.CI(n25978), .I0(n1380), 
            .I1(VCC_net), .CO(n25979));
    SB_LUT4 encoder0_position_23__I_0_add_937_12_lut (.I0(GND_net), .I1(n1381), 
            .I2(VCC_net), .I3(n25977), .O(n1434)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1000_3_lut (.I0(n1462), .I1(n1515), 
            .I2(n1480), .I3(GND_net), .O(n1540));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1000_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_12 (.CI(n25977), .I0(n1381), 
            .I1(VCC_net), .CO(n25978));
    SB_LUT4 encoder0_position_23__I_0_i998_3_lut (.I0(n1460), .I1(n1513), 
            .I2(n1480), .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_11_lut (.I0(GND_net), .I1(n1382), 
            .I2(VCC_net), .I3(n25976), .O(n1435)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_11 (.CI(n25976), .I0(n1382), 
            .I1(VCC_net), .CO(n25977));
    SB_LUT4 encoder0_position_23__I_0_i1002_3_lut (.I0(n1464), .I1(n1517), 
            .I2(n1480), .I3(GND_net), .O(n1542));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i993_3_lut (.I0(n1455), .I1(n1508), 
            .I2(n1480), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13648_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n30466), 
            .I3(GND_net), .O(n18228));   // verilog/coms.v(127[12] 300[6])
    defparam i13648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i992_3_lut (.I0(n1454), .I1(n1507), 
            .I2(n1480), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i997_3_lut (.I0(n1459), .I1(n1512), 
            .I2(n1480), .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1004_3_lut (.I0(n1466), .I1(n1519), 
            .I2(n1480), .I3(GND_net), .O(n1544));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13649_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n30466), 
            .I3(GND_net), .O(n18229));   // verilog/coms.v(127[12] 300[6])
    defparam i13649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i994_3_lut (.I0(n1456), .I1(n1509), 
            .I2(n1480), .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_10_lut (.I0(GND_net), .I1(n1383), 
            .I2(VCC_net), .I3(n25975), .O(n1436)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_10 (.CI(n25975), .I0(n1383), 
            .I1(VCC_net), .CO(n25976));
    SB_LUT4 encoder0_position_23__I_0_add_937_9_lut (.I0(GND_net), .I1(n1384), 
            .I2(VCC_net), .I3(n25974), .O(n1437)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_9 (.CI(n25974), .I0(n1384), 
            .I1(VCC_net), .CO(n25975));
    SB_LUT4 encoder0_position_23__I_0_add_937_8_lut (.I0(GND_net), .I1(n1385), 
            .I2(VCC_net), .I3(n25973), .O(n1438)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_8 (.CI(n25973), .I0(n1385), 
            .I1(VCC_net), .CO(n25974));
    SB_LUT4 encoder0_position_23__I_0_add_937_7_lut (.I0(GND_net), .I1(n1386), 
            .I2(GND_net), .I3(n25972), .O(n1439)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_7 (.CI(n25972), .I0(n1386), 
            .I1(GND_net), .CO(n25973));
    SB_LUT4 encoder0_position_23__I_0_add_937_6_lut (.I0(GND_net), .I1(n1387), 
            .I2(GND_net), .I3(n25971), .O(n1440)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1005_3_lut (.I0(n1467), .I1(n1520), 
            .I2(n1480), .I3(GND_net), .O(n1545));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i940_3_lut (.I0(n1377), .I1(n1430), 
            .I2(n1402), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13650_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n30466), 
            .I3(GND_net), .O(n18230));   // verilog/coms.v(127[12] 300[6])
    defparam i13650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i947_3_lut (.I0(n1384), .I1(n1437), 
            .I2(n1402), .I3(GND_net), .O(n1462));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i939_3_lut (.I0(n1376), .I1(n1429), 
            .I2(n1402), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i945_3_lut (.I0(n1382), .I1(n1435), 
            .I2(n1402), .I3(GND_net), .O(n1460));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i944_3_lut (.I0(n1381), .I1(n1434), 
            .I2(n1402), .I3(GND_net), .O(n1459));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i946_3_lut (.I0(n1383), .I1(n1436), 
            .I2(n1402), .I3(GND_net), .O(n1461));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i950_3_lut (.I0(n1387), .I1(n1440), 
            .I2(n1402), .I3(GND_net), .O(n1465));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i951_3_lut (.I0(n1388), .I1(n1441), 
            .I2(n1402), .I3(GND_net), .O(n1466));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i951_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_6 (.CI(n25971), .I0(n1387), 
            .I1(GND_net), .CO(n25972));
    SB_LUT4 encoder0_position_23__I_0_i942_3_lut (.I0(n1379), .I1(n1432), 
            .I2(n1402), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_5_lut (.I0(GND_net), .I1(n1388), 
            .I2(VCC_net), .I3(n25970), .O(n1441)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i941_3_lut (.I0(n1378), .I1(n1431), 
            .I2(n1402), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i941_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_5 (.CI(n25970), .I0(n1388), 
            .I1(VCC_net), .CO(n25971));
    SB_LUT4 encoder0_position_23__I_0_i948_3_lut (.I0(n1385), .I1(n1438), 
            .I2(n1402), .I3(GND_net), .O(n1463));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i943_3_lut (.I0(n1380), .I1(n1433), 
            .I2(n1402), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_4_lut (.I0(GND_net), .I1(n1389), 
            .I2(GND_net), .I3(n25969), .O(n1442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i949_3_lut (.I0(n1386), .I1(n1439), 
            .I2(n1402), .I3(GND_net), .O(n1464));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i892_3_lut (.I0(n1304), .I1(n1357), 
            .I2(n1324), .I3(GND_net), .O(n1382));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i886_3_lut (.I0(n1298), .I1(n1351), 
            .I2(n1324), .I3(GND_net), .O(n1376));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i891_3_lut (.I0(n1303), .I1(n1356), 
            .I2(n1324), .I3(GND_net), .O(n1381));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i895_3_lut (.I0(n1307), .I1(n1360), 
            .I2(n1324), .I3(GND_net), .O(n1385));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i887_3_lut (.I0(n1299), .I1(n1352), 
            .I2(n1324), .I3(GND_net), .O(n1377));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i890_3_lut (.I0(n1302), .I1(n1355), 
            .I2(n1324), .I3(GND_net), .O(n1380));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i890_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_615_9 (.CI(n25591), .I0(n35425), .I1(n18), .CO(n25592));
    SB_LUT4 encoder0_position_23__I_0_i893_3_lut (.I0(n1305), .I1(n1358), 
            .I2(n1324), .I3(GND_net), .O(n1383));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i898_3_lut (.I0(n1310), .I1(n1363), 
            .I2(n1324), .I3(GND_net), .O(n1388));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i898_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_937_4 (.CI(n25969), .I0(n1389), 
            .I1(GND_net), .CO(n25970));
    SB_LUT4 encoder0_position_23__I_0_i896_3_lut (.I0(n1308), .I1(n1361), 
            .I2(n1324), .I3(GND_net), .O(n1386));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_3_lut (.I0(GND_net), .I1(n1390), 
            .I2(VCC_net), .I3(n25968), .O(n1443)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_3 (.CI(n25968), .I0(n1390), 
            .I1(VCC_net), .CO(n25969));
    SB_LUT4 encoder0_position_23__I_0_i897_3_lut (.I0(n1309), .I1(n1362), 
            .I2(n1324), .I3(GND_net), .O(n1387));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_937_2_lut (.I0(GND_net), .I1(n923), 
            .I2(GND_net), .I3(VCC_net), .O(n1444)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i900_3_lut (.I0(n922), .I1(n1365), 
            .I2(n1324), .I3(GND_net), .O(n1390));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_8_lut (.I0(duty[6]), .I1(n35425), .I2(n19_adj_4796), 
            .I3(n25590), .O(pwm_setpoint_22__N_3[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_937_2 (.CI(VCC_net), .I0(n923), 
            .I1(GND_net), .CO(n25968));
    SB_LUT4 encoder0_position_23__I_0_i899_3_lut (.I0(n1311), .I1(n1364), 
            .I2(n1324), .I3(GND_net), .O(n1389));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i840_3_lut (.I0(n1227), .I1(n1280), 
            .I2(n1246), .I3(GND_net), .O(n1305));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i837_3_lut (.I0(n1224), .I1(n1277), 
            .I2(n1246), .I3(GND_net), .O(n1302));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i839_3_lut (.I0(n1226), .I1(n1279), 
            .I2(n1246), .I3(GND_net), .O(n1304));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i834_3_lut (.I0(n1221), .I1(n1274), 
            .I2(n1246), .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i833_3_lut (.I0(n1220), .I1(n1273), 
            .I2(n1246), .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i836_3_lut (.I0(n1223), .I1(n1276), 
            .I2(n1246), .I3(GND_net), .O(n1301));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_615_8 (.CI(n25590), .I0(n35425), .I1(n19_adj_4796), .CO(n25591));
    SB_LUT4 encoder0_position_23__I_0_i844_3_lut (.I0(n1231), .I1(n1284), 
            .I2(n1246), .I3(GND_net), .O(n1309));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i842_3_lut (.I0(n1229), .I1(n1282), 
            .I2(n1246), .I3(GND_net), .O(n1307));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i843_3_lut (.I0(n1230), .I1(n1283), 
            .I2(n1246), .I3(GND_net), .O(n1308));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i846_3_lut (.I0(n435), .I1(n1286), 
            .I2(n1246), .I3(GND_net), .O(n1311));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i845_3_lut (.I0(n1232), .I1(n1285), 
            .I2(n1246), .I3(GND_net), .O(n1310));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3158_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i780_3_lut (.I0(n1142), .I1(n1195), 
            .I2(n1168), .I3(GND_net), .O(n1220));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i786_3_lut (.I0(n1148), .I1(n1201), 
            .I2(n1168), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i781_3_lut (.I0(n1143), .I1(n1196), 
            .I2(n1168), .I3(GND_net), .O(n1221));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i787_3_lut (.I0(n1149), .I1(n1202), 
            .I2(n1168), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i788_3_lut (.I0(n1150), .I1(n1203), 
            .I2(n1168), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i782_3_lut (.I0(n1144), .I1(n1197), 
            .I2(n1168), .I3(GND_net), .O(n1222));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i789_3_lut (.I0(n1151), .I1(n1204), 
            .I2(n1168), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i784_3_lut (.I0(n1146), .I1(n1199), 
            .I2(n1168), .I3(GND_net), .O(n1224));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i783_3_lut (.I0(n1145), .I1(n1198), 
            .I2(n1168), .I3(GND_net), .O(n1223));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i728_3_lut (.I0(n1065), .I1(n1118), 
            .I2(n1090), .I3(GND_net), .O(n1143));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i727_3_lut (.I0(n1064), .I1(n1117), 
            .I2(n1090), .I3(GND_net), .O(n1142));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i734_3_lut (.I0(n1071), .I1(n1124), 
            .I2(n1090), .I3(GND_net), .O(n1149));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i730_3_lut (.I0(n1067), .I1(n1120), 
            .I2(n1090), .I3(GND_net), .O(n1145));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i730_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i735_3_lut (.I0(n1072), .I1(n1125), 
            .I2(n1090), .I3(GND_net), .O(n1150));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i732_3_lut (.I0(n1069), .I1(n1122), 
            .I2(n1090), .I3(GND_net), .O(n1147));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i729_3_lut (.I0(n1066), .I1(n1119), 
            .I2(n1090), .I3(GND_net), .O(n1144));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i733_3_lut (.I0(n1070), .I1(n1123), 
            .I2(n1090), .I3(GND_net), .O(n1148));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i731_3_lut (.I0(n1068), .I1(n1121), 
            .I2(n1090), .I3(GND_net), .O(n1146));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i679_3_lut (.I0(n991), .I1(n1044), 
            .I2(n1012), .I3(GND_net), .O(n1069));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i676_3_lut (.I0(n988), .I1(n1041), 
            .I2(n1012), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i677_3_lut (.I0(n989), .I1(n1042), 
            .I2(n1012), .I3(GND_net), .O(n1067));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i678_3_lut (.I0(n990), .I1(n1043), 
            .I2(n1012), .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i674_3_lut (.I0(n986), .I1(n1039), 
            .I2(n1012), .I3(GND_net), .O(n1064));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i675_3_lut (.I0(n987), .I1(n1040), 
            .I2(n1012), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i682_3_lut (.I0(n994), .I1(n1047), 
            .I2(n1012), .I3(GND_net), .O(n1072));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_687_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4875));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_i680_3_lut (.I0(n992), .I1(n1045), 
            .I2(n1012), .I3(GND_net), .O(n1070));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_615_7_lut (.I0(duty[5]), .I1(n35425), .I2(n20_adj_4797), 
            .I3(n25589), .O(pwm_setpoint_22__N_3[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_i681_3_lut (.I0(n993), .I1(n1046), 
            .I2(n1012), .I3(GND_net), .O(n1071));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i622_3_lut (.I0(n909), .I1(n962), 
            .I2(n934), .I3(GND_net), .O(n987));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i621_3_lut (.I0(n908), .I1(n961), 
            .I2(n934), .I3(GND_net), .O(n986));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i626_3_lut (.I0(n913), .I1(n966), 
            .I2(n934), .I3(GND_net), .O(n991));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i627_3_lut (.I0(n914), .I1(n967), 
            .I2(n934), .I3(GND_net), .O(n992));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i627_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i625_3_lut (.I0(n912), .I1(n965), 
            .I2(n934), .I3(GND_net), .O(n990));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i623_3_lut (.I0(n910), .I1(n963), 
            .I2(n934), .I3(GND_net), .O(n988));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_884_16_lut (.I0(GND_net), .I1(n1298), 
            .I2(VCC_net), .I3(n25958), .O(n1351)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i624_3_lut (.I0(n911), .I1(n964), 
            .I2(n934), .I3(GND_net), .O(n989));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i624_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i570_3_lut (.I0(n832), .I1(n885), 
            .I2(n856), .I3(GND_net), .O(n910));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i569_3_lut (.I0(n831), .I1(n884), 
            .I2(n856), .I3(GND_net), .O(n909));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_884_15_lut (.I0(GND_net), .I1(n1299), 
            .I2(VCC_net), .I3(n25957), .O(n1352)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_687_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4879));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_i571_3_lut (.I0(n833), .I1(n886), 
            .I2(n856), .I3(GND_net), .O(n911));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i571_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_884_15 (.CI(n25957), .I0(n1299), 
            .I1(VCC_net), .CO(n25958));
    SB_LUT4 encoder0_position_23__I_0_i572_3_lut (.I0(n834), .I1(n887), 
            .I2(n856), .I3(GND_net), .O(n912));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_884_14_lut (.I0(GND_net), .I1(n1300), 
            .I2(VCC_net), .I3(n25956), .O(n1353)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i568_3_lut (.I0(n830), .I1(n883), 
            .I2(n856), .I3(GND_net), .O(n908));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i573_3_lut (.I0(n835), .I1(n888), 
            .I2(n856), .I3(GND_net), .O(n913));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i516_3_lut (.I0(n753), .I1(n806), 
            .I2(n778), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i27955_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n34127));
    defparam i27955_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_23__I_0_i517_3_lut (.I0(n754), .I1(n807), 
            .I2(n778), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i520_3_lut (.I0(n757), .I1(n810), 
            .I2(n778), .I3(GND_net), .O(n835));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i518_3_lut (.I0(n755), .I1(n808), 
            .I2(n778), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i518_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_884_14 (.CI(n25956), .I0(n1300), 
            .I1(VCC_net), .CO(n25957));
    SB_LUT4 encoder0_position_23__I_0_i519_3_lut (.I0(n756), .I1(n809), 
            .I2(n778), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_884_13_lut (.I0(GND_net), .I1(n1301), 
            .I2(VCC_net), .I3(n25955), .O(n1354)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i522_3_lut (.I0(n516), .I1(n812), 
            .I2(n778), .I3(GND_net), .O(n837));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i522_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_884_13 (.CI(n25955), .I0(n1301), 
            .I1(VCC_net), .CO(n25956));
    SB_LUT4 encoder0_position_23__I_0_add_884_12_lut (.I0(GND_net), .I1(n1302), 
            .I2(VCC_net), .I3(n25954), .O(n1355)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_12 (.CI(n25954), .I0(n1302), 
            .I1(VCC_net), .CO(n25955));
    SB_LUT4 encoder0_position_23__I_0_add_884_11_lut (.I0(GND_net), .I1(n1303), 
            .I2(VCC_net), .I3(n25953), .O(n1356)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_11 (.CI(n25953), .I0(n1303), 
            .I1(VCC_net), .CO(n25954));
    SB_LUT4 encoder0_position_23__I_0_add_884_10_lut (.I0(GND_net), .I1(n1304), 
            .I2(VCC_net), .I3(n25952), .O(n1357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_10 (.CI(n25952), .I0(n1304), 
            .I1(VCC_net), .CO(n25953));
    SB_LUT4 encoder0_position_23__I_0_i521_3_lut (.I0(n758), .I1(n811), 
            .I2(n778), .I3(GND_net), .O(n836));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_884_9_lut (.I0(GND_net), .I1(n1305), 
            .I2(VCC_net), .I3(n25951), .O(n1358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_9 (.CI(n25951), .I0(n1305), 
            .I1(VCC_net), .CO(n25952));
    SB_LUT4 encoder0_position_23__I_0_add_884_8_lut (.I0(GND_net), .I1(n1306), 
            .I2(VCC_net), .I3(n25950), .O(n1359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_687_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4881));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_884_8 (.CI(n25950), .I0(n1306), 
            .I1(VCC_net), .CO(n25951));
    SB_LUT4 i18181_3_lut (.I0(n517), .I1(n836), .I2(n837), .I3(GND_net), 
            .O(n22757));
    defparam i18181_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1643 (.I0(n834), .I1(n833), .I2(n22757), .I3(n835), 
            .O(n32355));
    defparam i2_4_lut_adj_1643.LUT_INIT = 16'h8880;
    SB_LUT4 encoder0_position_23__I_0_add_884_7_lut (.I0(GND_net), .I1(n1307), 
            .I2(GND_net), .I3(n25949), .O(n1360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28933_4_lut (.I0(n32355), .I1(n830), .I2(n832), .I3(n831), 
            .O(n856));
    defparam i28933_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_23__I_0_add_884_7 (.CI(n25949), .I0(n1307), 
            .I1(GND_net), .CO(n25950));
    SB_LUT4 mux_3158_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4827), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i576_3_lut (.I0(n517), .I1(n891), 
            .I2(n856), .I3(GND_net), .O(n916));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i575_3_lut (.I0(n837), .I1(n890), 
            .I2(n856), .I3(GND_net), .O(n915));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_687_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4877));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_i574_3_lut (.I0(n836), .I1(n889), 
            .I2(n856), .I3(GND_net), .O(n914));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18357_4_lut (.I0(n518), .I1(n914), .I2(n915), .I3(n916), 
            .O(n22937));
    defparam i18357_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1644 (.I0(n913), .I1(n908), .I2(n912), .I3(n22937), 
            .O(n7_adj_4850));
    defparam i2_4_lut_adj_1644.LUT_INIT = 16'heccc;
    SB_LUT4 i28949_4_lut (.I0(n7_adj_4850), .I1(n911), .I2(n909), .I3(n910), 
            .O(n934));
    defparam i28949_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i27970_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n34142));
    defparam i27970_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 encoder0_position_23__I_0_add_884_6_lut (.I0(GND_net), .I1(n1308), 
            .I2(GND_net), .I3(n25948), .O(n1361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_6 (.CI(n25948), .I0(n1308), 
            .I1(GND_net), .CO(n25949));
    SB_LUT4 encoder0_position_23__I_0_add_884_5_lut (.I0(GND_net), .I1(n1309), 
            .I2(VCC_net), .I3(n25947), .O(n1362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_5 (.CI(n25947), .I0(n1309), 
            .I1(VCC_net), .CO(n25948));
    SB_CARRY add_615_7 (.CI(n25589), .I0(n35425), .I1(n20_adj_4797), .CO(n25590));
    SB_LUT4 encoder0_position_23__I_0_add_884_4_lut (.I0(GND_net), .I1(n1310), 
            .I2(GND_net), .I3(n25946), .O(n1363)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_4 (.CI(n25946), .I0(n1310), 
            .I1(GND_net), .CO(n25947));
    SB_LUT4 encoder0_position_23__I_0_add_884_3_lut (.I0(GND_net), .I1(n1311), 
            .I2(VCC_net), .I3(n25945), .O(n1364)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_3 (.CI(n25945), .I0(n1311), 
            .I1(VCC_net), .CO(n25946));
    SB_LUT4 encoder0_position_23__I_0_add_884_2_lut (.I0(GND_net), .I1(n922), 
            .I2(GND_net), .I3(VCC_net), .O(n1365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3158_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4785), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_2 (.CI(VCC_net), .I0(n922), 
            .I1(GND_net), .CO(n25945));
    SB_LUT4 encoder0_position_23__I_0_add_831_15_lut (.I0(GND_net), .I1(n1220), 
            .I2(VCC_net), .I3(n25944), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_831_14_lut (.I0(GND_net), .I1(n1221), 
            .I2(VCC_net), .I3(n25943), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_14 (.CI(n25943), .I0(n1221), 
            .I1(VCC_net), .CO(n25944));
    SB_LUT4 encoder0_position_23__I_0_add_831_13_lut (.I0(GND_net), .I1(n1222), 
            .I2(VCC_net), .I3(n25942), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_13 (.CI(n25942), .I0(n1222), 
            .I1(VCC_net), .CO(n25943));
    SB_LUT4 encoder0_position_23__I_0_add_831_12_lut (.I0(GND_net), .I1(n1223), 
            .I2(VCC_net), .I3(n25941), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_12 (.CI(n25941), .I0(n1223), 
            .I1(VCC_net), .CO(n25942));
    SB_LUT4 encoder0_position_23__I_0_add_831_11_lut (.I0(GND_net), .I1(n1224), 
            .I2(VCC_net), .I3(n25940), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_11 (.CI(n25940), .I0(n1224), 
            .I1(VCC_net), .CO(n25941));
    SB_LUT4 encoder0_position_23__I_0_i630_3_lut (.I0(n518), .I1(n970), 
            .I2(n934), .I3(GND_net), .O(n995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_831_10_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n25939), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_10 (.CI(n25939), .I0(n1225), 
            .I1(VCC_net), .CO(n25940));
    SB_LUT4 encoder0_position_23__I_0_i629_3_lut (.I0(n916), .I1(n969), 
            .I2(n934), .I3(GND_net), .O(n994));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i628_3_lut (.I0(n915), .I1(n968), 
            .I2(n934), .I3(GND_net), .O(n993));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i628_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18353_4_lut (.I0(n519), .I1(n993), .I2(n994), .I3(n995), 
            .O(n22933));
    defparam i18353_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_2_lut_adj_1645 (.I0(n989), .I1(n988), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4871));
    defparam i2_2_lut_adj_1645.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n990), .I1(n992), .I2(n991), .I3(n22933), 
            .O(n7_adj_4872));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'heaaa;
    SB_LUT4 i28967_4_lut (.I0(n986), .I1(n7_adj_4872), .I2(n987), .I3(n8_adj_4871), 
            .O(n1012));
    defparam i28967_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4849), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i684_3_lut (.I0(n519), .I1(n1049), 
            .I2(n1012), .I3(GND_net), .O(n1074));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i683_3_lut (.I0(n995), .I1(n1048), 
            .I2(n1012), .I3(GND_net), .O(n1073));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18168_3_lut (.I0(n433), .I1(n1073), .I2(n1074), .I3(GND_net), 
            .O(n22743));
    defparam i18168_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1647 (.I0(n1071), .I1(n1070), .I2(n22743), .I3(n1072), 
            .O(n31767));
    defparam i2_4_lut_adj_1647.LUT_INIT = 16'h8880;
    SB_LUT4 i5_4_lut_adj_1648 (.I0(n1065), .I1(n1064), .I2(n31767), .I3(n1068), 
            .O(n12_adj_4870));
    defparam i5_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i28983_4_lut (.I0(n1067), .I1(n12_adj_4870), .I2(n1066), .I3(n1069), 
            .O(n1090));
    defparam i28983_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4848), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n433));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i738_3_lut (.I0(n433), .I1(n1128), 
            .I2(n1090), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5007[1]), .I1(r_SM_Main_adj_5007[0]), 
            .I2(r_SM_Main_adj_5007[2]), .I3(r_SM_Main_2__N_3404[1]), .O(n35944));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 encoder0_position_23__I_0_i737_3_lut (.I0(n1074), .I1(n1127), 
            .I2(n1090), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i736_3_lut (.I0(n1073), .I1(n1126), 
            .I2(n1090), .I3(GND_net), .O(n1151));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18347_4_lut (.I0(n434), .I1(n1151), .I2(n1152), .I3(n1153), 
            .O(n22927));
    defparam i18347_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i6_4_lut_adj_1649 (.I0(n1146), .I1(n1148), .I2(n1144), .I3(n1147), 
            .O(n14_adj_4811));
    defparam i6_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n1150), .I1(n1145), .I2(n1149), .I3(n22927), 
            .O(n9_adj_4812));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'heccc;
    SB_LUT4 i29008_4_lut (.I0(n9_adj_4812), .I1(n14_adj_4811), .I2(n1142), 
            .I3(n1143), .O(n1168));
    defparam i29008_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4820), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n434));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i792_3_lut (.I0(n434), .I1(n1207), 
            .I2(n1168), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i791_3_lut (.I0(n1153), .I1(n1206), 
            .I2(n1168), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i790_3_lut (.I0(n1152), .I1(n1205), 
            .I2(n1168), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3158_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4847), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n435));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18345_4_lut (.I0(n435), .I1(n1230), .I2(n1231), .I3(n1232), 
            .O(n22925));
    defparam i18345_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i13690_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n32812), .I3(GND_net), .O(n18270));   // verilog/coms.v(127[12] 300[6])
    defparam i13690_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1651 (.I0(n1223), .I1(n1224), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4806));
    defparam i1_2_lut_adj_1651.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1652 (.I0(n1229), .I1(n1222), .I2(n1228), .I3(n22925), 
            .O(n12_adj_4805));
    defparam i3_4_lut_adj_1652.LUT_INIT = 16'heccc;
    SB_LUT4 i13691_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n32812), .I3(GND_net), .O(n18271));   // verilog/coms.v(127[12] 300[6])
    defparam i13691_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1653 (.I0(n1225), .I1(n1227), .I2(n1221), .I3(n10_adj_4806), 
            .O(n16_adj_4804));
    defparam i7_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i29109_4_lut (.I0(n1226), .I1(n16_adj_4804), .I2(n12_adj_4805), 
            .I3(n1220), .O(n1246));
    defparam i29109_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i785_3_lut (.I0(n1147), .I1(n1200), 
            .I2(n1168), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13692_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n32812), .I3(GND_net), .O(n18272));   // verilog/coms.v(127[12] 300[6])
    defparam i13692_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i838_3_lut (.I0(n1225), .I1(n1278), 
            .I2(n1246), .I3(GND_net), .O(n1303));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i841_3_lut (.I0(n1228), .I1(n1281), 
            .I2(n1246), .I3(GND_net), .O(n1306));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18339_3_lut (.I0(n922), .I1(n1310), .I2(n1311), .I3(GND_net), 
            .O(n22919));
    defparam i18339_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1654 (.I0(n1308), .I1(n1307), .I2(n22919), .I3(n1309), 
            .O(n32929));
    defparam i2_4_lut_adj_1654.LUT_INIT = 16'h8880;
    SB_LUT4 i13693_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n32812), .I3(GND_net), .O(n18273));   // verilog/coms.v(127[12] 300[6])
    defparam i13693_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1655 (.I0(n1300), .I1(n32929), .I2(n1306), .I3(n1303), 
            .O(n16_adj_4803));
    defparam i6_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i13694_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n32812), .I3(GND_net), .O(n18274));   // verilog/coms.v(127[12] 300[6])
    defparam i13694_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1656 (.I0(n1301), .I1(n1298), .I2(n1299), .I3(n1304), 
            .O(n17_adj_4802));
    defparam i7_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i29027_4_lut (.I0(n17_adj_4802), .I1(n1302), .I2(n16_adj_4803), 
            .I3(n1305), .O(n1324));
    defparam i29027_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i835_3_lut (.I0(n1222), .I1(n1275), 
            .I2(n1246), .I3(GND_net), .O(n1300));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i888_3_lut (.I0(n1300), .I1(n1353), 
            .I2(n1324), .I3(GND_net), .O(n1378));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13695_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n32812), .I3(GND_net), .O(n18275));   // verilog/coms.v(127[12] 300[6])
    defparam i13695_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i894_3_lut (.I0(n1306), .I1(n1359), 
            .I2(n1324), .I3(GND_net), .O(n1384));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i889_3_lut (.I0(n1301), .I1(n1354), 
            .I2(n1324), .I3(GND_net), .O(n1379));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13696_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n32812), .I3(GND_net), .O(n18276));   // verilog/coms.v(127[12] 300[6])
    defparam i13696_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18336_3_lut (.I0(n923), .I1(n1389), .I2(n1390), .I3(GND_net), 
            .O(n22915));
    defparam i18336_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1657 (.I0(n1387), .I1(n1386), .I2(n22915), .I3(n1388), 
            .O(n32238));
    defparam i2_4_lut_adj_1657.LUT_INIT = 16'h8880;
    SB_LUT4 i13697_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n32812), .I3(GND_net), .O(n18277));   // verilog/coms.v(127[12] 300[6])
    defparam i13697_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1658 (.I0(n1383), .I1(n1380), .I2(n1377), .I3(n32238), 
            .O(n18_adj_4937));
    defparam i7_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1385), .I1(n1381), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4938));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13698_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n32812), .I3(GND_net), .O(n18278));   // verilog/coms.v(127[12] 300[6])
    defparam i13698_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_4_lut_adj_1659 (.I0(n1379), .I1(n18_adj_4937), .I2(n1384), 
            .I3(n1378), .O(n20_adj_4936));
    defparam i9_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i13699_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n32812), .I3(GND_net), .O(n18279));   // verilog/coms.v(127[12] 300[6])
    defparam i13699_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29070_4_lut (.I0(n1376), .I1(n20_adj_4936), .I2(n16_adj_4938), 
            .I3(n1382), .O(n1402));
    defparam i29070_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4841), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i954_3_lut (.I0(n923), .I1(n1444), 
            .I2(n1402), .I3(GND_net), .O(n1469));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i953_3_lut (.I0(n1390), .I1(n1443), 
            .I2(n1402), .I3(GND_net), .O(n1468));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13700_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n32812), .I3(GND_net), .O(n18280));   // verilog/coms.v(127[12] 300[6])
    defparam i13700_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i952_3_lut (.I0(n1389), .I1(n1442), 
            .I2(n1402), .I3(GND_net), .O(n1467));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18430_4_lut (.I0(n924), .I1(n1467), .I2(n1468), .I3(n1469), 
            .O(n23011));
    defparam i18430_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i8_4_lut_adj_1660 (.I0(n1464), .I1(n1458), .I2(n1463), .I3(n1456), 
            .O(n20_adj_4818));
    defparam i8_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1661 (.I0(n1457), .I1(n1466), .I2(n1465), .I3(n23011), 
            .O(n13_adj_4821));
    defparam i1_4_lut_adj_1661.LUT_INIT = 16'heaaa;
    SB_LUT4 i13701_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n32812), .I3(GND_net), .O(n18281));   // verilog/coms.v(127[12] 300[6])
    defparam i13701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13702_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n32812), .I3(GND_net), .O(n18282));   // verilog/coms.v(127[12] 300[6])
    defparam i13702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13703_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n32812), .I3(GND_net), .O(n18283));   // verilog/coms.v(127[12] 300[6])
    defparam i13703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_2_lut (.I0(n1461), .I1(n1459), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4819));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_add_831_9_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n25938), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_9 (.CI(n25938), .I0(n1226), 
            .I1(VCC_net), .CO(n25939));
    SB_LUT4 i10_4_lut_adj_1662 (.I0(n13_adj_4821), .I1(n20_adj_4818), .I2(n1460), 
            .I3(n1454), .O(n22_adj_4817));
    defparam i10_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_831_8_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n25937), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_6_lut (.I0(duty[4]), .I1(n35425), .I2(n21_adj_4798), 
            .I3(n25588), .O(pwm_setpoint_22__N_3[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_831_8 (.CI(n25937), .I0(n1227), 
            .I1(VCC_net), .CO(n25938));
    SB_LUT4 i29091_4_lut (.I0(n1462), .I1(n22_adj_4817), .I2(n18_adj_4819), 
            .I3(n1455), .O(n1480));
    defparam i29091_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_add_831_7_lut (.I0(GND_net), .I1(n1228), 
            .I2(GND_net), .I3(n25936), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_7 (.CI(n25936), .I0(n1228), 
            .I1(GND_net), .CO(n25937));
    SB_LUT4 encoder0_position_23__I_0_add_831_6_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n25935), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_6 (.CI(n25935), .I0(n1229), 
            .I1(GND_net), .CO(n25936));
    SB_LUT4 encoder0_position_23__I_0_add_831_5_lut (.I0(GND_net), .I1(n1230), 
            .I2(VCC_net), .I3(n25934), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_5 (.CI(n25934), .I0(n1230), 
            .I1(VCC_net), .CO(n25935));
    SB_LUT4 encoder0_position_23__I_0_add_831_4_lut (.I0(GND_net), .I1(n1231), 
            .I2(GND_net), .I3(n25933), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_4 (.CI(n25933), .I0(n1231), 
            .I1(GND_net), .CO(n25934));
    SB_LUT4 mux_3158_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4836), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13704_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n32812), .I3(GND_net), .O(n18284));   // verilog/coms.v(127[12] 300[6])
    defparam i13704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1008_3_lut (.I0(n924), .I1(n1523), 
            .I2(n1480), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1007_3_lut (.I0(n1469), .I1(n1522), 
            .I2(n1480), .I3(GND_net), .O(n1547));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_831_3_lut (.I0(GND_net), .I1(n1232), 
            .I2(VCC_net), .I3(n25932), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_6 (.CI(n25588), .I0(n35425), .I1(n21_adj_4798), .CO(n25589));
    SB_CARRY encoder0_position_23__I_0_add_831_3 (.CI(n25932), .I0(n1232), 
            .I1(VCC_net), .CO(n25933));
    SB_LUT4 encoder0_position_23__I_0_add_831_2_lut (.I0(GND_net), .I1(n435), 
            .I2(GND_net), .I3(VCC_net), .O(n1286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_2 (.CI(VCC_net), .I0(n435), 
            .I1(GND_net), .CO(n25932));
    SB_LUT4 encoder0_position_23__I_0_add_778_14_lut (.I0(GND_net), .I1(n1142), 
            .I2(VCC_net), .I3(n25931), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13705_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n32812), .I3(GND_net), .O(n18285));   // verilog/coms.v(127[12] 300[6])
    defparam i13705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_13_lut (.I0(GND_net), .I1(n1143), 
            .I2(VCC_net), .I3(n25930), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_13 (.CI(n25930), .I0(n1143), 
            .I1(VCC_net), .CO(n25931));
    SB_LUT4 encoder0_position_23__I_0_add_778_12_lut (.I0(GND_net), .I1(n1144), 
            .I2(VCC_net), .I3(n25929), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_12 (.CI(n25929), .I0(n1144), 
            .I1(VCC_net), .CO(n25930));
    SB_LUT4 encoder0_position_23__I_0_add_778_11_lut (.I0(GND_net), .I1(n1145), 
            .I2(VCC_net), .I3(n25928), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_11 (.CI(n25928), .I0(n1145), 
            .I1(VCC_net), .CO(n25929));
    SB_LUT4 encoder0_position_23__I_0_add_778_10_lut (.I0(GND_net), .I1(n1146), 
            .I2(VCC_net), .I3(n25927), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_10 (.CI(n25927), .I0(n1146), 
            .I1(VCC_net), .CO(n25928));
    SB_LUT4 encoder0_position_23__I_0_add_778_9_lut (.I0(GND_net), .I1(n1147), 
            .I2(VCC_net), .I3(n25926), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_9 (.CI(n25926), .I0(n1147), 
            .I1(VCC_net), .CO(n25927));
    SB_LUT4 encoder0_position_23__I_0_add_778_8_lut (.I0(GND_net), .I1(n1148), 
            .I2(VCC_net), .I3(n25925), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_8 (.CI(n25925), .I0(n1148), 
            .I1(VCC_net), .CO(n25926));
    SB_LUT4 encoder0_position_23__I_0_add_778_7_lut (.I0(GND_net), .I1(n1149), 
            .I2(GND_net), .I3(n25924), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_615_5_lut (.I0(duty[3]), .I1(n35425), .I2(n22), .I3(n25587), 
            .O(pwm_setpoint_22__N_3[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_778_7 (.CI(n25924), .I0(n1149), 
            .I1(GND_net), .CO(n25925));
    SB_LUT4 encoder0_position_23__I_0_add_778_6_lut (.I0(GND_net), .I1(n1150), 
            .I2(GND_net), .I3(n25923), .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_615_5 (.CI(n25587), .I0(n35425), .I1(n22), .CO(n25588));
    SB_CARRY encoder0_position_23__I_0_add_778_6 (.CI(n25923), .I0(n1150), 
            .I1(GND_net), .CO(n25924));
    SB_LUT4 encoder0_position_23__I_0_add_778_5_lut (.I0(GND_net), .I1(n1151), 
            .I2(VCC_net), .I3(n25922), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_5 (.CI(n25922), .I0(n1151), 
            .I1(VCC_net), .CO(n25923));
    SB_LUT4 add_615_4_lut (.I0(duty[2]), .I1(n35425), .I2(n23_adj_4799), 
            .I3(n25586), .O(pwm_setpoint_22__N_3[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_615_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_778_4_lut (.I0(GND_net), .I1(n1152), 
            .I2(GND_net), .I3(n25921), .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_4 (.CI(n25921), .I0(n1152), 
            .I1(GND_net), .CO(n25922));
    SB_LUT4 encoder0_position_23__I_0_add_778_3_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n25920), .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1006_3_lut (.I0(n1468), .I1(n1521), 
            .I2(n1480), .I3(GND_net), .O(n1546));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1006_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_778_3 (.CI(n25920), .I0(n1153), 
            .I1(VCC_net), .CO(n25921));
    SB_LUT4 encoder0_position_23__I_0_add_778_2_lut (.I0(GND_net), .I1(n434), 
            .I2(GND_net), .I3(VCC_net), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_2 (.CI(VCC_net), .I0(n434), 
            .I1(GND_net), .CO(n25920));
    SB_LUT4 encoder0_position_23__I_0_add_725_13_lut (.I0(GND_net), .I1(n1064), 
            .I2(VCC_net), .I3(n25919), .O(n1117)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_12_lut (.I0(GND_net), .I1(n1065), 
            .I2(VCC_net), .I3(n25918), .O(n1118)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_12 (.CI(n25918), .I0(n1065), 
            .I1(VCC_net), .CO(n25919));
    SB_LUT4 encoder0_position_23__I_0_add_725_11_lut (.I0(GND_net), .I1(n1066), 
            .I2(VCC_net), .I3(n25917), .O(n1119)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_11 (.CI(n25917), .I0(n1066), 
            .I1(VCC_net), .CO(n25918));
    SB_LUT4 encoder0_position_23__I_0_add_725_10_lut (.I0(GND_net), .I1(n1067), 
            .I2(VCC_net), .I3(n25916), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_10 (.CI(n25916), .I0(n1067), 
            .I1(VCC_net), .CO(n25917));
    SB_LUT4 add_1733_7_lut (.I0(GND_net), .I1(n509), .I2(GND_net), .I3(n25654), 
            .O(n5273)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_9_lut (.I0(GND_net), .I1(n1068), 
            .I2(VCC_net), .I3(n25915), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_9 (.CI(n25915), .I0(n1068), 
            .I1(VCC_net), .CO(n25916));
    SB_LUT4 i18426_4_lut (.I0(n925), .I1(n1546), .I2(n1547), .I3(n1548), 
            .O(n23007));
    defparam i18426_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1663 (.I0(n1545), .I1(n1534), .I2(n1544), .I3(n23007), 
            .O(n17_adj_4933));
    defparam i4_4_lut_adj_1663.LUT_INIT = 16'heccc;
    SB_LUT4 i8_4_lut_adj_1664 (.I0(n1533), .I1(n1542), .I2(n1538), .I3(n1540), 
            .O(n21_adj_4930));
    defparam i8_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1539), .I1(n1536), .I2(n1543), .I3(GND_net), 
            .O(n20_adj_4931));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13706_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n32812), .I3(GND_net), .O(n18286));   // verilog/coms.v(127[12] 300[6])
    defparam i13706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13707_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n32812), .I3(GND_net), .O(n18287));   // verilog/coms.v(127[12] 300[6])
    defparam i13707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_1665 (.I0(n21_adj_4930), .I1(n17_adj_4933), .I2(n1537), 
            .I3(n1532), .O(n24_adj_4929));
    defparam i11_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 i13708_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n32812), .I3(GND_net), .O(n18288));   // verilog/coms.v(127[12] 300[6])
    defparam i13708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28917_4_lut (.I0(n1535), .I1(n24_adj_4929), .I2(n20_adj_4931), 
            .I3(n1541), .O(n1558));
    defparam i28917_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_725_8_lut (.I0(GND_net), .I1(n1069), 
            .I2(VCC_net), .I3(n25914), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13709_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n32812), .I3(GND_net), .O(n18289));   // verilog/coms.v(127[12] 300[6])
    defparam i13709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1062_3_lut (.I0(n925), .I1(n1602), 
            .I2(n1558), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1061_3_lut (.I0(n1548), .I1(n1601), 
            .I2(n1558), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13710_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n32812), .I3(GND_net), .O(n18290));   // verilog/coms.v(127[12] 300[6])
    defparam i13710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3158_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18324_3_lut (.I0(n926), .I1(n1626), .I2(n1627), .I3(GND_net), 
            .O(n22903));
    defparam i18324_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1666 (.I0(n1624), .I1(n1623), .I2(n22903), .I3(n1625), 
            .O(n32337));
    defparam i2_4_lut_adj_1666.LUT_INIT = 16'h8880;
    SB_LUT4 i13711_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n32812), .I3(GND_net), .O(n18291));   // verilog/coms.v(127[12] 300[6])
    defparam i13711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_2_lut (.I0(n1618), .I1(n1613), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4826));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1667 (.I0(n1614), .I1(n1612), .I2(n1615), .I3(n1617), 
            .O(n24_adj_4824));
    defparam i10_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_23__I_0_add_725_8 (.CI(n25914), .I0(n1069), 
            .I1(VCC_net), .CO(n25915));
    SB_LUT4 i8_4_lut_adj_1668 (.I0(n1610), .I1(n1622), .I2(n1620), .I3(n32337), 
            .O(n22_adj_4825));
    defparam i8_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1669 (.I0(n1616), .I1(n24_adj_4824), .I2(n18_adj_4826), 
            .I3(n1611), .O(n26));
    defparam i12_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_725_7_lut (.I0(GND_net), .I1(n1070), 
            .I2(GND_net), .I3(n25913), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13712_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n32812), .I3(GND_net), .O(n18292));   // verilog/coms.v(127[12] 300[6])
    defparam i13712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29050_4_lut (.I0(n1621), .I1(n26), .I2(n22_adj_4825), .I3(n1619), 
            .O(n1636));
    defparam i29050_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i13460_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18040));   // verilog/coms.v(127[12] 300[6])
    defparam i13460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1059_3_lut (.I0(n1546), .I1(n1599), 
            .I2(n1558), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1112_3_lut (.I0(n1624), .I1(n1677), 
            .I2(n1636), .I3(GND_net), .O(n1702));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1113_3_lut (.I0(n1625), .I1(n1678), 
            .I2(n1636), .I3(GND_net), .O(n1703));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1110_3_lut (.I0(n1622), .I1(n1675), 
            .I2(n1636), .I3(GND_net), .O(n1700));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13462_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n21943), 
            .I3(n16544), .O(n18042));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13462_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_23__I_0_add_725_7 (.CI(n25913), .I0(n1070), 
            .I1(GND_net), .CO(n25914));
    SB_LUT4 encoder0_position_23__I_0_add_725_6_lut (.I0(GND_net), .I1(n1071), 
            .I2(GND_net), .I3(n25912), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_6 (.CI(n25912), .I0(n1071), 
            .I1(GND_net), .CO(n25913));
    SB_LUT4 encoder0_position_23__I_0_add_725_5_lut (.I0(GND_net), .I1(n1072), 
            .I2(VCC_net), .I3(n25911), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_5 (.CI(n25911), .I0(n1072), 
            .I1(VCC_net), .CO(n25912));
    SB_LUT4 i18420_4_lut (.I0(n927), .I1(n1704), .I2(n1705), .I3(n1706), 
            .O(n23001));
    defparam i18420_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i11_4_lut_adj_1670 (.I0(n1688), .I1(n1695), .I2(n1692), .I3(n1701), 
            .O(n26_adj_4944));
    defparam i11_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 i13463_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n21943), 
            .I3(n16549), .O(n18043));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13463_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i4_4_lut_adj_1671 (.I0(n1700), .I1(n1703), .I2(n1702), .I3(n23001), 
            .O(n19_adj_4946));
    defparam i4_4_lut_adj_1671.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1672 (.I0(n1698), .I1(n1693), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4947));
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1673 (.I0(n1697), .I1(n1694), .I2(n1691), .I3(n1689), 
            .O(n24_adj_4945));
    defparam i9_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1674 (.I0(n19_adj_4946), .I1(n26_adj_4944), .I2(n1690), 
            .I3(n1696), .O(n28_adj_4943));
    defparam i13_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i13464_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4846), 
            .I3(n16544), .O(n18044));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13464_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29133_4_lut (.I0(n1699), .I1(n28_adj_4943), .I2(n24_adj_4945), 
            .I3(n16_adj_4947), .O(n1714));
    defparam i29133_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3158_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n927));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13465_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4846), 
            .I3(n16549), .O(n18045));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13465_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13466_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4840), 
            .I3(n16544), .O(n18046));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13466_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1170_3_lut (.I0(n927), .I1(n1760), 
            .I2(n1714), .I3(GND_net), .O(n1785));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1169_3_lut (.I0(n1706), .I1(n1759), 
            .I2(n1714), .I3(GND_net), .O(n1784));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18316_3_lut (.I0(n928), .I1(n1784), .I2(n1785), .I3(GND_net), 
            .O(n22895));
    defparam i18316_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1675 (.I0(n1782), .I1(n1781), .I2(n22895), .I3(n1783), 
            .O(n32029));
    defparam i2_4_lut_adj_1675.LUT_INIT = 16'h8880;
    SB_LUT4 i12_4_lut_adj_1676 (.I0(n1772), .I1(n1767), .I2(n1775), .I3(n1779), 
            .O(n28_adj_4894));
    defparam i12_4_lut_adj_1676.LUT_INIT = 16'hfffe;
    SB_LUT4 i13467_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4840), 
            .I3(n16549), .O(n18047));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13467_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10_4_lut_adj_1677 (.I0(n1770), .I1(n1773), .I2(n1766), .I3(n1771), 
            .O(n26_adj_4896));
    defparam i10_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i13713_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n13933), .I3(GND_net), .O(n18293));   // verilog/coms.v(127[12] 300[6])
    defparam i13713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1678 (.I0(n1778), .I1(n1777), .I2(n1774), .I3(n1768), 
            .O(n27_adj_4895));
    defparam i11_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 i13714_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n13933), .I3(GND_net), .O(n18294));   // verilog/coms.v(127[12] 300[6])
    defparam i13714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13715_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n13933), .I3(GND_net), .O(n18295));   // verilog/coms.v(127[12] 300[6])
    defparam i13715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1679 (.I0(n32029), .I1(n1776), .I2(n1769), .I3(n1780), 
            .O(n25_adj_4897));
    defparam i9_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 i29158_4_lut (.I0(n25_adj_4897), .I1(n27_adj_4895), .I2(n26_adj_4896), 
            .I3(n28_adj_4894), .O(n1792));
    defparam i29158_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i13716_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n13933), .I3(GND_net), .O(n18296));   // verilog/coms.v(127[12] 300[6])
    defparam i13716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3158_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4843), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1224_3_lut (.I0(n928), .I1(n1839), 
            .I2(n1792), .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1224_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1223_3_lut (.I0(n1785), .I1(n1838), 
            .I2(n1792), .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3158_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1680 (.I0(n1851), .I1(n1848), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4815));
    defparam i1_2_lut_adj_1680.LUT_INIT = 16'heeee;
    SB_LUT4 i18314_3_lut (.I0(n929), .I1(n1863), .I2(n1864), .I3(GND_net), 
            .O(n22893));
    defparam i18314_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1681 (.I0(n1861), .I1(n1860), .I2(n22893), .I3(n1862), 
            .O(n32360));
    defparam i2_4_lut_adj_1681.LUT_INIT = 16'h8880;
    SB_LUT4 i13_4_lut_adj_1682 (.I0(n1844), .I1(n1859), .I2(n1847), .I3(n18_adj_4815), 
            .O(n30_adj_4813));
    defparam i13_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1683 (.I0(n1852), .I1(n32360), .I2(n1845), .I3(n1850), 
            .O(n28_adj_4814));
    defparam i11_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i13717_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n13933), .I3(GND_net), .O(n18297));   // verilog/coms.v(127[12] 300[6])
    defparam i13717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13718_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n13933), .I3(GND_net), .O(n18298));   // verilog/coms.v(127[12] 300[6])
    defparam i13718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1684 (.I0(n1856), .I1(n1849), .I2(n1846), .I3(n1853), 
            .O(n29));
    defparam i12_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1685 (.I0(n1854), .I1(n1858), .I2(n1855), .I3(n1857), 
            .O(n27));
    defparam i10_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i29184_4_lut (.I0(n27), .I1(n29), .I2(n28_adj_4814), .I3(n30_adj_4813), 
            .O(n1870));
    defparam i29184_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i13719_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n13933), .I3(GND_net), .O(n18299));   // verilog/coms.v(127[12] 300[6])
    defparam i13719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1219_3_lut (.I0(n1781), .I1(n1834), 
            .I2(n1792), .I3(GND_net), .O(n1859));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1263_3_lut (.I0(n1850), .I1(n1903), 
            .I2(n1870), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1272_3_lut (.I0(n1859), .I1(n1912), 
            .I2(n1870), .I3(GND_net), .O(n1937));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1267_3_lut (.I0(n1854), .I1(n1907), 
            .I2(n1870), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13468_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4), .I3(n16544), 
            .O(n18048));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13468_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13469_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18049));   // verilog/coms.v(127[12] 300[6])
    defparam i13469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13470_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n32040), 
            .I3(GND_net), .O(n18050));   // verilog/coms.v(127[12] 300[6])
    defparam i13470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1260_3_lut (.I0(n1847), .I1(n1900), 
            .I2(n1870), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13471_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n32040), 
            .I3(GND_net), .O(n18051));   // verilog/coms.v(127[12] 300[6])
    defparam i13471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18408_4_lut (.I0(n930), .I1(n1941), .I2(n1942), .I3(n1943), 
            .O(n22989));
    defparam i18408_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i10_4_lut_adj_1686 (.I0(n1925), .I1(n1932), .I2(n1937), .I3(n1928), 
            .O(n28));
    defparam i10_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1687 (.I0(n1923), .I1(n1930), .I2(n1927), .I3(n1935), 
            .O(n31));
    defparam i13_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1688 (.I0(n1938), .I1(n1940), .I2(n1939), .I3(n22989), 
            .O(n22_adj_4800));
    defparam i4_4_lut_adj_1688.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut_adj_1689 (.I0(n1931), .I1(n1934), .I2(n1922), .I3(n1936), 
            .O(n30));
    defparam i12_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1690 (.I0(n31), .I1(n1924), .I2(n28), .I3(n1933), 
            .O(n34));
    defparam i16_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_LUT4 i13472_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n32812), .I3(GND_net), .O(n18052));   // verilog/coms.v(127[12] 300[6])
    defparam i13472_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_2_lut (.I0(n1926), .I1(n1929), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_4801));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29211_4_lut (.I0(n21_adj_4801), .I1(n34), .I2(n30), .I3(n22_adj_4800), 
            .O(n1948));
    defparam i29211_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n22632), 
            .I2(n16614), .I3(GND_net), .O(n63));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 encoder0_position_23__I_0_i1257_3_lut (.I0(n1844), .I1(n1897), 
            .I2(n1870), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1310_3_lut (.I0(n1922), .I1(n1975), 
            .I2(n1948), .I3(GND_net), .O(n2000));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_725_4_lut (.I0(GND_net), .I1(n1073), 
            .I2(GND_net), .I3(n25910), .O(n1126)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_4 (.CI(n25910), .I0(n1073), 
            .I1(GND_net), .CO(n25911));
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4790));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13720_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n13933), .I3(GND_net), .O(n18300));   // verilog/coms.v(127[12] 300[6])
    defparam i13720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13721_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n13933), .I3(GND_net), .O(n18301));   // verilog/coms.v(127[12] 300[6])
    defparam i13721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13722_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n13933), .I3(GND_net), .O(n18302));   // verilog/coms.v(127[12] 300[6])
    defparam i13722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13723_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n13933), .I3(GND_net), .O(n18303));   // verilog/coms.v(127[12] 300[6])
    defparam i13723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_725_3_lut (.I0(GND_net), .I1(n1074), 
            .I2(VCC_net), .I3(n25909), .O(n1127)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13724_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n13933), .I3(GND_net), .O(n18304));   // verilog/coms.v(127[12] 300[6])
    defparam i13724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13725_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n13933), .I3(GND_net), .O(n18305));   // verilog/coms.v(127[12] 300[6])
    defparam i13725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13726_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n13933), .I3(GND_net), .O(n18306));   // verilog/coms.v(127[12] 300[6])
    defparam i13726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13727_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n13933), .I3(GND_net), .O(n18307));   // verilog/coms.v(127[12] 300[6])
    defparam i13727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13728_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n13933), .I3(GND_net), .O(n18308));   // verilog/coms.v(127[12] 300[6])
    defparam i13728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13729_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n13933), .I3(GND_net), .O(n18309));   // verilog/coms.v(127[12] 300[6])
    defparam i13729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13730_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n13933), .I3(GND_net), .O(n18310));   // verilog/coms.v(127[12] 300[6])
    defparam i13730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13731_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n13933), .I3(GND_net), .O(n18311));   // verilog/coms.v(127[12] 300[6])
    defparam i13731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13732_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n13933), .I3(GND_net), .O(n18312));   // verilog/coms.v(127[12] 300[6])
    defparam i13732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13733_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n13933), .I3(GND_net), .O(n18313));   // verilog/coms.v(127[12] 300[6])
    defparam i13733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13734_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n13933), .I3(GND_net), .O(n18314));   // verilog/coms.v(127[12] 300[6])
    defparam i13734_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_725_3 (.CI(n25909), .I0(n1074), 
            .I1(VCC_net), .CO(n25910));
    SB_LUT4 encoder0_position_23__I_0_add_725_2_lut (.I0(GND_net), .I1(n433), 
            .I2(GND_net), .I3(VCC_net), .O(n1128)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13735_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n13933), .I3(GND_net), .O(n18315));   // verilog/coms.v(127[12] 300[6])
    defparam i13735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13736_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n13933), .I3(GND_net), .O(n18316));   // verilog/coms.v(127[12] 300[6])
    defparam i13736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4789));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13737_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13933), .I3(GND_net), .O(n18317));   // verilog/coms.v(127[12] 300[6])
    defparam i13737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1495_3_lut (.I0(n22965), .I1(n5522), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_26[0]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1495_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i28166_4_lut (.I0(n10_adj_4832), .I1(n21828), .I2(n21898), 
            .I3(state_7__N_3815[0]), .O(n34061));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i28166_4_lut.LUT_INIT = 16'hc8cc;
    SB_CARRY encoder0_position_23__I_0_add_725_2 (.CI(VCC_net), .I0(n433), 
            .I1(GND_net), .CO(n25909));
    SB_LUT4 i16_4_lut_adj_1691 (.I0(state_adj_5030[0]), .I1(n34061), .I2(n4604), 
            .I3(n21826), .O(n8_adj_4807));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i16_4_lut_adj_1691.LUT_INIT = 16'h3afa;
    SB_LUT4 i13743_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13933), .I3(GND_net), .O(n18323));   // verilog/coms.v(127[12] 300[6])
    defparam i13743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_672_12_lut (.I0(GND_net), .I1(n986), 
            .I2(VCC_net), .I3(n25908), .O(n1039)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_672_11_lut (.I0(GND_net), .I1(n987), 
            .I2(VCC_net), .I3(n25907), .O(n1040)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_11 (.CI(n25907), .I0(n987), 
            .I1(VCC_net), .CO(n25908));
    SB_LUT4 encoder0_position_23__I_0_add_672_10_lut (.I0(GND_net), .I1(n988), 
            .I2(VCC_net), .I3(n25906), .O(n1041)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_10 (.CI(n25906), .I0(n988), 
            .I1(VCC_net), .CO(n25907));
    SB_LUT4 encoder0_position_23__I_0_add_672_9_lut (.I0(GND_net), .I1(n989), 
            .I2(VCC_net), .I3(n25905), .O(n1042)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_9 (.CI(n25905), .I0(n989), 
            .I1(VCC_net), .CO(n25906));
    SB_LUT4 i13744_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13933), .I3(GND_net), .O(n18324));   // verilog/coms.v(127[12] 300[6])
    defparam i13744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_672_8_lut (.I0(GND_net), .I1(n990), 
            .I2(VCC_net), .I3(n25904), .O(n1043)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_8 (.CI(n25904), .I0(n990), 
            .I1(VCC_net), .CO(n25905));
    SB_LUT4 encoder0_position_23__I_0_add_672_7_lut (.I0(GND_net), .I1(n991), 
            .I2(GND_net), .I3(n25903), .O(n1044)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_7 (.CI(n25903), .I0(n991), 
            .I1(GND_net), .CO(n25904));
    SB_LUT4 encoder0_position_23__I_0_add_672_6_lut (.I0(GND_net), .I1(n992), 
            .I2(GND_net), .I3(n25902), .O(n1045)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_6 (.CI(n25902), .I0(n992), 
            .I1(GND_net), .CO(n25903));
    SB_LUT4 encoder0_position_23__I_0_add_672_5_lut (.I0(GND_net), .I1(n993), 
            .I2(VCC_net), .I3(n25901), .O(n1046)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13745_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13933), .I3(GND_net), .O(n18325));   // verilog/coms.v(127[12] 300[6])
    defparam i13745_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_672_5 (.CI(n25901), .I0(n993), 
            .I1(VCC_net), .CO(n25902));
    SB_LUT4 encoder0_position_23__I_0_add_672_4_lut (.I0(GND_net), .I1(n994), 
            .I2(GND_net), .I3(n25900), .O(n1047)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_4 (.CI(n25900), .I0(n994), 
            .I1(GND_net), .CO(n25901));
    SB_LUT4 encoder0_position_23__I_0_add_672_3_lut (.I0(GND_net), .I1(n995), 
            .I2(VCC_net), .I3(n25899), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_3 (.CI(n25899), .I0(n995), 
            .I1(VCC_net), .CO(n25900));
    SB_LUT4 encoder0_position_23__I_0_add_672_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n25899));
    SB_LUT4 i1_2_lut_adj_1692 (.I0(n16456), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n16458));
    defparam i1_2_lut_adj_1692.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_add_619_11_lut (.I0(GND_net), .I1(n908), 
            .I2(VCC_net), .I3(n25898), .O(n961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_619_10_lut (.I0(GND_net), .I1(n909), 
            .I2(VCC_net), .I3(n25897), .O(n962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27962_4_lut (.I0(n27_adj_4889), .I1(n15_adj_4883), .I2(n13_adj_4882), 
            .I3(n11_adj_4880), .O(n34134));
    defparam i27962_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_23__I_0_add_619_10 (.CI(n25897), .I0(n909), 
            .I1(VCC_net), .CO(n25898));
    SB_LUT4 encoder0_position_23__I_0_add_619_9_lut (.I0(GND_net), .I1(n910), 
            .I2(VCC_net), .I3(n25896), .O(n963)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_9 (.CI(n25896), .I0(n910), 
            .I1(VCC_net), .CO(n25897));
    SB_LUT4 encoder0_position_23__I_0_add_619_8_lut (.I0(GND_net), .I1(n911), 
            .I2(VCC_net), .I3(n25895), .O(n964)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28260_4_lut (.I0(n9_adj_4878), .I1(n7_adj_4876), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n34434));
    defparam i28260_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i28450_4_lut (.I0(n15_adj_4883), .I1(n13_adj_4882), .I2(n11_adj_4880), 
            .I3(n34434), .O(n34624));
    defparam i28450_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_23__I_0_add_619_8 (.CI(n25895), .I0(n911), 
            .I1(VCC_net), .CO(n25896));
    SB_LUT4 i28448_4_lut (.I0(n21_adj_4886), .I1(n19_adj_4885), .I2(n17_adj_4884), 
            .I3(n34624), .O(n34622));
    defparam i28448_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i27964_4_lut (.I0(n27_adj_4889), .I1(n25_adj_4888), .I2(n23_adj_4887), 
            .I3(n34622), .O(n34136));
    defparam i27964_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_619_7_lut (.I0(GND_net), .I1(n912), 
            .I2(GND_net), .I3(n25894), .O(n965)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_687_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4874));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_CARRY encoder0_position_23__I_0_add_619_7 (.CI(n25894), .I0(n912), 
            .I1(GND_net), .CO(n25895));
    SB_LUT4 encoder0_position_23__I_0_add_619_6_lut (.I0(GND_net), .I1(n913), 
            .I2(GND_net), .I3(n25893), .O(n966)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_6 (.CI(n25893), .I0(n913), 
            .I1(GND_net), .CO(n25894));
    SB_LUT4 encoder0_position_23__I_0_add_619_5_lut (.I0(GND_net), .I1(n914), 
            .I2(VCC_net), .I3(n25892), .O(n967)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28598_3_lut (.I0(n4_adj_4874), .I1(pwm_setpoint[13]), .I2(n27_adj_4889), 
            .I3(GND_net), .O(n34772));   // verilog/pwm.v(21[8:24])
    defparam i28598_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_5 (.CI(n25892), .I0(n914), 
            .I1(VCC_net), .CO(n25893));
    SB_LUT4 encoder0_position_23__I_0_add_619_4_lut (.I0(GND_net), .I1(n915), 
            .I2(GND_net), .I3(n25891), .O(n968)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_687_i30_3_lut (.I0(n12_adj_4881), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4891));   // verilog/pwm.v(21[8:24])
    defparam LessThan_687_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_4 (.CI(n25891), .I0(n915), 
            .I1(GND_net), .CO(n25892));
    SB_LUT4 encoder0_position_23__I_0_add_619_3_lut (.I0(GND_net), .I1(n916), 
            .I2(VCC_net), .I3(n25890), .O(n969)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_3 (.CI(n25890), .I0(n916), 
            .I1(VCC_net), .CO(n25891));
    SB_LUT4 i13746_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13933), .I3(GND_net), .O(n18326));   // verilog/coms.v(127[12] 300[6])
    defparam i13746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_2_lut (.I0(GND_net), .I1(n518), 
            .I2(GND_net), .I3(VCC_net), .O(n970)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_2 (.CI(VCC_net), .I0(n518), 
            .I1(GND_net), .CO(n25890));
    SB_LUT4 encoder0_position_23__I_0_add_566_10_lut (.I0(GND_net), .I1(n830), 
            .I2(VCC_net), .I3(n25889), .O(n883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_9_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n25888), .O(n884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_9 (.CI(n25888), .I0(n831), 
            .I1(VCC_net), .CO(n25889));
    SB_LUT4 encoder0_position_23__I_0_add_566_8_lut (.I0(GND_net), .I1(n832), 
            .I2(VCC_net), .I3(n25887), .O(n885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_8 (.CI(n25887), .I0(n832), 
            .I1(VCC_net), .CO(n25888));
    SB_LUT4 encoder0_position_23__I_0_add_566_7_lut (.I0(GND_net), .I1(n833), 
            .I2(GND_net), .I3(n25886), .O(n886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_7 (.CI(n25886), .I0(n833), 
            .I1(GND_net), .CO(n25887));
    SB_LUT4 i28599_3_lut (.I0(n34772), .I1(pwm_setpoint[14]), .I2(n29_adj_4890), 
            .I3(GND_net), .O(n34773));   // verilog/pwm.v(21[8:24])
    defparam i28599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_566_6_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(n25885), .O(n887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_6 (.CI(n25885), .I0(n834), 
            .I1(GND_net), .CO(n25886));
    SB_LUT4 encoder0_position_23__I_0_add_566_5_lut (.I0(GND_net), .I1(n835), 
            .I2(VCC_net), .I3(n25884), .O(n888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_5 (.CI(n25884), .I0(n835), 
            .I1(VCC_net), .CO(n25885));
    SB_LUT4 encoder0_position_23__I_0_add_566_4_lut (.I0(GND_net), .I1(n836), 
            .I2(GND_net), .I3(n25883), .O(n889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_4 (.CI(n25883), .I0(n836), 
            .I1(GND_net), .CO(n25884));
    SB_LUT4 i27958_4_lut (.I0(n33), .I1(n31_adj_4892), .I2(n29_adj_4890), 
            .I3(n34134), .O(n34130));
    defparam i27958_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_566_3_lut (.I0(GND_net), .I1(n837), 
            .I2(VCC_net), .I3(n25882), .O(n890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_3 (.CI(n25882), .I0(n837), 
            .I1(VCC_net), .CO(n25883));
    SB_LUT4 encoder0_position_23__I_0_add_566_2_lut (.I0(GND_net), .I1(n517), 
            .I2(GND_net), .I3(VCC_net), .O(n891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_2 (.CI(VCC_net), .I0(n517), 
            .I1(GND_net), .CO(n25882));
    SB_LUT4 i13747_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13933), .I3(GND_net), .O(n18327));   // verilog/coms.v(127[12] 300[6])
    defparam i13747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13748_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13933), .I3(GND_net), .O(n18328));   // verilog/coms.v(127[12] 300[6])
    defparam i13748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28697_4_lut (.I0(n30_adj_4891), .I1(n10_adj_4879), .I2(n35), 
            .I3(n34127), .O(n34871));   // verilog/pwm.v(21[8:24])
    defparam i28697_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13749_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13933), .I3(GND_net), .O(n18329));   // verilog/coms.v(127[12] 300[6])
    defparam i13749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13750_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13933), .I3(GND_net), .O(n18330));   // verilog/coms.v(127[12] 300[6])
    defparam i13750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13751_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13933), .I3(GND_net), .O(n18331));   // verilog/coms.v(127[12] 300[6])
    defparam i13751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13752_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13933), .I3(GND_net), .O(n18332));   // verilog/coms.v(127[12] 300[6])
    defparam i13752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13753_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13933), .I3(GND_net), .O(n18333));   // verilog/coms.v(127[12] 300[6])
    defparam i13753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13754_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13933), .I3(GND_net), .O(n18334));   // verilog/coms.v(127[12] 300[6])
    defparam i13754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13755_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13933), .I3(GND_net), .O(n18335));   // verilog/coms.v(127[12] 300[6])
    defparam i13755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28573_3_lut (.I0(n34773), .I1(pwm_setpoint[15]), .I2(n31_adj_4892), 
            .I3(GND_net), .O(n34747));   // verilog/pwm.v(21[8:24])
    defparam i28573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13756_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13933), .I3(GND_net), .O(n18336));   // verilog/coms.v(127[12] 300[6])
    defparam i13756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13757_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13933), .I3(GND_net), .O(n18337));   // verilog/coms.v(127[12] 300[6])
    defparam i13757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13758_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13933), .I3(GND_net), .O(n18338));   // verilog/coms.v(127[12] 300[6])
    defparam i13758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3158_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4831), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1733_6_lut (.I0(n33075), .I1(n510), .I2(GND_net), .I3(n25653), 
            .O(n33988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_6_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i13759_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13933), .I3(GND_net), .O(n18339));   // verilog/coms.v(127[12] 300[6])
    defparam i13759_3_lut.LUT_INIT = 16'hcaca;
    GND i1 (.Y(GND_net));
    SB_CARRY add_1733_6 (.CI(n25653), .I0(n510), .I1(GND_net), .CO(n25654));
    SB_LUT4 i13760_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13933), .I3(GND_net), .O(n18340));   // verilog/coms.v(127[12] 300[6])
    defparam i13760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13475_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n32040), .I3(GND_net), .O(n18055));   // verilog/coms.v(127[12] 300[6])
    defparam i13475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1733_5_lut (.I0(GND_net), .I1(n511), .I2(VCC_net), .I3(n25652), 
            .O(n5275)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_26[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_CARRY add_1733_5 (.CI(n25652), .I0(n511), .I1(VCC_net), .CO(n25653));
    SB_LUT4 i26907_1_lut (.I0(n4_adj_4927), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n33075));
    defparam i26907_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3158_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4829), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n510));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3158_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n3_adj_4816), .I3(n25855), .O(displacement_23__N_50[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28600_3_lut (.I0(n6_adj_4875), .I1(pwm_setpoint[10]), .I2(n21_adj_4886), 
            .I3(GND_net), .O(n34774));   // verilog/pwm.v(21[8:24])
    defparam i28600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28601_3_lut (.I0(n34774), .I1(pwm_setpoint[11]), .I2(n23_adj_4887), 
            .I3(GND_net), .O(n34775));   // verilog/pwm.v(21[8:24])
    defparam i28601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4816), .I3(n25854), .O(displacement_23__N_50[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n25854), .I0(encoder1_position[22]), 
            .I1(n3_adj_4816), .CO(n25855));
    SB_LUT4 i28250_4_lut (.I0(n23_adj_4887), .I1(n21_adj_4886), .I2(n19_adj_4885), 
            .I3(n34142), .O(n34424));
    defparam i28250_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n3_adj_4816), .I3(n25853), .O(displacement_23__N_50[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n25853), .I0(encoder1_position[21]), 
            .I1(n3_adj_4816), .CO(n25854));
    SB_CARRY add_615_4 (.CI(n25586), .I0(n35425), .I1(n23_adj_4799), .CO(n25587));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4787), .I3(n25852), .O(displacement_23__N_50[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_4899), .I3(n26460), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1733_4_lut (.I0(GND_net), .I1(n425), .I2(GND_net), .I3(n25651), 
            .O(n5276)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4900), .I3(n26459), .O(n3_adj_4829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_25 (.CI(n26459), 
            .I0(GND_net), .I1(n3_adj_4900), .CO(n26460));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4901), .I3(n26458), .O(n4_adj_4831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1733_4 (.CI(n25651), .I0(n425), .I1(GND_net), .CO(n25652));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_24 (.CI(n26458), 
            .I0(GND_net), .I1(n4_adj_4901), .CO(n26459));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4902), .I3(n26457), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1733_3_lut (.I0(GND_net), .I1(n513), .I2(VCC_net), .I3(n25650), 
            .O(n5277)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_23 (.CI(n26457), 
            .I0(GND_net), .I1(n5_adj_4902), .CO(n26458));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4903), .I3(n26456), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_22 (.CI(n26456), 
            .I0(GND_net), .I1(n6_adj_4903), .CO(n26457));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4904), .I3(n26455), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_21 (.CI(n26455), 
            .I0(GND_net), .I1(n7_adj_4904), .CO(n26456));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_4905), .I3(n26454), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_20 (.CI(n26454), 
            .I0(GND_net), .I1(n8_adj_4905), .CO(n26455));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_4906), .I3(n26453), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_19 (.CI(n26453), 
            .I0(GND_net), .I1(n9_adj_4906), .CO(n26454));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_4907), .I3(n26452), .O(n10_adj_4827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_18 (.CI(n26452), 
            .I0(GND_net), .I1(n10_adj_4907), .CO(n26453));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_4908), .I3(n26451), .O(n11_adj_4785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_17 (.CI(n26451), 
            .I0(GND_net), .I1(n11_adj_4908), .CO(n26452));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_4909), .I3(n26450), .O(n12_adj_4849)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_16 (.CI(n26450), 
            .I0(GND_net), .I1(n12_adj_4909), .CO(n26451));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_4910), .I3(n26449), .O(n13_adj_4848)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n25852), .I0(encoder1_position[20]), 
            .I1(n5_adj_4787), .CO(n25853));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_15 (.CI(n26449), 
            .I0(GND_net), .I1(n13_adj_4910), .CO(n26450));
    SB_CARRY add_1733_3 (.CI(n25650), .I0(n513), .I1(VCC_net), .CO(n25651));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_4911), .I3(n26448), .O(n14_adj_4820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4786), .I3(n25851), .O(displacement_23__N_50[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_14 (.CI(n26448), 
            .I0(GND_net), .I1(n14_adj_4911), .CO(n26449));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_4912), .I3(n26447), .O(n15_adj_4847)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n25851), .I0(encoder1_position[19]), 
            .I1(n6_adj_4786), .CO(n25852));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_13 (.CI(n26447), 
            .I0(GND_net), .I1(n15_adj_4912), .CO(n26448));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_4913), .I3(n26446), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_12 (.CI(n26446), 
            .I0(GND_net), .I1(n16_adj_4913), .CO(n26447));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_4914), .I3(n26445), .O(n17_adj_4841)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_11 (.CI(n26445), 
            .I0(GND_net), .I1(n17_adj_4914), .CO(n26446));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_4915), .I3(n26444), .O(n18_adj_4836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_59_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4835), .I3(n15_adj_4828), .O(motor_state_23__N_74[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_59_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_10 (.CI(n26444), 
            .I0(GND_net), .I1(n18_adj_4915), .CO(n26445));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_4916), .I3(n26443), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_9 (.CI(n26443), 
            .I0(GND_net), .I1(n19_adj_4916), .CO(n26444));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_4917), .I3(n26442), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_8 (.CI(n26442), 
            .I0(GND_net), .I1(n20_adj_4917), .CO(n26443));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_4918), .I3(n26441), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_7 (.CI(n26441), 
            .I0(GND_net), .I1(n21_adj_4918), .CO(n26442));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_4919), .I3(n26440), .O(n22_adj_4843)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_6 (.CI(n26440), 
            .I0(GND_net), .I1(n22_adj_4919), .CO(n26441));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_4920), .I3(n26439), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_5 (.CI(n26439), 
            .I0(GND_net), .I1(n23_adj_4920), .CO(n26440));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_4921), .I3(n26438), .O(n24_adj_4839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_4 (.CI(n26438), 
            .I0(GND_net), .I1(n24_adj_4921), .CO(n26439));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_4922), .I3(n26437), .O(n25_adj_4842)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_3 (.CI(n26437), 
            .I0(GND_net), .I1(n25_adj_4922), .CO(n26438));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n26437));
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4851), .I3(n25850), .O(displacement_23__N_50[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n25850), .I0(encoder1_position[18]), 
            .I1(n7_adj_4851), .CO(n25851));
    SB_LUT4 add_1733_2_lut (.I0(GND_net), .I1(n514), .I2(GND_net), .I3(VCC_net), 
            .O(n5278)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1733_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4852), .I3(n25849), .O(displacement_23__N_50[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n25849), .I0(encoder1_position[17]), 
            .I1(n8_adj_4852), .CO(n25850));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4853), .I3(n25848), .O(displacement_23__N_50[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n25848), .I0(encoder1_position[16]), 
            .I1(n9_adj_4853), .CO(n25849));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4854), .I3(n25847), .O(displacement_23__N_50[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n25847), .I0(encoder1_position[15]), 
            .I1(n10_adj_4854), .CO(n25848));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4855), .I3(n25846), .O(displacement_23__N_50[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n25846), .I0(encoder1_position[14]), 
            .I1(n11_adj_4855), .CO(n25847));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4856), .I3(n25845), .O(displacement_23__N_50[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n25845), .I0(encoder1_position[13]), 
            .I1(n12_adj_4856), .CO(n25846));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4857), .I3(n25844), .O(displacement_23__N_50[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n25844), .I0(encoder1_position[12]), 
            .I1(n13_adj_4857), .CO(n25845));
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4858), .I3(n25843), .O(displacement_23__N_50[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n25843), .I0(encoder1_position[11]), 
            .I1(n14_adj_4858), .CO(n25844));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4859), .I3(n25842), .O(displacement_23__N_50[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n25842), .I0(encoder1_position[10]), 
            .I1(n15_adj_4859), .CO(n25843));
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4860), .I3(n25841), .O(displacement_23__N_50[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n25841), .I0(encoder1_position[9]), 
            .I1(n16_adj_4860), .CO(n25842));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4861), .I3(n25840), .O(displacement_23__N_50[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n25840), .I0(encoder1_position[8]), 
            .I1(n17_adj_4861), .CO(n25841));
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4862), .I3(n25839), .O(displacement_23__N_50[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n25839), .I0(encoder1_position[7]), 
            .I1(n18_adj_4862), .CO(n25840));
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4863), .I3(n25838), .O(displacement_23__N_50[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n25838), .I0(encoder1_position[6]), 
            .I1(n19_adj_4863), .CO(n25839));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4864), .I3(n25837), .O(displacement_23__N_50[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n25837), .I0(encoder1_position[5]), 
            .I1(n20_adj_4864), .CO(n25838));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4865), .I3(n25836), .O(displacement_23__N_50[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13761_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13933), .I3(GND_net), .O(n18341));   // verilog/coms.v(127[12] 300[6])
    defparam i13761_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n25836), .I0(encoder1_position[4]), 
            .I1(n21_adj_4865), .CO(n25837));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4866), .I3(n25835), .O(displacement_23__N_50[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n25835), .I0(encoder1_position[3]), 
            .I1(n22_adj_4866), .CO(n25836));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4867), .I3(n25834), .O(displacement_23__N_50[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n25834), .I0(encoder1_position[2]), 
            .I1(n23_adj_4867), .CO(n25835));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4868), .I3(n25833), .O(displacement_23__N_50[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n25833), .I0(encoder1_position[1]), 
            .I1(n24_adj_4868), .CO(n25834));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4869), .I3(VCC_net), .O(displacement_23__N_50[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4869), .CO(n25833));
    SB_LUT4 i13762_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13933), .I3(GND_net), .O(n18342));   // verilog/coms.v(127[12] 300[6])
    defparam i13762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13763_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13933), .I3(GND_net), .O(n18343));   // verilog/coms.v(127[12] 300[6])
    defparam i13763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13764_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13933), .I3(GND_net), .O(n18344));   // verilog/coms.v(127[12] 300[6])
    defparam i13764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13765_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13933), .I3(GND_net), .O(n18345));   // verilog/coms.v(127[12] 300[6])
    defparam i13765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13766_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13933), 
            .I3(GND_net), .O(n18346));   // verilog/coms.v(127[12] 300[6])
    defparam i13766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28492_3_lut (.I0(n8_adj_4877), .I1(pwm_setpoint[9]), .I2(n19_adj_4885), 
            .I3(GND_net), .O(n34666));   // verilog/pwm.v(21[8:24])
    defparam i28492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28571_3_lut (.I0(n34775), .I1(pwm_setpoint[12]), .I2(n25_adj_4888), 
            .I3(GND_net), .O(n34745));   // verilog/pwm.v(21[8:24])
    defparam i28571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13767_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13933), 
            .I3(GND_net), .O(n18347));   // verilog/coms.v(127[12] 300[6])
    defparam i13767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25067_2_lut (.I0(n16606), .I1(n3303), .I2(GND_net), .I3(GND_net), 
            .O(n31225));
    defparam i25067_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1693 (.I0(n30480), .I1(n16613), .I2(n31225), 
            .I3(n771), .O(n33043));
    defparam i3_4_lut_adj_1693.LUT_INIT = 16'hafbf;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n63), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n33043), .I3(n13810), .O(n29947));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'hd5f5;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4788));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_4_lut (.I0(n16613), .I1(n63_adj_4873), .I2(n771), 
            .I3(n19_adj_4893), .O(n5_adj_4932));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcc04;
    SB_LUT4 i13477_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n32962), 
            .I3(GND_net), .O(n18057));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13477_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13768_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13933), 
            .I3(GND_net), .O(n18348));   // verilog/coms.v(127[12] 300[6])
    defparam i13768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13769_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13933), 
            .I3(GND_net), .O(n18349));   // verilog/coms.v(127[12] 300[6])
    defparam i13769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13770_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13933), 
            .I3(GND_net), .O(n18350));   // verilog/coms.v(127[12] 300[6])
    defparam i13770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13771_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13933), 
            .I3(GND_net), .O(n18351));   // verilog/coms.v(127[12] 300[6])
    defparam i13771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13772_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13933), 
            .I3(GND_net), .O(n18352));   // verilog/coms.v(127[12] 300[6])
    defparam i13772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13773_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13933), 
            .I3(GND_net), .O(n18353));   // verilog/coms.v(127[12] 300[6])
    defparam i13773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13774_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13933), 
            .I3(GND_net), .O(n18354));   // verilog/coms.v(127[12] 300[6])
    defparam i13774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13775_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13933), 
            .I3(GND_net), .O(n18355));   // verilog/coms.v(127[12] 300[6])
    defparam i13775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13776_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13933), 
            .I3(GND_net), .O(n18356));   // verilog/coms.v(127[12] 300[6])
    defparam i13776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13777_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13933), 
            .I3(GND_net), .O(n18357));   // verilog/coms.v(127[12] 300[6])
    defparam i13777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13778_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13933), 
            .I3(GND_net), .O(n18358));   // verilog/coms.v(127[12] 300[6])
    defparam i13778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13779_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13933), 
            .I3(GND_net), .O(n18359));   // verilog/coms.v(127[12] 300[6])
    defparam i13779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13780_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13933), 
            .I3(GND_net), .O(n18360));   // verilog/coms.v(127[12] 300[6])
    defparam i13780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13781_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13933), 
            .I3(GND_net), .O(n18361));   // verilog/coms.v(127[12] 300[6])
    defparam i13781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13782_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13933), 
            .I3(GND_net), .O(n18362));   // verilog/coms.v(127[12] 300[6])
    defparam i13782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13783_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13933), 
            .I3(GND_net), .O(n18363));   // verilog/coms.v(127[12] 300[6])
    defparam i13783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13784_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13933), 
            .I3(GND_net), .O(n18364));   // verilog/coms.v(127[12] 300[6])
    defparam i13784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13785_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13933), 
            .I3(GND_net), .O(n18365));   // verilog/coms.v(127[12] 300[6])
    defparam i13785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13786_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13933), 
            .I3(GND_net), .O(n18366));   // verilog/coms.v(127[12] 300[6])
    defparam i13786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13787_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13933), 
            .I3(GND_net), .O(n18367));   // verilog/coms.v(127[12] 300[6])
    defparam i13787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13788_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13933), 
            .I3(GND_net), .O(n18368));   // verilog/coms.v(127[12] 300[6])
    defparam i13788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13789_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13933), 
            .I3(GND_net), .O(n18369));   // verilog/coms.v(127[12] 300[6])
    defparam i13789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13790_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13933), .I3(GND_net), .O(n18370));   // verilog/coms.v(127[12] 300[6])
    defparam i13790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13791_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13933), .I3(GND_net), .O(n18371));   // verilog/coms.v(127[12] 300[6])
    defparam i13791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13792_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13933), .I3(GND_net), .O(n18372));   // verilog/coms.v(127[12] 300[6])
    defparam i13792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13793_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13933), .I3(GND_net), .O(n18373));   // verilog/coms.v(127[12] 300[6])
    defparam i13793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13794_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13933), .I3(GND_net), .O(n18374));   // verilog/coms.v(127[12] 300[6])
    defparam i13794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13795_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13933), .I3(GND_net), .O(n18375));   // verilog/coms.v(127[12] 300[6])
    defparam i13795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13796_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13933), .I3(GND_net), .O(n18376));   // verilog/coms.v(127[12] 300[6])
    defparam i13796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13797_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13933), .I3(GND_net), .O(n18377));   // verilog/coms.v(127[12] 300[6])
    defparam i13797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13798_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13933), .I3(GND_net), .O(n18378));   // verilog/coms.v(127[12] 300[6])
    defparam i13798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13799_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13933), .I3(GND_net), .O(n18379));   // verilog/coms.v(127[12] 300[6])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13800_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13933), .I3(GND_net), .O(n18380));   // verilog/coms.v(127[12] 300[6])
    defparam i13800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13801_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13933), .I3(GND_net), .O(n18381));   // verilog/coms.v(127[12] 300[6])
    defparam i13801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13802_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13933), .I3(GND_net), .O(n18382));   // verilog/coms.v(127[12] 300[6])
    defparam i13802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13803_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13933), .I3(GND_net), .O(n18383));   // verilog/coms.v(127[12] 300[6])
    defparam i13803_3_lut.LUT_INIT = 16'hcaca;
    motorControl control (.\Kp[2] (Kp[2]), .GND_net(GND_net), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .IntegralLimit({IntegralLimit}), .\Kp[5] (Kp[5]), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .PWMLimit({PWMLimit}), 
            .\Ki[0] (Ki[0]), .\Ki[14] (Ki[14]), .duty({duty}), .clk32MHz(clk32MHz), 
            .\Kp[15] (Kp[15]), .VCC_net(VCC_net), .\Ki[15] (Ki[15]), .\Ki[1] (Ki[1]), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Ki[6] (Ki[6]), .\Ki[12] (Ki[12]), .setpoint({setpoint}), 
            .motor_state({motor_state}), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .n35425(n35425), .\Ki[11] (Ki[11]), 
            .\Ki[13] (Ki[13])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_LUT4 i13804_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13933), .I3(GND_net), .O(n18384));   // verilog/coms.v(127[12] 300[6])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13805_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13933), .I3(GND_net), .O(n18385));   // verilog/coms.v(127[12] 300[6])
    defparam i13805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13806_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13933), .I3(GND_net), .O(n18386));   // verilog/coms.v(127[12] 300[6])
    defparam i13806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13807_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13933), .I3(GND_net), .O(n18387));   // verilog/coms.v(127[12] 300[6])
    defparam i13807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13808_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13933), .I3(GND_net), .O(n18388));   // verilog/coms.v(127[12] 300[6])
    defparam i13808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13809_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13933), .I3(GND_net), .O(n18389));   // verilog/coms.v(127[12] 300[6])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13810_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13933), .I3(GND_net), .O(n18390));   // verilog/coms.v(127[12] 300[6])
    defparam i13810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13811_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13933), .I3(GND_net), .O(n18391));   // verilog/coms.v(127[12] 300[6])
    defparam i13811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13812_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13933), .I3(GND_net), .O(n18392));   // verilog/coms.v(127[12] 300[6])
    defparam i13812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13813_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13933), .I3(GND_net), .O(n18393));   // verilog/coms.v(127[12] 300[6])
    defparam i13813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13814_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13933), .I3(GND_net), .O(n18394));   // verilog/coms.v(127[12] 300[6])
    defparam i13814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13815_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13933), .I3(GND_net), .O(n18395));   // verilog/coms.v(127[12] 300[6])
    defparam i13815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13816_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13933), .I3(GND_net), .O(n18396));   // verilog/coms.v(127[12] 300[6])
    defparam i13816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13817_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13933), .I3(GND_net), .O(n18397));   // verilog/coms.v(127[12] 300[6])
    defparam i13817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13818_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13933), .I3(GND_net), .O(n18398));   // verilog/coms.v(127[12] 300[6])
    defparam i13818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13819_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13933), .I3(GND_net), .O(n18399));   // verilog/coms.v(127[12] 300[6])
    defparam i13819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13820_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13933), .I3(GND_net), .O(n18400));   // verilog/coms.v(127[12] 300[6])
    defparam i13820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28536_4_lut (.I0(n33), .I1(n31_adj_4892), .I2(n29_adj_4890), 
            .I3(n34136), .O(n34710));
    defparam i28536_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13821_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13933), .I3(GND_net), .O(n18401));   // verilog/coms.v(127[12] 300[6])
    defparam i13821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13822_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13933), .I3(GND_net), .O(n18402));   // verilog/coms.v(127[12] 300[6])
    defparam i13822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13823_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13933), .I3(GND_net), .O(n18403));   // verilog/coms.v(127[12] 300[6])
    defparam i13823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13824_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13933), .I3(GND_net), .O(n18404));   // verilog/coms.v(127[12] 300[6])
    defparam i13824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28744_4_lut (.I0(n34747), .I1(n34871), .I2(n35), .I3(n34130), 
            .O(n34918));   // verilog/pwm.v(21[8:24])
    defparam i28744_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13825_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13933), .I3(GND_net), .O(n18405));   // verilog/coms.v(127[12] 300[6])
    defparam i13825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13826_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13933), .I3(GND_net), .O(n18406));   // verilog/coms.v(127[12] 300[6])
    defparam i13826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13827_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13933), .I3(GND_net), .O(n18407));   // verilog/coms.v(127[12] 300[6])
    defparam i13827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13828_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13933), .I3(GND_net), .O(n18408));   // verilog/coms.v(127[12] 300[6])
    defparam i13828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13829_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13933), .I3(GND_net), .O(n18409));   // verilog/coms.v(127[12] 300[6])
    defparam i13829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13830_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13933), .I3(GND_net), .O(n18410));   // verilog/coms.v(127[12] 300[6])
    defparam i13830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13831_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13933), .I3(GND_net), .O(n18411));   // verilog/coms.v(127[12] 300[6])
    defparam i13831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13832_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13933), .I3(GND_net), .O(n18412));   // verilog/coms.v(127[12] 300[6])
    defparam i13832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13833_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13933), .I3(GND_net), .O(n18413));   // verilog/coms.v(127[12] 300[6])
    defparam i13833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13834_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13933), .I3(GND_net), .O(n18414));   // verilog/coms.v(127[12] 300[6])
    defparam i13834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13835_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13933), .I3(GND_net), .O(n18415));   // verilog/coms.v(127[12] 300[6])
    defparam i13835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13836_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13933), .I3(GND_net), .O(n18416));   // verilog/coms.v(127[12] 300[6])
    defparam i13836_3_lut.LUT_INIT = 16'hcaca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4833, 
            quadB_debounced_adj_4834}), .ENCODER1_A_c_1(ENCODER1_A_c_1), 
            .reg_B({reg_B_adj_5018}), .n33025(n33025), .VCC_net(VCC_net), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n18059(n18059), .n18544(n18544)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    SB_LUT4 i13837_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13933), .I3(GND_net), .O(n18417));   // verilog/coms.v(127[12] 300[6])
    defparam i13837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13838_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n13933), .I3(GND_net), .O(n18418));   // verilog/coms.v(127[12] 300[6])
    defparam i13838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28594_4_lut (.I0(n34745), .I1(n34666), .I2(n25_adj_4888), 
            .I3(n34424), .O(n34768));   // verilog/pwm.v(21[8:24])
    defparam i28594_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13839_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n13933), .I3(GND_net), .O(n18419));   // verilog/coms.v(127[12] 300[6])
    defparam i13839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13840_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n13933), .I3(GND_net), .O(n18420));   // verilog/coms.v(127[12] 300[6])
    defparam i13840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13841_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n13933), .I3(GND_net), .O(n18421));   // verilog/coms.v(127[12] 300[6])
    defparam i13841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13842_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n13933), .I3(GND_net), .O(n18422));   // verilog/coms.v(127[12] 300[6])
    defparam i13842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13843_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n13933), .I3(GND_net), .O(n18423));   // verilog/coms.v(127[12] 300[6])
    defparam i13843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13844_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n13933), .I3(GND_net), .O(n18424));   // verilog/coms.v(127[12] 300[6])
    defparam i13844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13845_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n13933), .I3(GND_net), .O(n18425));   // verilog/coms.v(127[12] 300[6])
    defparam i13845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13846_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n13933), .I3(GND_net), .O(n18426));   // verilog/coms.v(127[12] 300[6])
    defparam i13846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13847_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n13933), .I3(GND_net), .O(n18427));   // verilog/coms.v(127[12] 300[6])
    defparam i13847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13848_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n13933), .I3(GND_net), .O(n18428));   // verilog/coms.v(127[12] 300[6])
    defparam i13848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13849_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n13933), .I3(GND_net), .O(n18429));   // verilog/coms.v(127[12] 300[6])
    defparam i13849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13850_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n13933), .I3(GND_net), .O(n18430));   // verilog/coms.v(127[12] 300[6])
    defparam i13850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13851_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n13933), .I3(GND_net), .O(n18431));   // verilog/coms.v(127[12] 300[6])
    defparam i13851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13852_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n13933), .I3(GND_net), .O(n18432));   // verilog/coms.v(127[12] 300[6])
    defparam i13852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13853_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n13933), .I3(GND_net), .O(n18433));   // verilog/coms.v(127[12] 300[6])
    defparam i13853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13854_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[22]), 
            .I2(n13933), .I3(GND_net), .O(n18434));   // verilog/coms.v(127[12] 300[6])
    defparam i13854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13855_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n13933), .I3(GND_net), .O(n18435));   // verilog/coms.v(127[12] 300[6])
    defparam i13855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13856_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[22]), 
            .I2(n13933), .I3(GND_net), .O(n18436));   // verilog/coms.v(127[12] 300[6])
    defparam i13856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13478_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5007[1]), .I2(n9799), 
            .I3(n4_adj_4823), .O(n18058));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13478_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i28748_4_lut (.I0(n34768), .I1(n34918), .I2(n35), .I3(n34710), 
            .O(n34922));   // verilog/pwm.v(21[8:24])
    defparam i28748_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28749_3_lut (.I0(n34922), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n34923));   // verilog/pwm.v(21[8:24])
    defparam i28749_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28747_3_lut (.I0(n34923), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n34921));   // verilog/pwm.v(21[8:24])
    defparam i28747_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13857_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n13933), .I3(GND_net), .O(n18437));   // verilog/coms.v(127[12] 300[6])
    defparam i13857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28677_3_lut (.I0(n34921), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n34851));   // verilog/pwm.v(21[8:24])
    defparam i28677_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13858_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n13933), .I3(GND_net), .O(n18438));   // verilog/coms.v(127[12] 300[6])
    defparam i13858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13859_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n13933), .I3(GND_net), .O(n18439));   // verilog/coms.v(127[12] 300[6])
    defparam i13859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13860_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n13933), .I3(GND_net), .O(n18440));   // verilog/coms.v(127[12] 300[6])
    defparam i13860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28678_3_lut (.I0(n34851), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n34852));   // verilog/pwm.v(21[8:24])
    defparam i28678_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13861_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n13933), .I3(GND_net), .O(n18441));   // verilog/coms.v(127[12] 300[6])
    defparam i13861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13862_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13933), .I3(GND_net), .O(n18442));   // verilog/coms.v(127[12] 300[6])
    defparam i13862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13863_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13933), .I3(GND_net), .O(n18443));   // verilog/coms.v(127[12] 300[6])
    defparam i13863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13864_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13933), .I3(GND_net), .O(n18444));   // verilog/coms.v(127[12] 300[6])
    defparam i13864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13865_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13933), .I3(GND_net), .O(n18445));   // verilog/coms.v(127[12] 300[6])
    defparam i13865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13866_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13933), .I3(GND_net), .O(n18446));   // verilog/coms.v(127[12] 300[6])
    defparam i13866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13867_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13933), .I3(GND_net), .O(n18447));   // verilog/coms.v(127[12] 300[6])
    defparam i13867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28579_3_lut (.I0(n34852), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n34753));   // verilog/pwm.v(21[8:24])
    defparam i28579_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13870_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n32040), 
            .I3(GND_net), .O(n18450));   // verilog/coms.v(127[12] 300[6])
    defparam i13870_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.\state[2] (state_adj_5030[2]), .\state[0] (state_adj_5030[0]), 
           .\state[3] (state_adj_5030[3]), .GND_net(GND_net), .n21828(n21828), 
           .n21898(n21898), .n4604(n4604), .n21826(n21826), .CLK_c(CLK_c), 
           .scl_enable(scl_enable), .\state_7__N_3815[0] (state_7__N_3815[0]), 
           .sda_enable(sda_enable), .VCC_net(VCC_net), .n5019(n5019), 
           .n34058(n34058), .\state_7__N_3831[3] (state_7__N_3831[3]), .n10(n10_adj_4832), 
           .n5(n5_adj_4808), .n882({scl}), .n8(n8_adj_4807), .n11(n11)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(244[10] 254[6])
    SB_LUT4 i13871_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n32040), 
            .I3(GND_net), .O(n18451));   // verilog/coms.v(127[12] 300[6])
    defparam i13871_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13872_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n32040), 
            .I3(GND_net), .O(n18452));   // verilog/coms.v(127[12] 300[6])
    defparam i13872_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13873_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n32040), 
            .I3(GND_net), .O(n18453));   // verilog/coms.v(127[12] 300[6])
    defparam i13873_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13874_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n32040), 
            .I3(GND_net), .O(n18454));   // verilog/coms.v(127[12] 300[6])
    defparam i13874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13875_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n32040), 
            .I3(GND_net), .O(n18455));   // verilog/coms.v(127[12] 300[6])
    defparam i13875_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13876_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n32040), 
            .I3(GND_net), .O(n18456));   // verilog/coms.v(127[12] 300[6])
    defparam i13876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13877_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n32040), 
            .I3(GND_net), .O(n18457));   // verilog/coms.v(127[12] 300[6])
    defparam i13877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13878_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n32040), 
            .I3(GND_net), .O(n18458));   // verilog/coms.v(127[12] 300[6])
    defparam i13878_3_lut.LUT_INIT = 16'hacac;
    pwm PWM (.n34753(n34753), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n16458(n16458), .GND_net(GND_net), .pwm_counter({pwm_counter}), 
        .n16456(n16456)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    SB_LUT4 i13879_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n32040), 
            .I3(GND_net), .O(n18459));   // verilog/coms.v(127[12] 300[6])
    defparam i13879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13880_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n32040), 
            .I3(GND_net), .O(n18460));   // verilog/coms.v(127[12] 300[6])
    defparam i13880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13881_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n32040), 
            .I3(GND_net), .O(n18461));   // verilog/coms.v(127[12] 300[6])
    defparam i13881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13882_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n32040), 
            .I3(GND_net), .O(n18462));   // verilog/coms.v(127[12] 300[6])
    defparam i13882_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13883_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n32040), 
            .I3(GND_net), .O(n18463));   // verilog/coms.v(127[12] 300[6])
    defparam i13883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13884_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n32040), 
            .I3(GND_net), .O(n18464));   // verilog/coms.v(127[12] 300[6])
    defparam i13884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13885_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n32040), 
            .I3(GND_net), .O(n18465));   // verilog/coms.v(127[12] 300[6])
    defparam i13885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13886_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n32040), 
            .I3(GND_net), .O(n18466));   // verilog/coms.v(127[12] 300[6])
    defparam i13886_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.clk32MHz(clk32MHz), .GND_net(GND_net), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n30471(n30471), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[5] ({Open_0, Open_1, \data_out_frame[5] [5:2], 
         Open_2, Open_3}), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[5][7] (\data_out_frame[5] [7]), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .\data_out_frame[5][6] (\data_out_frame[5] [6]), 
         .n30475(n30475), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n22632(n22632), .\data_in_frame[1] ({Open_4, Open_5, \data_in_frame[1] [5:4], 
         Open_6, Open_7, Open_8, Open_9}), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[1][6] (\data_in_frame[1] [6]), .\data_in_frame[1][7] (\data_in_frame[1] [7]), 
         .n16613(n16613), .n4922(n4922), .n122(n122), .n16606(n16606), 
         .n3303(n3303), .n63(n63_adj_4873), .n5(n5_adj_4898), .n36350(n36350), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .n63_adj_3(n63), .n2696(n2696), 
         .n4452(n4452), .n16621(n16621), .n13810(n13810), .n771(n771), 
         .n9711(n9711), .n123(n123), .\FRAME_MATCHER.state_31__N_2579[1] (\FRAME_MATCHER.state_31__N_2579 [1]), 
         .\data_in[0] ({\data_in[0] }), .\data_in[1] ({\data_in[1] }), .\data_in[2] ({\data_in[2] }), 
         .\data_in[3] ({\data_in[3] }), .rx_data({rx_data}), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .control_mode({Open_10, Open_11, Open_12, Open_13, control_mode[3:2], 
         Open_14, Open_15}), .n32040(n32040), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .rx_data_ready(rx_data_ready), .setpoint({setpoint}), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n18102(n18102), .n18101(n18101), .n18100(n18100), .n16614(n16614), 
         .n18099(n18099), .n18098(n18098), .\control_mode[6] (control_mode[6]), 
         .\control_mode[7] (control_mode[7]), .\control_mode[4] (control_mode[4]), 
         .\control_mode[5] (control_mode[5]), .n15(n15_adj_4828), .\state[2] (state_adj_5030[2]), 
         .\state[3] (state_adj_5030[3]), .n10(n10_adj_4832), .n15_adj_4(n15_adj_4835), 
         .tx_active(tx_active), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n18097(n18097), .n18096(n18096), .n18095(n18095), .DE_c(DE_c), 
         .n18091(n18091), .n18090(n18090), .n18089(n18089), .n18088(n18088), 
         .n18087(n18087), .PWMLimit({PWMLimit}), .n18086(n18086), .n18085(n18085), 
         .n18084(n18084), .n18083(n18083), .n18082(n18082), .n18081(n18081), 
         .n18080(n18080), .n18079(n18079), .n18078(n18078), .n18077(n18077), 
         .n18076(n18076), .n18075(n18075), .n18074(n18074), .n18073(n18073), 
         .n18072(n18072), .n18071(n18071), .n18070(n18070), .n18069(n18069), 
         .n18068(n18068), .n18067(n18067), .n18066(n18066), .n18065(n18065), 
         .n35879(n35879), .n35882(n35882), .LED_c(LED_c), .n32812(n32812), 
         .\state[0] (state_adj_5030[0]), .n5019(n5019), .n18536(n18536), 
         .IntegralLimit({IntegralLimit}), .n18535(n18535), .n18534(n18534), 
         .n18533(n18533), .n18532(n18532), .n18531(n18531), .n18530(n18530), 
         .n18529(n18529), .n18528(n18528), .n18527(n18527), .n18526(n18526), 
         .n18525(n18525), .n18524(n18524), .n18523(n18523), .n18522(n18522), 
         .n18521(n18521), .n18520(n18520), .n18519(n18519), .n18518(n18518), 
         .n18517(n18517), .n18516(n18516), .n18515(n18515), .n18514(n18514), 
         .n18513(n18513), .n18512(n18512), .n18511(n18511), .n18510(n18510), 
         .n18509(n18509), .n18508(n18508), .n18507(n18507), .n18506(n18506), 
         .n18505(n18505), .n18504(n18504), .n18503(n18503), .n18502(n18502), 
         .n18501(n18501), .n18500(n18500), .n18499(n18499), .n18498(n18498), 
         .n18497(n18497), .n18496(n18496), .n18495(n18495), .n18494(n18494), 
         .n18493(n18493), .n18492(n18492), .n18491(n18491), .n18490(n18490), 
         .n18489(n18489), .n18485(n18485), .n18484(n18484), .n18483(n18483), 
         .n18482(n18482), .n18481(n18481), .n18480(n18480), .n18479(n18479), 
         .\Kp[1] (Kp[1]), .n18478(n18478), .\Kp[2] (Kp[2]), .n18477(n18477), 
         .\Kp[3] (Kp[3]), .n18476(n18476), .\Kp[4] (Kp[4]), .n18475(n18475), 
         .\Kp[5] (Kp[5]), .n18474(n18474), .\Kp[6] (Kp[6]), .n18473(n18473), 
         .\Kp[7] (Kp[7]), .n18472(n18472), .\Kp[8] (Kp[8]), .n18471(n18471), 
         .\Kp[9] (Kp[9]), .n18470(n18470), .\Kp[10] (Kp[10]), .n18469(n18469), 
         .\Kp[11] (Kp[11]), .n18468(n18468), .\Kp[12] (Kp[12]), .n18467(n18467), 
         .\Kp[13] (Kp[13]), .n18466(n18466), .\Kp[14] (Kp[14]), .n18465(n18465), 
         .\Kp[15] (Kp[15]), .n18464(n18464), .\Ki[1] (Ki[1]), .n18463(n18463), 
         .\Ki[2] (Ki[2]), .n18462(n18462), .\Ki[3] (Ki[3]), .n18461(n18461), 
         .\Ki[4] (Ki[4]), .n18460(n18460), .\Ki[5] (Ki[5]), .n18459(n18459), 
         .\Ki[6] (Ki[6]), .n18458(n18458), .\Ki[7] (Ki[7]), .n18457(n18457), 
         .\Ki[8] (Ki[8]), .n18456(n18456), .\Ki[9] (Ki[9]), .n18455(n18455), 
         .\Ki[10] (Ki[10]), .n18454(n18454), .\Ki[11] (Ki[11]), .n18453(n18453), 
         .\Ki[12] (Ki[12]), .n18452(n18452), .\Ki[13] (Ki[13]), .n18451(n18451), 
         .\Ki[14] (Ki[14]), .n18450(n18450), .\Ki[15] (Ki[15]), .n18447(n18447), 
         .n18446(n18446), .n18445(n18445), .n18444(n18444), .n18443(n18443), 
         .n18442(n18442), .n18441(n18441), .n18440(n18440), .n18439(n18439), 
         .n18438(n18438), .n18437(n18437), .n18436(n18436), .n18435(n18435), 
         .n18434(n18434), .n18433(n18433), .n18432(n18432), .n18431(n18431), 
         .n18430(n18430), .n18429(n18429), .n18428(n18428), .n18427(n18427), 
         .n18426(n18426), .n18425(n18425), .n18424(n18424), .n18423(n18423), 
         .n18422(n18422), .n18421(n18421), .n18420(n18420), .n18419(n18419), 
         .n18418(n18418), .n18417(n18417), .n18416(n18416), .n18415(n18415), 
         .n18414(n18414), .n18413(n18413), .n18412(n18412), .n18411(n18411), 
         .n18410(n18410), .n18409(n18409), .n18408(n18408), .n18407(n18407), 
         .n18406(n18406), .n18405(n18405), .n18404(n18404), .n18403(n18403), 
         .n18402(n18402), .n18401(n18401), .n18400(n18400), .n18399(n18399), 
         .n18398(n18398), .n18397(n18397), .n18396(n18396), .n18395(n18395), 
         .n18394(n18394), .n18393(n18393), .n18392(n18392), .n18391(n18391), 
         .n18390(n18390), .n18389(n18389), .n18388(n18388), .n18387(n18387), 
         .n18386(n18386), .n18385(n18385), .n18384(n18384), .n18383(n18383), 
         .n18382(n18382), .n18381(n18381), .n18380(n18380), .n18379(n18379), 
         .n18378(n18378), .n18377(n18377), .n18376(n18376), .n18375(n18375), 
         .n18374(n18374), .n18373(n18373), .n18372(n18372), .n18371(n18371), 
         .n18370(n18370), .n18369(n18369), .n18368(n18368), .n18367(n18367), 
         .n18366(n18366), .n18365(n18365), .n18364(n18364), .n18363(n18363), 
         .n18362(n18362), .n18361(n18361), .n18360(n18360), .n18359(n18359), 
         .n18358(n18358), .n18357(n18357), .n18356(n18356), .n18355(n18355), 
         .n18354(n18354), .n18353(n18353), .n18352(n18352), .n18351(n18351), 
         .n18350(n18350), .n18349(n18349), .n18348(n18348), .n29947(n29947), 
         .n18347(n18347), .n18346(n18346), .n18345(n18345), .n18344(n18344), 
         .n18343(n18343), .n18342(n18342), .n18341(n18341), .n18055(n18055), 
         .n18340(n18340), .n18339(n18339), .n18338(n18338), .n18337(n18337), 
         .n18336(n18336), .n18335(n18335), .n18334(n18334), .n18333(n18333), 
         .n18332(n18332), .n18331(n18331), .n18330(n18330), .n18329(n18329), 
         .n18328(n18328), .n18327(n18327), .n18326(n18326), .n18325(n18325), 
         .n18324(n18324), .n18323(n18323), .n18317(n18317), .n18316(n18316), 
         .n18315(n18315), .n18314(n18314), .n18313(n18313), .n18312(n18312), 
         .n18311(n18311), .n18310(n18310), .n18309(n18309), .n18308(n18308), 
         .n18307(n18307), .n18306(n18306), .n18305(n18305), .n18304(n18304), 
         .n18303(n18303), .n18302(n18302), .n18301(n18301), .n18300(n18300), 
         .n18052(n18052), .neopxl_color({neopxl_color}), .n18051(n18051), 
         .\Ki[0] (Ki[0]), .n18050(n18050), .\Kp[0] (Kp[0]), .n18049(n18049), 
         .n18299(n18299), .n18298(n18298), .n18297(n18297), .n18296(n18296), 
         .n18295(n18295), .n18294(n18294), .n18293(n18293), .n18040(n18040), 
         .n18292(n18292), .n18291(n18291), .n18290(n18290), .n18289(n18289), 
         .n18288(n18288), .n18287(n18287), .n18286(n18286), .n18285(n18285), 
         .n18284(n18284), .n18283(n18283), .n18282(n18282), .n18281(n18281), 
         .n18280(n18280), .n18279(n18279), .n18278(n18278), .n18277(n18277), 
         .n18276(n18276), .n18275(n18275), .n18274(n18274), .n18273(n18273), 
         .n18272(n18272), .n18271(n18271), .n18270(n18270), .n18230(n18230), 
         .n18229(n18229), .n18228(n18228), .n18227(n18227), .n18226(n18226), 
         .n18225(n18225), .n18224(n18224), .n18223(n18223), .n18166(n18166), 
         .n18165(n18165), .n18164(n18164), .n18163(n18163), .n18162(n18162), 
         .n18161(n18161), .n18160(n18160), .n18159(n18159), .n19(n19_adj_4893), 
         .\motor_state_23__N_74[0] (motor_state_23__N_74[0]), .\encoder0_position_scaled[0] (encoder0_position_scaled[0]), 
         .motor_state({motor_state}), .\motor_state_23__N_74[1] (motor_state_23__N_74[1]), 
         .\encoder0_position_scaled[1] (encoder0_position_scaled[1]), .\motor_state_23__N_74[2] (motor_state_23__N_74[2]), 
         .\encoder0_position_scaled[2] (encoder0_position_scaled[2]), .\motor_state_23__N_74[3] (motor_state_23__N_74[3]), 
         .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), .\motor_state_23__N_74[4] (motor_state_23__N_74[4]), 
         .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), .\motor_state_23__N_74[5] (motor_state_23__N_74[5]), 
         .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), .\motor_state_23__N_74[6] (motor_state_23__N_74[6]), 
         .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), .\motor_state_23__N_74[7] (motor_state_23__N_74[7]), 
         .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), .\motor_state_23__N_74[8] (motor_state_23__N_74[8]), 
         .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), .\motor_state_23__N_74[9] (motor_state_23__N_74[9]), 
         .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), .\motor_state_23__N_74[10] (motor_state_23__N_74[10]), 
         .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), .\motor_state_23__N_74[11] (motor_state_23__N_74[11]), 
         .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), .\motor_state_23__N_74[12] (motor_state_23__N_74[12]), 
         .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), .\motor_state_23__N_74[13] (motor_state_23__N_74[13]), 
         .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), .\motor_state_23__N_74[14] (motor_state_23__N_74[14]), 
         .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), .\motor_state_23__N_74[15] (motor_state_23__N_74[15]), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .\motor_state_23__N_74[16] (motor_state_23__N_74[16]), 
         .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), .\motor_state_23__N_74[17] (motor_state_23__N_74[17]), 
         .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), .\motor_state_23__N_74[18] (motor_state_23__N_74[18]), 
         .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), .\motor_state_23__N_74[19] (motor_state_23__N_74[19]), 
         .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), .\motor_state_23__N_74[20] (motor_state_23__N_74[20]), 
         .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), .\motor_state_23__N_74[21] (motor_state_23__N_74[21]), 
         .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), .\motor_state_23__N_74[23] (motor_state_23__N_74[23]), 
         .\motor_state_23__N_74[22] (motor_state_23__N_74[22]), .n13933(n13933), 
         .n30466(n30466), .VCC_net(VCC_net), .n17831(n17831), .n17982(n17982), 
         .r_SM_Main({r_SM_Main_adj_5007}), .\r_SM_Main_2__N_3404[1] (r_SM_Main_2__N_3404[1]), 
         .tx_o(tx_o), .\r_Bit_Index[0] (r_Bit_Index_adj_5009[0]), .n4(n4_adj_4823), 
         .n18322(n18322), .n18058(n18058), .n35944(n35944), .n9799(n9799), 
         .tx_enable(tx_enable), .n17825(n17825), .n17980(n17980), .\r_Bit_Index[0]_adj_5 (r_Bit_Index[0]), 
         .n16549(n16549), .n4_adj_6(n4), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
         .n18488(n18488), .n21943(n21943), .n4_adj_7(n4_adj_4846), .n4_adj_8(n4_adj_4840), 
         .n16544(n16544), .n18540(n18540), .n18048(n18048), .n18047(n18047), 
         .n18046(n18046), .n18045(n18045), .n18044(n18044), .n18043(n18043), 
         .n18042(n18042)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    SB_LUT4 i13887_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n32040), 
            .I3(GND_net), .O(n18467));   // verilog/coms.v(127[12] 300[6])
    defparam i13887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13888_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n32040), 
            .I3(GND_net), .O(n18468));   // verilog/coms.v(127[12] 300[6])
    defparam i13888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13889_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n32040), 
            .I3(GND_net), .O(n18469));   // verilog/coms.v(127[12] 300[6])
    defparam i13889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13890_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n32040), 
            .I3(GND_net), .O(n18470));   // verilog/coms.v(127[12] 300[6])
    defparam i13890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13891_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n32040), 
            .I3(GND_net), .O(n18471));   // verilog/coms.v(127[12] 300[6])
    defparam i13891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13892_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n32040), 
            .I3(GND_net), .O(n18472));   // verilog/coms.v(127[12] 300[6])
    defparam i13892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13893_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n32040), 
            .I3(GND_net), .O(n18473));   // verilog/coms.v(127[12] 300[6])
    defparam i13893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13894_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n32040), 
            .I3(GND_net), .O(n18474));   // verilog/coms.v(127[12] 300[6])
    defparam i13894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13895_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n32040), 
            .I3(GND_net), .O(n18475));   // verilog/coms.v(127[12] 300[6])
    defparam i13895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13896_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n32040), 
            .I3(GND_net), .O(n18476));   // verilog/coms.v(127[12] 300[6])
    defparam i13896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13897_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n32040), 
            .I3(GND_net), .O(n18477));   // verilog/coms.v(127[12] 300[6])
    defparam i13897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13898_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n32040), 
            .I3(GND_net), .O(n18478));   // verilog/coms.v(127[12] 300[6])
    defparam i13898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13899_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n32040), 
            .I3(GND_net), .O(n18479));   // verilog/coms.v(127[12] 300[6])
    defparam i13899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13900_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18480));   // verilog/coms.v(127[12] 300[6])
    defparam i13900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13901_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18481));   // verilog/coms.v(127[12] 300[6])
    defparam i13901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13902_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18482));   // verilog/coms.v(127[12] 300[6])
    defparam i13902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13903_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18483));   // verilog/coms.v(127[12] 300[6])
    defparam i13903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13904_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18484));   // verilog/coms.v(127[12] 300[6])
    defparam i13904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13905_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18485));   // verilog/coms.v(127[12] 300[6])
    defparam i13905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13909_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18489));   // verilog/coms.v(127[12] 300[6])
    defparam i13909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13910_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18490));   // verilog/coms.v(127[12] 300[6])
    defparam i13910_3_lut.LUT_INIT = 16'hcaca;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, clk32MHz, 
            data_o, VCC_net, reg_B, n32962, ENCODER0_B_c_0, n18541, 
            n18057, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    input VCC_net;
    output [1:0]reg_B;
    output n32962;
    input ENCODER0_B_c_0;
    input n18541;
    input n18057;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2906;
    
    wire n2902, n25692, n25693, n25691, n25690, count_enable, B_delayed, 
        A_delayed, n25689, n25688, n25687, n25686, n25685, n25684, 
        n25683, n25682, n25681, n25680, n25679, count_direction, 
        n25678, n25701, n25700, n25699, n25698, n25697, n25696, 
        n25695, n25694;
    
    SB_LUT4 add_684_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2902), 
            .I3(n25692), .O(n2906[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_16 (.CI(n25692), .I0(encoder0_position[14]), .I1(n2902), 
            .CO(n25693));
    SB_LUT4 add_684_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2902), 
            .I3(n25691), .O(n2906[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_15 (.CI(n25691), .I0(encoder0_position[13]), .I1(n2902), 
            .CO(n25692));
    SB_LUT4 add_684_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2902), 
            .I3(n25690), .O(n2906[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[0]));   // quad.v(35[10] 41[6])
    SB_CARRY add_684_14 (.CI(n25690), .I0(encoder0_position[12]), .I1(n2902), 
            .CO(n25691));
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_684_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2902), 
            .I3(n25689), .O(n2906[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_13 (.CI(n25689), .I0(encoder0_position[11]), .I1(n2902), 
            .CO(n25690));
    SB_LUT4 add_684_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2902), 
            .I3(n25688), .O(n2906[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_12 (.CI(n25688), .I0(encoder0_position[10]), .I1(n2902), 
            .CO(n25689));
    SB_LUT4 add_684_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2902), 
            .I3(n25687), .O(n2906[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_11 (.CI(n25687), .I0(encoder0_position[9]), .I1(n2902), 
            .CO(n25688));
    SB_LUT4 add_684_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2902), 
            .I3(n25686), .O(n2906[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_10 (.CI(n25686), .I0(encoder0_position[8]), .I1(n2902), 
            .CO(n25687));
    SB_LUT4 add_684_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2902), 
            .I3(n25685), .O(n2906[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_9 (.CI(n25685), .I0(encoder0_position[7]), .I1(n2902), 
            .CO(n25686));
    SB_LUT4 add_684_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2902), 
            .I3(n25684), .O(n2906[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_8 (.CI(n25684), .I0(encoder0_position[6]), .I1(n2902), 
            .CO(n25685));
    SB_LUT4 add_684_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2902), 
            .I3(n25683), .O(n2906[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[3]));   // quad.v(35[10] 41[6])
    SB_CARRY add_684_7 (.CI(n25683), .I0(encoder0_position[5]), .I1(n2902), 
            .CO(n25684));
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2906[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_684_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2902), 
            .I3(n25682), .O(n2906[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_6 (.CI(n25682), .I0(encoder0_position[4]), .I1(n2902), 
            .CO(n25683));
    SB_LUT4 add_684_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2902), 
            .I3(n25681), .O(n2906[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_5 (.CI(n25681), .I0(encoder0_position[3]), .I1(n2902), 
            .CO(n25682));
    SB_LUT4 add_684_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2902), 
            .I3(n25680), .O(n2906[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_4 (.CI(n25680), .I0(encoder0_position[2]), .I1(n2902), 
            .CO(n25681));
    SB_LUT4 add_684_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2902), 
            .I3(n25679), .O(n2906[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_3 (.CI(n25679), .I0(encoder0_position[1]), .I1(n2902), 
            .CO(n25680));
    SB_LUT4 add_684_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n25678), .O(n2906[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_2 (.CI(n25678), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n25679));
    SB_CARRY add_684_1 (.CI(GND_net), .I0(n2902), .I1(n2902), .CO(n25678));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1097_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2902));   // quad.v(37[5] 40[8])
    defparam i1097_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_684_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2902), 
            .I3(n25701), .O(n2906[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_684_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2902), 
            .I3(n25700), .O(n2906[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_24 (.CI(n25700), .I0(encoder0_position[22]), .I1(n2902), 
            .CO(n25701));
    SB_LUT4 add_684_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2902), 
            .I3(n25699), .O(n2906[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_23 (.CI(n25699), .I0(encoder0_position[21]), .I1(n2902), 
            .CO(n25700));
    SB_LUT4 add_684_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2902), 
            .I3(n25698), .O(n2906[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_22 (.CI(n25698), .I0(encoder0_position[20]), .I1(n2902), 
            .CO(n25699));
    SB_LUT4 add_684_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2902), 
            .I3(n25697), .O(n2906[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_21 (.CI(n25697), .I0(encoder0_position[19]), .I1(n2902), 
            .CO(n25698));
    SB_LUT4 add_684_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2902), 
            .I3(n25696), .O(n2906[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_20 (.CI(n25696), .I0(encoder0_position[18]), .I1(n2902), 
            .CO(n25697));
    SB_LUT4 add_684_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2902), 
            .I3(n25695), .O(n2906[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_19 (.CI(n25695), .I0(encoder0_position[17]), .I1(n2902), 
            .CO(n25696));
    SB_LUT4 add_684_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2902), 
            .I3(n25694), .O(n2906[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_18 (.CI(n25694), .I0(encoder0_position[16]), .I1(n2902), 
            .CO(n25695));
    SB_LUT4 add_684_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2902), 
            .I3(n25693), .O(n2906[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_684_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_684_17 (.CI(n25693), .I0(encoder0_position[15]), .I1(n2902), 
            .CO(n25694));
    \grp_debouncer(2,100)_U0  debounce (.GND_net(GND_net), .VCC_net(VCC_net), 
            .reg_B({reg_B}), .clk32MHz(clk32MHz), .n32962(n32962), .ENCODER0_B_c_0(ENCODER0_B_c_0), 
            .n18541(n18541), .data_o({data_o}), .n18057(n18057), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (GND_net, VCC_net, reg_B, clk32MHz, 
            n32962, ENCODER0_B_c_0, n18541, data_o, n18057, ENCODER0_A_c_1);
    input GND_net;
    input VCC_net;
    output [1:0]reg_B;
    input clk32MHz;
    output n32962;
    input ENCODER0_B_c_0;
    input n18541;
    output [1:0]data_o;
    input n18057;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]n33;
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n26324, n26325, n26323;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n12, n2, cnt_next_6__N_3647, n26326, n26328, n26327;
    
    SB_LUT4 cnt_reg_1467_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n26324), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1467_add_4_4 (.CI(n26324), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n26325));
    SB_LUT4 cnt_reg_1467_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n26323), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1467_add_4_3 (.CI(n26323), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n26324));
    SB_LUT4 cnt_reg_1467_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1467_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n26323));
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[4]), .I3(cnt_reg[2]), 
            .O(n32962));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n32962), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_CARRY cnt_reg_1467_add_4_5 (.CI(n26325), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n26326));
    SB_LUT4 cnt_reg_1467_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n26328), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1467_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n26327), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1467_add_4_7 (.CI(n26327), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n26328));
    SB_LUT4 cnt_reg_1467_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n26326), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1467_add_4_6 (.CI(n26326), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n26327));
    SB_LUT4 cnt_reg_1467_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n26325), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1467_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR cnt_reg_1467__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18541));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18057));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1467__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1467__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1467__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1467__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1467__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1467__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (GND_net, clk32MHz, \state[1] , n29331, n17813, n31208, 
            VCC_net, timer, \neo_pixel_transmitter.t0 , neopxl_color, 
            LED_c, \state_3__N_319[1] , n18064, n18060, n18575, n18574, 
            n18573, n18572, n18571, n18570, n18569, n18568, n18567, 
            n18566, n18565, n18564, n18563, n18562, n18561, n18560, 
            n18559, n18558, n18557, n18556, n18555, n18554, n18553, 
            n18552, n18551, n18550, n18549, n18548, n18547, n18546, 
            n18545, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk32MHz;
    output \state[1] ;
    output n29331;
    output n17813;
    output n31208;
    input VCC_net;
    output [31:0]timer;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input [23:0]neopxl_color;
    input LED_c;
    output \state_3__N_319[1] ;
    input n18064;
    input n18060;
    input n18575;
    input n18574;
    input n18573;
    input n18572;
    input n18571;
    input n18570;
    input n18569;
    input n18568;
    input n18567;
    input n18566;
    input n18565;
    input n18564;
    input n18563;
    input n18562;
    input n18561;
    input n18560;
    input n18559;
    input n18558;
    input n18557;
    input n18556;
    input n18555;
    input n18554;
    input n18553;
    input n18552;
    input n18551;
    input n18550;
    input n18549;
    input n18548;
    input n18547;
    input n18546;
    input n18545;
    output NEOPXL_c;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n26355, n2793, n2819, n26356, n2;
    wire [31:0]n971;
    
    wire n1007, n3102, n3100, n36, n3099, n3107, n3094, n3105, 
        n46, n3089, n3093, n3085, n3095, n42, n3084, n3096, 
        n3083, n3103, n44, n2893, n2794, n26354, n2894, n2795, 
        n26353, \neo_pixel_transmitter.done_N_527 , n35736, \neo_pixel_transmitter.done , 
        n3097;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n3109, n31, n3091, n3092, n50, start_N_518, n7, start, 
        n3087, n3101, n3104, n48, n3106, n3086, n49, n3108, 
        n3088, n3090, n3098, n47, n3116, n3017, n35426, n35423;
    wire [31:0]n255;
    
    wire n17772, n17985, n2895, n2796, n26352, n2984, n2885, n2918, 
        n26307, n2985, n2886, n26306, n1006, n1928, n35434, n16468, 
        n31237, n27197;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n31346, n7_adj_4634, n31372, n16534, n2986, n2887, n26305, 
        n2987, n2888, n26304, n1895, n1902, n1899, n1897, n26, 
        n1907, n1909, n19, n2999, n3009, n30, n3008, n2988, 
        n42_adj_4635, n2990, n2998, n3004, n2995, n40, n3000, 
        n2996, n2993, n45, n1908, n1900, n16, n2992, n2994, 
        n3005, n44_adj_4636, n1904, n1901, n1906, n1898, n24, 
        n2997, n3007, n3006, n2989, n43, n1905, n1903, n28, 
        n3003, n2991, n47_adj_4637, n3002, n3001, n49_adj_4638, 
        n1896, n1829, n35433, n25, n27, n26_adj_4639, n28_adj_4640, 
        n37, n906, n1005, n2889, n26303, n608, n708, n31212, 
        n22673, n739, n15144, n27721, n31167, n807, n838, n60, 
        n905, n31210, n33145, n17881, n15162, n1009, n1008, n33157, 
        n6, n1037, n4, n2890, n26302, n2891, n26301, n2892, 
        n26300, n26299, n26298, n2896, n2797, n26351, n26297, 
        n26296, n2897, n26295, n22763, n1053, n14233, n2898, n26294, 
        n2899, n26293, n2900, n26292, n2901, n26291, n2798, n26350, 
        n2902, n26290, n1806, n1803, n1798, n1805, n24_adj_4641, 
        n1808, n1804, n1802, n1807, n22, n1800, n1799, n1797, 
        n1801, n23, n1796, n1809, n21, n1730, n35432, n1699, 
        n1709, n17, n1698, n1707, n1703, n1705, n21_adj_4642, 
        n1704, n1701, n1708, n20, n1702, n1697, n24_adj_4643, 
        n1700, n1706, n1631, n35431, n2903, n26289, n2904, n26288, 
        n2905, n26287, n2906, n26286, n2907, n26285, n2908, n26284, 
        n2909, n35424, n26283, n2799, n26349, n29, n36_adj_4644, 
        n30_adj_4645, n16589, n2800, n26348, n1608, n1606, n1604, 
        n1603, n20_adj_4646, n1602, n1609, n13, n1598, n1600, 
        n18, n1605, n1599, n22_adj_4647, n1601, n1607, n1334, 
        n35430, n31233, n2801, n26347, n2802, n26346, n1304, n1305, 
        n10, n1303, n1309, n12, n1306, n1308, n1302, n16_adj_4648, 
        n1307, n1301;
    wire [31:0]n133;
    
    wire n26251, n26250, n26249;
    wire [31:0]n1;
    
    wire n27382, n27729, n30476;
    wire [31:0]one_wire_N_470;
    
    wire n27418, n111, n116, n16_adj_4650, n18_adj_4651, n9, n26248, 
        n26247, n26246, n26245, n26244, n26243, n2803, n26345, 
        n26242, n26241, n26240, n2720, n35445, n26239, n26238, 
        n2804, n26344, n26237, n25527, n26236, n26235, n26234, 
        n26233, n26232, n26231, n2693, n2704, n28_adj_4661, n2805, 
        n26343, n26230, n26229, n26228, n2699, n2706, n2694, n2691, 
        n38, n26227, n26226, n26225, n26224, n2709, n22793, n2701, 
        n2696, n2697, n36_adj_4662, n2700, n2705, n42_adj_4663, 
        n2702, n2690, n2689, n2708, n40_adj_4664, n2687, n2703, 
        n2695, n41, n2688, n2698, n2692, n2707, n39, n26223, 
        n2806, n26342, n26222, n25519, n1103, n25642, n1104, n25641, 
        n2807, n26341, n1235, n35444, n26221, n26220, n26219, 
        n1205, n1208, n1202, n1206, n14, n26218, n1207, n1209, 
        n9_adj_4665, n26217, n26216, n26215, n26214, n1105, n25640, 
        n25528, n1203, n1204, n2621, n35443, n26213, n26212, n25547, 
        n26211, n26210, n26209, n26208, n2808, n26340, n26207, 
        n2809, n26339, n26206, n26205, n26204, n26203, n26202, 
        n26201, n25546, n26200, n26199, n26198, n25545, n26197, 
        n26196, n26195, n63, n26194, n61, n26193, n59, n26192, 
        n57, n26191, n55, n26190, n1106, n25639, n53, n26189, 
        n51, n26188, n49_adj_4666, n26187, n47_adj_4668, n26186, 
        n1107, n25638, n45_adj_4669, n26185, n43_adj_4670, n26184, 
        n41_adj_4671, n26183, n39_adj_4673, n26182, n2591, n2608, 
        n2601, n2605, n36_adj_4674, n2606, n2609, n25_adj_4676, 
        n2593, n2596, n2600, n2590, n34, n2594, n2589, n40_adj_4677, 
        n2602, n2588, n2604, n2607, n38_adj_4678, n2598, n2603, 
        n39_adj_4679, n37_adj_4680, n26181, n2592, n2597, n2595, 
        n2599, n37_adj_4681, n35, n26180, n33_adj_4682, n26179, 
        n2522, n35442, n31_adj_4684, n26178, n29_adj_4685, n26177, 
        n27_adj_4687, n26176, n25_adj_4688, n26175, n2491, n2504, 
        n24_adj_4689, n2496, n2505, n2500, n2499, n34_adj_4690, 
        n2497, n2509, n22_adj_4691, n1108, n35427, n25637, n23_adj_4692, 
        n26174, n21_adj_4693, n26173, n2490, n2494, n38_adj_4694, 
        n1109, n19_adj_4695, n26172, n17_adj_4696, n26171, n15, 
        n26170, n13_adj_4697, n26169, n11, n35428, n26168, n3209, 
        n22_adj_4698, n25801, n1136, n26167, n26166, n26165, n26164, 
        n26163, n2501, n2502, n2506, n2492, n36_adj_4700, n26162, 
        n25526, n2495, n2498, n2493, n37_adj_4701, n25800, n35429, 
        n26161, n2507, n2508, n2503, n2489, n35_adj_4702, n25799, 
        n25798, n21_adj_4705, n25797, n25796, n25795, n25520, n25794, 
        n25544, n25525, n2423, n35441, n25543, n25518, n25524, 
        n25542, n25793, n25792, n25541, n25540, n2404, n2407, 
        n22_adj_4715, n2400, n2397, n2402, n2393, n32_adj_4716, 
        n2409, n22787, n2391, n2398, n36_adj_4717, n25791, n2392, 
        n2396, n2390, n2408, n34_adj_4718, n2405, n2406, n2399, 
        n35_adj_4719, n2401, n2403, n2394, n2395, n33_adj_4720, 
        n25790, n25539, n24_adj_4721, n25789, n25788, n33_adj_4722, 
        n41_adj_4723, n38_adj_4724, n43_adj_4725, n40_adj_4726, n46_adj_4727, 
        n39_adj_4728, n47_adj_4729, n23_adj_4730, n25787, n2324, n35440, 
        n25786, n25785, n25784, n25783, n25782, n25781, n25780, 
        n25779, n25538, n25778, n25537, n25523, n25777, n25776, 
        n25775, n25774, n35597, n33265, n35591, n33268, n2302, 
        n2292, n22_adj_4731, n2299, n2309, n30_adj_4732, n35585, 
        n33271, n2294, n2306, n2297, n34_adj_4733, n25517, n2301, 
        n2307, n2291, n2305, n32_adj_4734, n2298, n2295, n2304, 
        n2300, n33_adj_4735, n25773, n2308, n2296, n2303, n2293, 
        n31_adj_4736, n25772, n46_adj_4737, n44_adj_4738, n35537, 
        n35540, n45_adj_4739, n35531, n35534, n43_adj_4740, n25522, 
        n2225, n35439, n25536, n25771, n4_adj_4741, n42_adj_4742, 
        n35519, n40_adj_4743, n34700, n48_adj_4744, n25535, n1400, 
        n25967, n1401, n25966, n52, n1402, n25965, n25534, n1403, 
        n25964, n25521, n25533, n1404, n25963, n1405, n25962, 
        n1406, n25961, n1407, n25960, n34034, n1408, n25959, n1409, 
        n34387, n34388, n33056, n25532, n26604, n26603, n26602, 
        n26601, n26600, n2193, n2194, n2206, n2204, n28_adj_4745, 
        n26599, n26598, n26597, n2203, n2209, n32_adj_4746, n2208, 
        n2201, n2192, n2196, n30_adj_4747, n26596, n2195, n2207, 
        n2205, n2199, n31_adj_4748, n2202, n2197, n2198, n2200, 
        n29_adj_4749, n26595, n26594, n26593, n26592, n26591, n26590, 
        n26589, n26588, n26587, n26586, n26585, n26584, n26583, 
        n26582, n26581, n26580, n26579, n26578, n26577, n25531, 
        n26576, n26575, n26574, n26573, n26572, n26571, n26570, 
        n26569, n2126, n35437, n51_adj_4750, n26568, n26567, n26566, 
        n1994, n26565, n1995, n26564, n1996, n26563, n1997, n26562, 
        n1998, n26561, n1999, n26560, n2000, n26559, n2001, n26558, 
        n2002, n26557, n2003, n26556, n25530, n25529, n2004, n26555, 
        n2005, n26554, n2006, n26553, n2007, n26552, n2008, n26551, 
        n2009, n2093, n2027, n26550;
    wire [3:0]state_3__N_319;
    
    wire n2094, n26549, n2095, n26548, n2096, n26547, n22097, 
        n12_adj_4751, n2786, n40_adj_4752, n2788, n38_adj_4753, n2787, 
        n39_adj_4754, n2790, n37_adj_4755, n34_adj_4756, n2789, n2792, 
        n42_adj_4757, n46_adj_4758, n2791, n33_adj_4759, n1039, n1499, 
        n1433, n25881, n1500, n25880, n1501, n25879, n1502, n25878, 
        n1503, n25877, n1504, n25876, n22737, n2097, n26546, n1505, 
        n25875, n2098, n26545, n2099, n26544, n2100, n26543, n1506, 
        n25874, n2101, n26542, n1507, n25873, n2102, n26541, n2103, 
        n26540, n2104, n26539, n2105, n26538, n2106, n26537, n2107, 
        n26536, n2108, n35435, n26535, n2109, n26534, n26533, 
        n26532, n1508, n35436, n25872, n1509, n1532, n35438, n25871, 
        n25870, n25869, n25868, n25867, \neo_pixel_transmitter.done_N_533 , 
        n31384, n25866, n26531, n26530, n25865, n26529, n25864, 
        n26528, n25863, n25862, n25861, n26527, n4820, n25860, 
        n26526, n26525, n26524, n26523, n26522, n26521, n26520, 
        n25859, n26519, n26518, n26517, n34056, n26516, n26515, 
        n31350, n26514, n26513, n26512, n26511, n25858, n26510, 
        n26509, n26508, n26507, n26506, n26505, n26504, n26503, 
        n26502, n25857, n26501, n25856, n26500, n26499, n26498, 
        n18_adj_4760, n26497, n26496, n26495, n26494, n26493, n26492, 
        n20_adj_4761, n26491, n15_adj_4762, n26490, n26489, n26488, 
        n26487, n26486, n26485, n26484, n26483, n26482, n26481, 
        n18_adj_4763, n26480, n22779, n26479, n26478, n26477, n26476, 
        n26475, n26474, n26473, n30_adj_4764, n26472, n26471, n28_adj_4765, 
        n26470, n29_adj_4766, n26469, n26468, n26467, n26466, n26465, 
        n26464, n26463, n27_adj_4767, n26462, n26461, n26436, n26435, 
        n26434, n26433, n26432, n26431, n26430, n26429, n26428, 
        n26427, n26426, n26425, n26424, n26423, n26422, n26421, 
        n26420, n26419, n26418, n26417, n26416, n26415, n26414, 
        n26413, n26412, n26411, n26410, n26409, n26408, n26407, 
        n26406, n26405, n26404, n26403, n26402, n26401, n26400, 
        n26399, n26398, n26397, n26396, n26395, n26394, n26393, 
        n26392, n26391, n26390, n26389, n26388, n26387, n26386, 
        n26385, n26384, n26383, n26382, n26381, n26380, n26379, 
        n26378, n26377, n26376, n26375, n26374, n26373, n26372, 
        n26371, n26370, n26369, n26368, n26367, n26366, n26365, 
        n26364, n26363, n26362, n26361, n26360, n26359, n26358, 
        n26357, n22815, n16_adj_4768, n17_adj_4769, n35447, n35450, 
        n14_adj_4770, n33986, n31304, n14_adj_4771, n13_adj_4772, 
        n20_adj_4773, n19_adj_4774, n6_adj_4775, n32361, n32_adj_4776, 
        n30_adj_4777, n31_adj_4778, n29_adj_4779;
    wire [4:0]color_bit_N_513;
    
    wire n34030, n18_adj_4780, n28_adj_4781, n26_adj_4782, n27_adj_4783, 
        n25_adj_4784;
    
    SB_CARRY mod_5_add_1942_19 (.CI(n26355), .I0(n2793), .I1(n2819), .CO(n26356));
    SB_LUT4 i28801_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i28801_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i9_2_lut (.I0(n3102), .I1(n3100), .I2(GND_net), .I3(GND_net), 
            .O(n36));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut (.I0(n3099), .I1(n3107), .I2(n3094), .I3(n3105), 
            .O(n46));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n3089), .I1(n3093), .I2(n3085), .I3(n3095), 
            .O(n42));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n3084), .I1(n3096), .I2(n3083), .I3(n3103), 
            .O(n44));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n26354), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n26354), .I0(n2794), .I1(n2819), .CO(n26355));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n26353), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n35736), .D(\neo_pixel_transmitter.done_N_527 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i4_3_lut (.I0(n3097), .I1(bit_ctr[4]), .I2(n3109), .I3(GND_net), 
            .O(n31));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i23_4_lut (.I0(n3091), .I1(n46), .I2(n36), .I3(n3092), .O(n50));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(n7), .D(start_N_518));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i21_4_lut (.I0(n3087), .I1(n42), .I2(n3101), .I3(n3104), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n31), .I1(n44), .I2(n3106), .I3(n3086), .O(n49));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n3108), .I1(n3088), .I2(n3090), .I3(n3098), 
            .O(n47));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n47), .I1(n49), .I2(n48), .I3(n50), .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29254_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35426));
    defparam i29254_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29251_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35423));
    defparam i29251_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n17772), 
            .D(n255[18]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n17772), 
            .D(n255[17]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n17772), 
            .D(n255[16]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n17772), 
            .D(n255[15]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n17772), 
            .D(n255[14]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n17772), 
            .D(n255[13]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n17772), 
            .D(n255[12]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n17772), 
            .D(n255[11]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n17772), 
            .D(n255[10]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n17772), 
            .D(n255[9]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n17772), 
            .D(n255[8]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n17772), 
            .D(n255[7]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n17772), 
            .D(n255[6]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n17772), 
            .D(n255[5]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n17772), 
            .D(n255[4]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n17772), 
            .D(n255[3]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n17772), 
            .D(n255[2]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n17772), 
            .D(n255[1]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n17772), 
            .D(n255[25]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n17772), 
            .D(n255[24]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n17772), 
            .D(n255[27]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_17 (.CI(n26353), .I0(n2795), .I1(n2819), .CO(n26354));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n26352), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n26307), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n26306), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28799_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i28799_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i29262_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35434));
    defparam i29262_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25182_4_lut (.I0(n16468), .I1(n31237), .I2(n27197), .I3(state[0]), 
            .O(n31346));
    defparam i25182_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut_adj_1494 (.I0(n31346), .I1(\state[1] ), .I2(start), 
            .I3(\neo_pixel_transmitter.done ), .O(n7_adj_4634));
    defparam i20_4_lut_adj_1494.LUT_INIT = 16'hcfcd;
    SB_LUT4 i1_4_lut (.I0(n31372), .I1(n7_adj_4634), .I2(n16534), .I3(\state[1] ), 
            .O(n29331));
    defparam i1_4_lut.LUT_INIT = 16'hccc4;
    SB_CARRY mod_5_add_2009_26 (.CI(n26306), .I0(n2886), .I1(n2918), .CO(n26307));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n26305), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n26305), .I0(n2887), .I1(n2918), .CO(n26306));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n26304), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1495 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19));
    defparam i4_3_lut_adj_1495.LUT_INIT = 16'heaea;
    SB_LUT4 i4_3_lut_adj_1496 (.I0(n2999), .I1(bit_ctr[5]), .I2(n3009), 
            .I3(GND_net), .O(n30));
    defparam i4_3_lut_adj_1496.LUT_INIT = 16'heaea;
    SB_LUT4 i16_4_lut (.I0(n2986), .I1(n3008), .I2(n2988), .I3(n2987), 
            .O(n42_adj_4635));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2990), .I1(n2998), .I2(n3004), .I3(n2995), 
            .O(n40));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1497 (.I0(n2985), .I1(n3000), .I2(n2996), .I3(n2993), 
            .O(n45));
    defparam i19_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut (.I0(n2992), .I1(n2994), .I2(n3005), .I3(n2984), 
            .O(n44_adj_4636));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1498 (.I0(n2997), .I1(n3007), .I2(n3006), .I3(n2989), 
            .O(n43));
    defparam i17_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n19), .I1(n26), .I2(n1905), .I3(n1903), .O(n28));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1499 (.I0(n3003), .I1(n42_adj_4635), .I2(n30), 
            .I3(n2991), .O(n47_adj_4637));
    defparam i21_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1500 (.I0(n45), .I1(n3002), .I2(n40), .I3(n3001), 
            .O(n49_adj_4638));
    defparam i23_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_adj_4638), .I1(n47_adj_4637), .I2(n43), 
            .I3(n44_adj_4636), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1501 (.I0(n1896), .I1(n28), .I2(n24), .I3(n16), 
            .O(n1928));
    defparam i14_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i29261_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35433));
    defparam i29261_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_24 (.CI(n26304), .I0(n2888), .I1(n2918), .CO(n26305));
    SB_LUT4 i17_4_lut_adj_1502 (.I0(n25), .I1(n27), .I2(n26_adj_4639), 
            .I3(n28_adj_4640), .O(n37));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n26303), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n26303), .I0(n2889), .I1(n2918), .CO(n26304));
    SB_LUT4 i18088_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i18088_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n31212), .I3(n22673), 
            .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n15144));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i28146_3_lut (.I0(n27721), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n31167));
    defparam i28146_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n31212), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i26973_3_lut (.I0(n906), .I1(n905), .I2(n31210), .I3(GND_net), 
            .O(n33145));
    defparam i26973_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n17881), .I1(n33145), .I2(bit_ctr[26]), .I3(n15162), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 i1_2_lut_adj_1504 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n15162));
    defparam i1_2_lut_adj_1504.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n15162), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26985_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n33157));
    defparam i26985_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n2), .I1(n6), .I2(n1005), .I3(n33157), .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i28811_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(22[26:36])
    defparam i28811_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n26302), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n26302), .I0(n2890), .I1(n2918), .CO(n26303));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n26301), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n26301), .I0(n2891), .I1(n2918), .CO(n26302));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n26300), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n26300), .I0(n2892), .I1(n2918), .CO(n26301));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n26299), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n26299), .I0(n2893), .I1(n2918), .CO(n26300));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n26298), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n26298), .I0(n2894), .I1(n2918), .CO(n26299));
    SB_CARRY mod_5_add_1942_16 (.CI(n26352), .I0(n2796), .I1(n2819), .CO(n26353));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n26351), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n26297), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n26297), .I0(n2895), .I1(n2918), .CO(n26298));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n26296), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n26296), .I0(n2896), .I1(n2918), .CO(n26297));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n26295), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i255_2_lut (.I0(n22763), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1053));   // verilog/neopixel.v(103[9] 111[12])
    defparam i255_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1505 (.I0(state[0]), .I1(n14233), .I2(n1053), 
            .I3(\state[1] ), .O(n17813));
    defparam i1_4_lut_adj_1505.LUT_INIT = 16'haf33;
    SB_LUT4 i15_4_lut_adj_1506 (.I0(n14233), .I1(n1053), .I2(\state[1] ), 
            .I3(state[0]), .O(n31208));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1506.LUT_INIT = 16'h0535;
    SB_CARRY mod_5_add_2009_15 (.CI(n26295), .I0(n2897), .I1(n2918), .CO(n26296));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n26294), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n26294), .I0(n2898), .I1(n2918), .CO(n26295));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n26293), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n26351), .I0(n2797), .I1(n2819), .CO(n26352));
    SB_CARRY mod_5_add_2009_13 (.CI(n26293), .I0(n2899), .I1(n2918), .CO(n26294));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n26292), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n26292), .I0(n2900), .I1(n2918), .CO(n26293));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n26291), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n26350), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n26291), .I0(n2901), .I1(n2918), .CO(n26292));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n26290), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n26290), .I0(n2902), .I1(n2918), .CO(n26291));
    SB_LUT4 i10_4_lut (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4641));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1507 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23));
    defparam i9_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1508 (.I0(n21), .I1(n23), .I2(n22), .I3(n24_adj_4641), 
            .O(n1829));
    defparam i13_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i29260_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35432));
    defparam i29260_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1509 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17));
    defparam i4_3_lut_adj_1509.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1510 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4642));
    defparam i8_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1511 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20));
    defparam i7_3_lut_adj_1511.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1512 (.I0(n21_adj_4642), .I1(n17), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4643));
    defparam i11_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n1700), .I1(n24_adj_4643), .I2(n20), .I3(n1706), 
            .O(n1730));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29259_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35431));
    defparam i29259_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n26289), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n26289), .I0(n2903), .I1(n2918), .CO(n26290));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n26288), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n26288), .I0(n2904), .I1(n2918), .CO(n26289));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n26287), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n26287), .I0(n2905), .I1(n2918), .CO(n26288));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n26286), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n26350), .I0(n2798), .I1(n2819), .CO(n26351));
    SB_CARRY mod_5_add_2009_6 (.CI(n26286), .I0(n2906), .I1(n2918), .CO(n26287));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n26285), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n26285), .I0(n2907), .I1(n2918), .CO(n26286));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n26284), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n26284), .I0(n2908), .I1(n2918), .CO(n26285));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n35424), 
            .I3(n26283), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n26283), .I0(n2909), .I1(n35424), .CO(n26284));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n35424), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n35424), 
            .CO(n26283));
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n17772), 
            .D(n255[21]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n17772), 
            .D(n255[20]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n26349), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19_4_lut_adj_1513 (.I0(n37), .I1(n29), .I2(n36_adj_4644), 
            .I3(n30_adj_4645), .O(n16589));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_13 (.CI(n26349), .I0(n2799), .I1(n2819), .CO(n26350));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n26348), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i8_4_lut_adj_1514 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4646));
    defparam i8_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), .I3(GND_net), 
            .O(n13));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1515 (.I0(n13), .I1(n20_adj_4646), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4647));
    defparam i10_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1516 (.I0(n1601), .I1(n22_adj_4647), .I2(n18), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n17772), 
            .D(n255[19]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_12 (.CI(n26348), .I0(n2800), .I1(n2819), .CO(n26349));
    SB_LUT4 i29258_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35430));
    defparam i29258_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25075_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n31233));
    defparam i25075_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n26347), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n26347), .I0(n2801), .I1(n2819), .CO(n26348));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n26346), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10));
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10), 
            .O(n16_adj_4648));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1518 (.I0(n1307), .I1(n16_adj_4648), .I2(n12), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1461_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n26251), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1461_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n26250), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n17772), 
            .D(n255[23]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1461_add_4_32 (.CI(n26250), .I0(GND_net), .I1(timer[30]), 
            .CO(n26251));
    SB_LUT4 timer_1461_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n26249), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(bit_ctr[3]), .I1(n27382), .I2(GND_net), 
            .I3(GND_net), .O(n27729));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1461_add_4_31 (.CI(n26249), .I0(GND_net), .I1(timer[29]), 
            .CO(n26250));
    SB_LUT4 i28750_2_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n30476));
    defparam i28750_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1520 (.I0(one_wire_N_470[4]), .I1(one_wire_N_470[3]), 
            .I2(n30476), .I3(n27418), .O(n111));
    defparam i1_4_lut_adj_1520.LUT_INIT = 16'h5155;
    SB_LUT4 i1_4_lut_adj_1521 (.I0(n111), .I1(n30476), .I2(one_wire_N_470[2]), 
            .I3(one_wire_N_470[3]), .O(n116));
    defparam i1_4_lut_adj_1521.LUT_INIT = 16'haeee;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_470[8]), .I1(one_wire_N_470[10]), .I2(n31233), 
            .I3(n116), .O(n16_adj_4650));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i8_3_lut (.I0(one_wire_N_470[5]), .I1(n16_adj_4650), .I2(n16589), 
            .I3(GND_net), .O(n18_adj_4651));
    defparam i8_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3_4_lut_adj_1522 (.I0(n9), .I1(one_wire_N_470[11]), .I2(n18_adj_4651), 
            .I3(one_wire_N_470[7]), .O(n35736));
    defparam i3_4_lut_adj_1522.LUT_INIT = 16'hffef;
    SB_LUT4 mux_724_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_527 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_724_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 timer_1461_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n26248), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_30 (.CI(n26248), .I0(GND_net), .I1(timer[28]), 
            .CO(n26249));
    SB_LUT4 timer_1461_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n26247), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_29 (.CI(n26247), .I0(GND_net), .I1(timer[27]), 
            .CO(n26248));
    SB_LUT4 timer_1461_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n26246), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_10 (.CI(n26346), .I0(n2802), .I1(n2819), .CO(n26347));
    SB_CARRY timer_1461_add_4_28 (.CI(n26246), .I0(GND_net), .I1(timer[26]), 
            .CO(n26247));
    SB_LUT4 timer_1461_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n26245), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_27 (.CI(n26245), .I0(GND_net), .I1(timer[25]), 
            .CO(n26246));
    SB_LUT4 timer_1461_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n26244), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_26 (.CI(n26244), .I0(GND_net), .I1(timer[24]), 
            .CO(n26245));
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1461_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n26243), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n26345), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1461_add_4_25 (.CI(n26243), .I0(GND_net), .I1(timer[23]), 
            .CO(n26244));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1461_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n26242), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1461_add_4_24 (.CI(n26242), .I0(GND_net), .I1(timer[22]), 
            .CO(n26243));
    SB_LUT4 timer_1461_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n26241), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_23 (.CI(n26241), .I0(GND_net), .I1(timer[21]), 
            .CO(n26242));
    SB_LUT4 timer_1461_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n26240), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_22 (.CI(n26240), .I0(GND_net), .I1(timer[20]), 
            .CO(n26241));
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_9 (.CI(n26345), .I0(n2803), .I1(n2819), .CO(n26346));
    SB_LUT4 i29273_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35445));
    defparam i29273_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1461_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n26239), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_21 (.CI(n26239), .I0(GND_net), .I1(timer[19]), 
            .CO(n26240));
    SB_LUT4 timer_1461_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n26238), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_20 (.CI(n26238), .I0(GND_net), .I1(timer[18]), 
            .CO(n26239));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n26344), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1461_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n26237), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_8 (.CI(n26344), .I0(n2804), .I1(n2819), .CO(n26345));
    SB_CARRY timer_1461_add_4_19 (.CI(n26237), .I0(GND_net), .I1(timer[17]), 
            .CO(n26238));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n25527), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1461_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n26236), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_18 (.CI(n26236), .I0(GND_net), .I1(timer[16]), 
            .CO(n26237));
    SB_LUT4 timer_1461_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n26235), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_17 (.CI(n26235), .I0(GND_net), .I1(timer[15]), 
            .CO(n26236));
    SB_LUT4 timer_1461_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n26234), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_16 (.CI(n26234), .I0(GND_net), .I1(timer[14]), 
            .CO(n26235));
    SB_LUT4 timer_1461_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n26233), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_15 (.CI(n26233), .I0(GND_net), .I1(timer[13]), 
            .CO(n26234));
    SB_LUT4 timer_1461_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n26232), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_14 (.CI(n26232), .I0(GND_net), .I1(timer[12]), 
            .CO(n26233));
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1461_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n26231), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1461_add_4_13 (.CI(n26231), .I0(GND_net), .I1(timer[11]), 
            .CO(n26232));
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4661));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n26343), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1461_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n26230), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_12 (.CI(n26230), .I0(GND_net), .I1(timer[10]), 
            .CO(n26231));
    SB_LUT4 timer_1461_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n26229), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_11 (.CI(n26229), .I0(GND_net), .I1(timer[9]), 
            .CO(n26230));
    SB_LUT4 timer_1461_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n26228), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_10 (.CI(n26228), .I0(GND_net), .I1(timer[8]), 
            .CO(n26229));
    SB_LUT4 i15_4_lut_adj_1523 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1461_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n26227), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_9 (.CI(n26227), .I0(GND_net), .I1(timer[7]), 
            .CO(n26228));
    SB_LUT4 timer_1461_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n26226), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_8 (.CI(n26226), .I0(GND_net), .I1(timer[6]), 
            .CO(n26227));
    SB_LUT4 timer_1461_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n26225), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_7 (.CI(n26225), .I0(GND_net), .I1(timer[5]), 
            .CO(n26226));
    SB_LUT4 timer_1461_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n26224), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18216_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n22793));
    defparam i18216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1942_7 (.CI(n26343), .I0(n2805), .I1(n2819), .CO(n26344));
    SB_CARRY timer_1461_add_4_6 (.CI(n26224), .I0(GND_net), .I1(timer[4]), 
            .CO(n26225));
    SB_LUT4 i13_4_lut_adj_1524 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n22793), 
            .O(n36_adj_4662));
    defparam i13_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1525 (.I0(n2700), .I1(n38), .I2(n28_adj_4661), 
            .I3(n2705), .O(n42_adj_4663));
    defparam i19_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1526 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4664));
    defparam i17_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1527 (.I0(n2687), .I1(n36_adj_4662), .I2(n2703), 
            .I3(n2695), .O(n41));
    defparam i18_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1528 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39));
    defparam i16_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1461_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n26223), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n26342), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1461_add_4_5 (.CI(n26223), .I0(GND_net), .I1(timer[3]), 
            .CO(n26224));
    SB_LUT4 i22_4_lut_adj_1529 (.I0(n39), .I1(n41), .I2(n40_adj_4664), 
            .I3(n42_adj_4663), .O(n2720));
    defparam i22_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1942_6 (.CI(n26342), .I0(n2806), .I1(n2819), .CO(n26343));
    SB_LUT4 timer_1461_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n26222), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n25519), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4), .I1(n4), .I2(n1037), .I3(n25642), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n25641), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n26341), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i29272_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35444));
    defparam i29272_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1461_add_4_4 (.CI(n26222), .I0(GND_net), .I1(timer[2]), 
            .CO(n26223));
    SB_LUT4 timer_1461_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n26221), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_3 (.CI(n26221), .I0(GND_net), .I1(timer[1]), 
            .CO(n26222));
    SB_LUT4 timer_1461_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1461_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1461_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n26221));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n26220), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n26219), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1530 (.I0(n1205), .I1(n1208), .I2(n1202), .I3(n1206), 
            .O(n14));
    defparam i6_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_27 (.CI(n26219), .I0(n2985), .I1(n3017), .CO(n26220));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n26218), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n26218), .I0(n2986), .I1(n3017), .CO(n26219));
    SB_CARRY mod_5_add_1942_5 (.CI(n26341), .I0(n2807), .I1(n2819), .CO(n26342));
    SB_LUT4 i1_3_lut_adj_1531 (.I0(bit_ctr[23]), .I1(n1207), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4665));
    defparam i1_3_lut_adj_1531.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n26217), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n26217), .I0(n2987), .I1(n3017), .CO(n26218));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n26216), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n26216), .I0(n2988), .I1(n3017), .CO(n26217));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n26215), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n26215), .I0(n2989), .I1(n3017), .CO(n26216));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n26214), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n25641), .I0(n1005), .I1(n1037), .CO(n25642));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n25640), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n25527), .I0(bit_ctr[11]), .I1(GND_net), .CO(n25528));
    SB_LUT4 i7_4_lut_adj_1532 (.I0(n9_adj_4665), .I1(n14), .I2(n1203), 
            .I3(n1204), .O(n1235));
    defparam i7_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i29271_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35443));
    defparam i29271_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_736_6 (.CI(n25640), .I0(n1006), .I1(n1037), .CO(n25641));
    SB_CARRY mod_5_add_2076_22 (.CI(n26214), .I0(n2990), .I1(n3017), .CO(n26215));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n26213), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n26213), .I0(n2991), .I1(n3017), .CO(n26214));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n26212), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n26212), .I0(n2992), .I1(n3017), .CO(n26213));
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n25547), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n26211), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n26211), .I0(n2993), .I1(n3017), .CO(n26212));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n26210), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n26210), .I0(n2994), .I1(n3017), .CO(n26211));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n26209), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n26209), .I0(n2995), .I1(n3017), .CO(n26210));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n26208), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n26340), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n26208), .I0(n2996), .I1(n3017), .CO(n26209));
    SB_CARRY mod_5_add_1942_4 (.CI(n26340), .I0(n2808), .I1(n2819), .CO(n26341));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n26207), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n35423), 
            .I3(n26339), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_15 (.CI(n26207), .I0(n2997), .I1(n3017), .CO(n26208));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n26206), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n26206), .I0(n2998), .I1(n3017), .CO(n26207));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n26205), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n26205), .I0(n2999), .I1(n3017), .CO(n26206));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n26204), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n26204), .I0(n3000), .I1(n3017), .CO(n26205));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n26203), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n26203), .I0(n3001), .I1(n3017), .CO(n26204));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n26202), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n26202), .I0(n3002), .I1(n3017), .CO(n26203));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n26201), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n26201), .I0(n3003), .I1(n3017), .CO(n26202));
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n25546), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n26200), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n26200), .I0(n3004), .I1(n3017), .CO(n26201));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n26199), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n26199), .I0(n3005), .I1(n3017), .CO(n26200));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n26198), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n25546), .I0(bit_ctr[30]), .I1(GND_net), .CO(n25547));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n25545), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_6 (.CI(n26198), .I0(n3006), .I1(n3017), .CO(n26199));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n26197), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n26197), .I0(n3007), .I1(n3017), .CO(n26198));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n26196), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n26196), .I0(n3008), .I1(n3017), .CO(n26197));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n35426), 
            .I3(n26195), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n26195), .I0(n3009), .I1(n35426), .CO(n26196));
    SB_CARRY mod_5_add_1942_3 (.CI(n26339), .I0(n2809), .I1(n35423), .CO(n26340));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n35426), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n35423), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n35426), 
            .CO(n26195));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n26194), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n26193), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n35423), 
            .CO(n26339));
    SB_CARRY mod_5_add_2143_28 (.CI(n26193), .I0(n3084), .I1(n3116), .CO(n26194));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n26192), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n26192), .I0(n3085), .I1(n3116), .CO(n26193));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n26191), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n26191), .I0(n3086), .I1(n3116), .CO(n26192));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n26190), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n26190), .I0(n3087), .I1(n3116), .CO(n26191));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n25639), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n26189), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n26189), .I0(n3088), .I1(n3116), .CO(n26190));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n26188), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n26188), .I0(n3089), .I1(n3116), .CO(n26189));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n26187), .O(n49_adj_4666)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n26187), .I0(n3090), .I1(n3116), .CO(n26188));
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n26186), .O(n47_adj_4668)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n26186), .I0(n3091), .I1(n3116), .CO(n26187));
    SB_CARRY mod_5_add_736_5 (.CI(n25639), .I0(n1007), .I1(n1037), .CO(n25640));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n25638), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n26185), .O(n45_adj_4669)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n26185), .I0(n3092), .I1(n3116), .CO(n26186));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n26184), .O(n43_adj_4670)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n26184), .I0(n3093), .I1(n3116), .CO(n26185));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n26183), .O(n41_adj_4671)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n26183), .I0(n3094), .I1(n3116), .CO(n26184));
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n26182), .O(n39_adj_4673)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1533 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4674));
    defparam i14_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_3_lut_adj_1534 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4676));
    defparam i3_3_lut_adj_1534.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_2143_17 (.CI(n26182), .I0(n3095), .I1(n3116), .CO(n26183));
    SB_LUT4 i12_4_lut_adj_1535 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34));
    defparam i12_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1536 (.I0(n25_adj_4676), .I1(n36_adj_4674), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4677));
    defparam i18_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1537 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4678));
    defparam i16_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4679));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n26181), .O(n37_adj_4680)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n17772), 
            .D(n255[0]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i15_4_lut_adj_1538 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4681));
    defparam i15_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1539 (.I0(n37_adj_4681), .I1(n39_adj_4679), .I2(n38_adj_4678), 
            .I3(n40_adj_4677), .O(n2621));
    defparam i21_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_16 (.CI(n26181), .I0(n3096), .I1(n3116), .CO(n26182));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n26180), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n26180), .I0(n3097), .I1(n3116), .CO(n26181));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n26179), .O(n33_adj_4682)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29270_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35442));
    defparam i29270_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_736_4 (.CI(n25638), .I0(n1008), .I1(n1037), .CO(n25639));
    SB_CARRY mod_5_add_2143_14 (.CI(n26179), .I0(n3098), .I1(n3116), .CO(n26180));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n26178), .O(n31_adj_4684)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n26178), .I0(n3099), .I1(n3116), .CO(n26179));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n26177), .O(n29_adj_4685)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n26177), .I0(n3100), .I1(n3116), .CO(n26178));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n26176), .O(n27_adj_4687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n26176), .I0(n3101), .I1(n3116), .CO(n26177));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n26175), .O(n25_adj_4688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4689));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1540 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4690));
    defparam i13_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_10 (.CI(n26175), .I0(n3102), .I1(n3116), .CO(n26176));
    SB_LUT4 i1_3_lut_adj_1541 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4691));
    defparam i1_3_lut_adj_1541.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n35427), 
            .I3(n25637), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n26174), .O(n23_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n26174), .I0(n3103), .I1(n3116), .CO(n26175));
    SB_CARRY mod_5_add_736_3 (.CI(n25637), .I0(n1009), .I1(n35427), .CO(n25638));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n26173), .O(n21_adj_4693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n26173), .I0(n3104), .I1(n3116), .CO(n26174));
    SB_LUT4 i17_4_lut_adj_1542 (.I0(n2490), .I1(n34_adj_4690), .I2(n24_adj_4689), 
            .I3(n2494), .O(n38_adj_4694));
    defparam i17_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n35427), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n26172), .O(n19_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n26172), .I0(n3105), .I1(n3116), .CO(n26173));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n26171), .O(n17_adj_4696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n26171), .I0(n3106), .I1(n3116), .CO(n26172));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n26170), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n26170), .I0(n3107), .I1(n3116), .CO(n26171));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n26169), .O(n13_adj_4697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n26169), .I0(n3108), .I1(n3116), .CO(n26170));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n35428), 
            .I3(n26168), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n26168), .I0(n3109), .I1(n35428), .CO(n26169));
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n35427), 
            .CO(n25637));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n35428), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n35428), 
            .CO(n26168));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_470[22]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n25801), .O(n22_adj_4698)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n26167), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n26166), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n26166), .I0(n1104), .I1(n1136), .CO(n26167));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n26165), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n26165), .I0(n1105), .I1(n1136), .CO(n26166));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n26164), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n26164), .I0(n1106), .I1(n1136), .CO(n26165));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n26163), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1543 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4700));
    defparam i15_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_5 (.CI(n26163), .I0(n1107), .I1(n1136), .CO(n26164));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n26162), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n25526), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1544 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4691), 
            .O(n37_adj_4701));
    defparam i16_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_803_4 (.CI(n26162), .I0(n1108), .I1(n1136), .CO(n26163));
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_470[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n25800), .O(n26_adj_4639)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n35429), 
            .I3(n26161), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n26161), .I0(n1109), .I1(n35429), .CO(n26162));
    SB_CARRY sub_14_add_2_32 (.CI(n25800), .I0(timer[30]), .I1(n1[30]), 
            .CO(n25801));
    SB_LUT4 i14_4_lut_adj_1545 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4702));
    defparam i14_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n35429), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n35429), 
            .CO(n26161));
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20_4_lut_adj_1546 (.I0(n35_adj_4702), .I1(n37_adj_4701), .I2(n36_adj_4700), 
            .I3(n38_adj_4694), .O(n2522));
    defparam i20_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_470[25]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n25799), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n25799), .I0(timer[29]), .I1(n1[29]), 
            .CO(n25800));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_470[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n25798), .O(n28_adj_4640)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n25798), .I0(timer[28]), .I1(n1[28]), 
            .CO(n25799));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_470[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n25797), .O(n21_adj_4705)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n25797), .I0(timer[27]), .I1(n1[27]), 
            .CO(n25798));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n25796), .O(one_wire_N_470[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n25796), .I0(timer[26]), .I1(n1[26]), 
            .CO(n25797));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n25795), .O(one_wire_N_470[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_12 (.CI(n25526), .I0(bit_ctr[10]), .I1(GND_net), .CO(n25527));
    SB_CARRY add_21_5 (.CI(n25519), .I0(bit_ctr[3]), .I1(GND_net), .CO(n25520));
    SB_CARRY sub_14_add_2_27 (.CI(n25795), .I0(timer[25]), .I1(n1[25]), 
            .CO(n25796));
    SB_CARRY add_21_31 (.CI(n25545), .I0(bit_ctr[29]), .I1(GND_net), .CO(n25546));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n25794), .O(one_wire_N_470[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n25544), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n25544), .I0(bit_ctr[28]), .I1(GND_net), .CO(n25545));
    SB_CARRY sub_14_add_2_26 (.CI(n25794), .I0(timer[24]), .I1(n1[24]), 
            .CO(n25795));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n25525), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29269_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35441));
    defparam i29269_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n25543), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n25518), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n17772), 
            .D(n255[22]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_4 (.CI(n25518), .I0(bit_ctr[2]), .I1(GND_net), .CO(n25519));
    SB_CARRY add_21_11 (.CI(n25525), .I0(bit_ctr[9]), .I1(GND_net), .CO(n25526));
    SB_CARRY add_21_29 (.CI(n25543), .I0(bit_ctr[27]), .I1(GND_net), .CO(n25544));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n25524), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n25542), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_470[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n25793), .O(n30_adj_4645)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n25793), .I0(timer[23]), .I1(n1[23]), 
            .CO(n25794));
    SB_CARRY add_21_28 (.CI(n25542), .I0(bit_ctr[26]), .I1(GND_net), .CO(n25543));
    SB_CARRY add_21_10 (.CI(n25524), .I0(bit_ctr[8]), .I1(GND_net), .CO(n25525));
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n25792), .O(one_wire_N_470[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n25541), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n25541), .I0(bit_ctr[25]), .I1(GND_net), .CO(n25542));
    SB_CARRY sub_14_add_2_24 (.CI(n25792), .I0(timer[22]), .I1(n1[22]), 
            .CO(n25793));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n25540), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(n2404), .I1(n2407), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4715));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1547 (.I0(n2400), .I1(n2397), .I2(n2402), .I3(n2393), 
            .O(n32_adj_4716));
    defparam i12_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i18210_2_lut (.I0(bit_ctr[11]), .I1(n2409), .I2(GND_net), 
            .I3(GND_net), .O(n22787));
    defparam i18210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16_4_lut_adj_1548 (.I0(n2391), .I1(n32_adj_4716), .I2(n22_adj_4715), 
            .I3(n2398), .O(n36_adj_4717));
    defparam i16_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_470[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n25791), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i14_4_lut_adj_1549 (.I0(n2392), .I1(n2396), .I2(n2390), .I3(n2408), 
            .O(n34_adj_4718));
    defparam i14_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1550 (.I0(n2405), .I1(n2406), .I2(n22787), .I3(n2399), 
            .O(n35_adj_4719));
    defparam i15_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_23 (.CI(n25791), .I0(timer[21]), .I1(n1[21]), 
            .CO(n25792));
    SB_LUT4 i13_4_lut_adj_1551 (.I0(n2401), .I1(n2403), .I2(n2394), .I3(n2395), 
            .O(n33_adj_4720));
    defparam i13_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_470[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n25790), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i19_4_lut_adj_1552 (.I0(n33_adj_4720), .I1(n35_adj_4719), .I2(n34_adj_4718), 
            .I3(n36_adj_4717), .O(n2423));
    defparam i19_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_26 (.CI(n25540), .I0(bit_ctr[24]), .I1(GND_net), .CO(n25541));
    SB_CARRY sub_14_add_2_22 (.CI(n25790), .I0(timer[20]), .I1(n1[20]), 
            .CO(n25791));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n25539), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_21_lut (.I0(one_wire_N_470[12]), .I1(timer[19]), 
            .I2(n1[19]), .I3(n25789), .O(n24_adj_4721)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n25789), .I0(timer[19]), .I1(n1[19]), 
            .CO(n25790));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n25788), .O(one_wire_N_470[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF timer_1461__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i29252_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35424));
    defparam i29252_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_3_lut_adj_1553 (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), 
            .I3(GND_net), .O(n33_adj_4722));
    defparam i8_3_lut_adj_1553.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1554 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4723));
    defparam i16_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4724));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1555 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_4725));
    defparam i18_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1556 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4726));
    defparam i15_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1557 (.I0(n41_adj_4723), .I1(n33_adj_4722), .I2(n2889), 
            .I3(n2901), .O(n46_adj_4727));
    defparam i21_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1558 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4728));
    defparam i14_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1559 (.I0(n43_adj_4725), .I1(n2904), .I2(n38_adj_4724), 
            .I3(n2893), .O(n47_adj_4729));
    defparam i22_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4729), .I1(n39_adj_4728), .I2(n46_adj_4727), 
            .I3(n40_adj_4726), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_25 (.CI(n25539), .I0(bit_ctr[23]), .I1(GND_net), .CO(n25540));
    SB_CARRY sub_14_add_2_20 (.CI(n25788), .I0(timer[18]), .I1(n1[18]), 
            .CO(n25789));
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_470[13]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n25787), .O(n23_adj_4730)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n25787), .I0(timer[17]), .I1(n1[17]), 
            .CO(n25788));
    SB_LUT4 i29268_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35440));
    defparam i29268_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n25786), .O(one_wire_N_470[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n25786), .I0(timer[16]), .I1(n1[16]), 
            .CO(n25787));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n25785), .O(one_wire_N_470[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_17 (.CI(n25785), .I0(timer[15]), .I1(n1[15]), 
            .CO(n25786));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n25784), .O(one_wire_N_470[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n25784), .I0(timer[14]), .I1(n1[14]), 
            .CO(n25785));
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n25783), .O(one_wire_N_470[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_15 (.CI(n25783), .I0(timer[13]), .I1(n1[13]), 
            .CO(n25784));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n25782), .O(one_wire_N_470[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_14 (.CI(n25782), .I0(timer[12]), .I1(n1[12]), 
            .CO(n25783));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n25781), .O(one_wire_N_470[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_13 (.CI(n25781), .I0(timer[11]), .I1(n1[11]), 
            .CO(n25782));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n25780), .O(one_wire_N_470[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n25780), .I0(timer[10]), .I1(n1[10]), 
            .CO(n25781));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n25779), .O(one_wire_N_470[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_11 (.CI(n25779), .I0(timer[9]), .I1(n1[9]), 
            .CO(n25780));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n25538), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n25778), .O(one_wire_N_470[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n25538), .I0(bit_ctr[22]), .I1(GND_net), .CO(n25539));
    SB_CARRY sub_14_add_2_10 (.CI(n25778), .I0(timer[8]), .I1(n1[8]), 
            .CO(n25779));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n25537), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n25523), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n25777), .O(one_wire_N_470[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n25777), .I0(timer[7]), .I1(n1[7]), .CO(n25778));
    SB_CARRY add_21_23 (.CI(n25537), .I0(bit_ctr[21]), .I1(GND_net), .CO(n25538));
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_470[9]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n25776), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_8 (.CI(n25776), .I0(timer[6]), .I1(n1[6]), .CO(n25777));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n25775), .O(one_wire_N_470[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n25523), .I0(bit_ctr[7]), .I1(GND_net), .CO(n25524));
    SB_CARRY sub_14_add_2_7 (.CI(n25775), .I0(timer[5]), .I1(n1[5]), .CO(n25776));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n25774), .O(one_wire_N_470[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n35597));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n35597_bdd_4_lut (.I0(n35597), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n33265));
    defparam n35597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29397 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n35591));
    defparam bit_ctr_0__bdd_4_lut_29397.LUT_INIT = 16'he4aa;
    SB_LUT4 n35591_bdd_4_lut (.I0(n35591), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n33268));
    defparam n35591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_2_lut_adj_1560 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4731));
    defparam i3_2_lut_adj_1560.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1561 (.I0(bit_ctr[12]), .I1(n22_adj_4731), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4732));
    defparam i11_4_lut_adj_1561.LUT_INIT = 16'hfefc;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29392 (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n35585));
    defparam bit_ctr_0__bdd_4_lut_29392.LUT_INIT = 16'he4aa;
    SB_LUT4 n35585_bdd_4_lut (.I0(n35585), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n33271));
    defparam n35585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_1562 (.I0(n2294), .I1(n30_adj_4732), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4733));
    defparam i15_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n25517), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n25774), .I0(timer[4]), .I1(n1[4]), .CO(n25775));
    SB_LUT4 i13_4_lut_adj_1563 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4734));
    defparam i13_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1564 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4735));
    defparam i14_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n25773), .O(one_wire_N_470[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1565 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4736));
    defparam i12_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1566 (.I0(n31_adj_4736), .I1(n33_adj_4735), .I2(n32_adj_4734), 
            .I3(n34_adj_4733), .O(n2324));
    defparam i18_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_5 (.CI(n25773), .I0(timer[3]), .I1(n1[3]), .CO(n25774));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n25772), .O(one_wire_N_470[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n25772), .I0(timer[2]), .I1(n1[2]), .CO(n25773));
    SB_LUT4 i19_4_lut_adj_1567 (.I0(bit_ctr[23]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46_adj_4737));
    defparam i19_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1568 (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[25]), 
            .I3(bit_ctr[10]), .O(n44_adj_4738));
    defparam i17_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29387 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n35537));
    defparam bit_ctr_0__bdd_4_lut_29387.LUT_INIT = 16'he4aa;
    SB_LUT4 n35537_bdd_4_lut (.I0(n35537), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n35540));
    defparam n35537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i18_4_lut_adj_1569 (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45_adj_4739));
    defparam i18_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29348 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n35531));
    defparam bit_ctr_0__bdd_4_lut_29348.LUT_INIT = 16'he4aa;
    SB_LUT4 n35531_bdd_4_lut (.I0(n35531), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n35534));
    defparam n35531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16_4_lut_adj_1570 (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43_adj_4740));
    defparam i16_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n25522), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29267_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35439));
    defparam i29267_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_8 (.CI(n25522), .I0(bit_ctr[6]), .I1(GND_net), .CO(n25523));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n25536), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4741), .I1(timer[1]), .I2(n1[1]), 
            .I3(n25771), .O(n27418)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_22 (.CI(n25536), .I0(bit_ctr[20]), .I1(GND_net), .CO(n25537));
    SB_LUT4 i15_4_lut_adj_1571 (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42_adj_4742));
    defparam i15_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_29343 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n35519));
    defparam bit_ctr_0__bdd_4_lut_29343.LUT_INIT = 16'he4aa;
    SB_LUT4 i13_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(GND_net), .O(n40_adj_4743));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 n35519_bdd_4_lut (.I0(n35519), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n34700));
    defparam n35519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i21_4_lut_adj_1572 (.I0(bit_ctr[26]), .I1(n42_adj_4742), .I2(bit_ctr[13]), 
            .I3(bit_ctr[22]), .O(n48_adj_4744));
    defparam i21_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_3 (.CI(n25771), .I0(timer[1]), .I1(n1[1]), .CO(n25772));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_470[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4741)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n25771));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n22673), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n27721));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n22673), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n25535), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n25967), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n25966), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25_4_lut_adj_1573 (.I0(n43_adj_4740), .I1(n45_adj_4739), .I2(n44_adj_4738), 
            .I3(n46_adj_4737), .O(n52));
    defparam i25_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_937_10 (.CI(n25966), .I0(n1302), .I1(n1334), .CO(n25967));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n25965), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_21 (.CI(n25535), .I0(bit_ctr[19]), .I1(GND_net), .CO(n25536));
    SB_CARRY add_21_3 (.CI(n25517), .I0(bit_ctr[1]), .I1(GND_net), .CO(n25518));
    SB_CARRY mod_5_add_937_9 (.CI(n25965), .I0(n1303), .I1(n1334), .CO(n25966));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n25534), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n25964), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n25521), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5016_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n31167), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i5016_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_CARRY add_21_20 (.CI(n25534), .I0(bit_ctr[18]), .I1(GND_net), .CO(n25535));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n25533), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_8 (.CI(n25964), .I0(n1304), .I1(n1334), .CO(n25965));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n25963), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n25963), .I0(n1305), .I1(n1334), .CO(n25964));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n25962), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n25962), .I0(n1306), .I1(n1334), .CO(n25963));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n25961), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n25961), .I0(n1307), .I1(n1334), .CO(n25962));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n25960), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_19 (.CI(n25533), .I0(bit_ctr[17]), .I1(GND_net), .CO(n25534));
    SB_CARRY mod_5_add_937_4 (.CI(n25960), .I0(n1308), .I1(n1334), .CO(n25961));
    SB_LUT4 i27922_3_lut_4_lut (.I0(n27197), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n16468), .O(n34034));
    defparam i27922_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n35430), 
            .I3(n25959), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n25959), .I0(n1309), .I1(n35430), .CO(n25960));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n35430), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n35430), 
            .CO(n25959));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n25517));
    SB_LUT4 i28214_3_lut_4_lut (.I0(n16468), .I1(n34387), .I2(start), 
            .I3(\state[1] ), .O(n34388));
    defparam i28214_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n22763), .I1(\state[1] ), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n33056));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n25532), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_319[1] ), .O(n17985));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n26604), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n26603), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n26603), .I0(n1599), .I1(n1631), .CO(n26604));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n26602), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n26602), .I0(n1600), .I1(n1631), .CO(n26603));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n26601), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n26601), .I0(n1601), .I1(n1631), .CO(n26602));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n26600), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut_adj_1574 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4745));
    defparam i10_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_10 (.CI(n26600), .I0(n1602), .I1(n1631), .CO(n26601));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n26599), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n26599), .I0(n1603), .I1(n1631), .CO(n26600));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n26598), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n26598), .I0(n1604), .I1(n1631), .CO(n26599));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n26597), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1575 (.I0(n2203), .I1(n28_adj_4745), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4746));
    defparam i14_4_lut_adj_1575.LUT_INIT = 16'hfeee;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n17772), 
            .D(n255[31]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i12_4_lut_adj_1576 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4747));
    defparam i12_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_7 (.CI(n26597), .I0(n1605), .I1(n1631), .CO(n26598));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n26596), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1577 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4748));
    defparam i13_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1578 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4749));
    defparam i11_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1138_6 (.CI(n26596), .I0(n1606), .I1(n1631), .CO(n26597));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n26595), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n26595), .I0(n1607), .I1(n1631), .CO(n26596));
    SB_LUT4 i17_4_lut_adj_1579 (.I0(n29_adj_4749), .I1(n31_adj_4748), .I2(n30_adj_4747), 
            .I3(n32_adj_4746), .O(n2225));
    defparam i17_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n26594), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n26594), .I0(n1608), .I1(n1631), .CO(n26595));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n35431), 
            .I3(n26593), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n26593), .I0(n1609), .I1(n35431), .CO(n26594));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n35431), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n35431), 
            .CO(n26593));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n26592), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n26591), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n26591), .I0(n1698), .I1(n1730), .CO(n26592));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n26590), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n26590), .I0(n1699), .I1(n1730), .CO(n26591));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n26589), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n26589), .I0(n1700), .I1(n1730), .CO(n26590));
    SB_CARRY add_21_18 (.CI(n25532), .I0(bit_ctr[16]), .I1(GND_net), .CO(n25533));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n26588), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n26588), .I0(n1701), .I1(n1730), .CO(n26589));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n26587), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n26587), .I0(n1702), .I1(n1730), .CO(n26588));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n26586), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n26586), .I0(n1703), .I1(n1730), .CO(n26587));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n26585), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n26585), .I0(n1704), .I1(n1730), .CO(n26586));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n26584), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n26584), .I0(n1705), .I1(n1730), .CO(n26585));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n26583), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n26583), .I0(n1706), .I1(n1730), .CO(n26584));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n26582), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n26582), .I0(n1707), .I1(n1730), .CO(n26583));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n26581), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n26581), .I0(n1708), .I1(n1730), .CO(n26582));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n35432), 
            .I3(n26580), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n26580), .I0(n1709), .I1(n35432), .CO(n26581));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n35432), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n35432), 
            .CO(n26580));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n26579), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n26578), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n26578), .I0(n1797), .I1(n1829), .CO(n26579));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n26577), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n25531), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_14 (.CI(n26577), .I0(n1798), .I1(n1829), .CO(n26578));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n26576), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n26576), .I0(n1799), .I1(n1829), .CO(n26577));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n26575), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n26575), .I0(n1800), .I1(n1829), .CO(n26576));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n26574), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_7 (.CI(n25521), .I0(bit_ctr[5]), .I1(GND_net), .CO(n25522));
    SB_CARRY mod_5_add_1272_11 (.CI(n26574), .I0(n1801), .I1(n1829), .CO(n26575));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n26573), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n26573), .I0(n1802), .I1(n1829), .CO(n26574));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n26572), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n26572), .I0(n1803), .I1(n1829), .CO(n26573));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n26571), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n26571), .I0(n1804), .I1(n1829), .CO(n26572));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n26570), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n26570), .I0(n1805), .I1(n1829), .CO(n26571));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n26569), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n26569), .I0(n1806), .I1(n1829), .CO(n26570));
    SB_LUT4 i29265_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35437));
    defparam i29265_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24_4_lut_adj_1580 (.I0(bit_ctr[30]), .I1(n48_adj_4744), .I2(n40_adj_4743), 
            .I3(bit_ctr[24]), .O(n51_adj_4750));
    defparam i24_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(bit_ctr[3]), .I1(n51_adj_4750), .I2(bit_ctr[4]), 
            .I3(n52), .O(\state_3__N_319[1] ));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'hffec;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n18064));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n17772), 
            .D(n255[30]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n26568), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n26568), .I0(n1807), .I1(n1829), .CO(n26569));
    SB_LUT4 i1_2_lut_adj_1582 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n16534));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'hbbbb;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n26567), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n26567), .I0(n1808), .I1(n1829), .CO(n26568));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n35433), 
            .I3(n26566), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n26566), .I0(n1809), .I1(n35433), .CO(n26567));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n35433), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n35433), 
            .CO(n26566));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n26565), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n26564), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n26564), .I0(n1896), .I1(n1928), .CO(n26565));
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n18060));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1461__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n26563), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n26563), .I0(n1897), .I1(n1928), .CO(n26564));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n26562), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n26562), .I0(n1898), .I1(n1928), .CO(n26563));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n26561), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n26561), .I0(n1899), .I1(n1928), .CO(n26562));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n26560), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n26560), .I0(n1900), .I1(n1928), .CO(n26561));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n26559), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_17 (.CI(n25531), .I0(bit_ctr[15]), .I1(GND_net), .CO(n25532));
    SB_CARRY mod_5_add_1339_11 (.CI(n26559), .I0(n1901), .I1(n1928), .CO(n26560));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n25520), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n26558), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n26558), .I0(n1902), .I1(n1928), .CO(n26559));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n26557), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n26557), .I0(n1903), .I1(n1928), .CO(n26558));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n26556), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n25530), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n26556), .I0(n1904), .I1(n1928), .CO(n26557));
    SB_CARRY add_21_16 (.CI(n25530), .I0(bit_ctr[14]), .I1(GND_net), .CO(n25531));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n25529), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n25529), .I0(bit_ctr[13]), .I1(GND_net), .CO(n25530));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n25528), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n26555), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n26555), .I0(n1905), .I1(n1928), .CO(n26556));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n26554), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n26554), .I0(n1906), .I1(n1928), .CO(n26555));
    SB_CARRY add_21_14 (.CI(n25528), .I0(bit_ctr[12]), .I1(GND_net), .CO(n25529));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n26553), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n26553), .I0(n1907), .I1(n1928), .CO(n26554));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n26552), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n26552), .I0(n1908), .I1(n1928), .CO(n26553));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n35434), 
            .I3(n26551), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n26551), .I0(n1909), .I1(n35434), .CO(n26552));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n35434), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n35434), 
            .CO(n26551));
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n18575));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n18574));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i29257_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35429));
    defparam i29257_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n18573));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n18572));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n18571));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n18570));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n18569));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n18568));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n18567));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n18566));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n18565));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n18564));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n18563));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n18562));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n18561));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n18560));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n18559));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n18558));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n18557));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n18556));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n18555));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n18554));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n18553));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n18552));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n18551));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n18550));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n18549));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n18548));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n18547));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n18546));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n18545));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n26550), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk32MHz), .E(n17813), .D(state_3__N_319[0]), 
            .S(n31208));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n26549), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n26549), .I0(n1995), .I1(n2027), .CO(n26550));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n26548), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n26548), .I0(n1996), .I1(n2027), .CO(n26549));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n26547), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17524_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n22097));
    defparam i17524_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1107), .I1(n1104), .I2(n22097), .I3(n1108), 
            .O(n12_adj_4751));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1583 (.I0(n1105), .I1(n12_adj_4751), .I2(n1103), 
            .I3(n1106), .O(n1136));
    defparam i6_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29256_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35428));
    defparam i29256_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_15 (.CI(n26547), .I0(n1997), .I1(n2027), .CO(n26548));
    SB_LUT4 i16_4_lut_adj_1584 (.I0(n2786), .I1(n2798), .I2(n2794), .I3(n2795), 
            .O(n40_adj_4752));
    defparam i16_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1585 (.I0(n2796), .I1(n2799), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4753));
    defparam i14_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1586 (.I0(n2803), .I1(n2805), .I2(n2787), .I3(n2793), 
            .O(n39_adj_4754));
    defparam i15_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1587 (.I0(n2804), .I1(n2802), .I2(n2790), .I3(n2800), 
            .O(n37_adj_4755));
    defparam i13_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2807), .I1(n2801), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4756));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1588 (.I0(n2789), .I1(n2792), .I2(n2797), .I3(n2806), 
            .O(n42_adj_4757));
    defparam i18_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1589 (.I0(n37_adj_4755), .I1(n39_adj_4754), .I2(n38_adj_4753), 
            .I3(n40_adj_4752), .O(n46_adj_4758));
    defparam i22_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2791), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4759));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1590 (.I0(n33_adj_4759), .I1(n46_adj_4758), .I2(n42_adj_4757), 
            .I3(n34_adj_4756), .O(n2819));
    defparam i23_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i241_2_lut (.I0(LED_c), .I1(\state_3__N_319[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1039));   // verilog/neopixel.v(40[18] 45[12])
    defparam i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n25881), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n25880), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n25880), .I0(n1401), .I1(n1433), .CO(n25881));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n25879), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n25879), .I0(n1402), .I1(n1433), .CO(n25880));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n25878), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n25878), .I0(n1403), .I1(n1433), .CO(n25879));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n25877), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n25877), .I0(n1404), .I1(n1433), .CO(n25878));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n25876), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n25876), .I0(n1405), .I1(n1433), .CO(n25877));
    SB_LUT4 i2_2_lut_adj_1591 (.I0(n16468), .I1(n31237), .I2(GND_net), 
            .I3(GND_net), .O(n22737));
    defparam i2_2_lut_adj_1591.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n26546), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n25875), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n25875), .I0(n1406), .I1(n1433), .CO(n25876));
    SB_CARRY mod_5_add_1406_14 (.CI(n26546), .I0(n1998), .I1(n2027), .CO(n26547));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n26545), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n26545), .I0(n1999), .I1(n2027), .CO(n26546));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n26544), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n26544), .I0(n2000), .I1(n2027), .CO(n26545));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n26543), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n26543), .I0(n2001), .I1(n2027), .CO(n26544));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n25874), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n25874), .I0(n1407), .I1(n1433), .CO(n25875));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n26542), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n26542), .I0(n2002), .I1(n2027), .CO(n26543));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n25873), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n26541), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n26541), .I0(n2003), .I1(n2027), .CO(n26542));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n26540), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n26540), .I0(n2004), .I1(n2027), .CO(n26541));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n26539), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n26539), .I0(n2005), .I1(n2027), .CO(n26540));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n26538), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n26538), .I0(n2006), .I1(n2027), .CO(n26539));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n26537), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n26537), .I0(n2007), .I1(n2027), .CO(n26538));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n26536), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n26536), .I0(n2008), .I1(n2027), .CO(n26537));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n35435), 
            .I3(n26535), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_3 (.CI(n26535), .I0(n2009), .I1(n35435), .CO(n26536));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n35435), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n35435), 
            .CO(n26535));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n26534), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n26533), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n26533), .I0(n2094), .I1(n2126), .CO(n26534));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n26532), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n25873), .I0(n1408), .I1(n1433), .CO(n25874));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n35436), 
            .I3(n25872), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n25872), .I0(n1409), .I1(n35436), .CO(n25873));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n35436), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i29266_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35438));
    defparam i29266_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n35436), 
            .CO(n25872));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n25871), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n25870), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n25870), .I0(n1500), .I1(n1532), .CO(n25871));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n25869), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n25869), .I0(n1501), .I1(n1532), .CO(n25870));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n25868), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n25868), .I0(n1502), .I1(n1532), .CO(n25869));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n25867), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n26532), .I0(n2095), .I1(n2126), .CO(n26533));
    SB_CARRY mod_5_add_1071_9 (.CI(n25867), .I0(n1503), .I1(n1532), .CO(n25868));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n31384), .D(\neo_pixel_transmitter.done_N_533 ), 
            .R(n33056));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n25866), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n26531), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n25866), .I0(n1504), .I1(n1532), .CO(n25867));
    SB_CARRY mod_5_add_1473_16 (.CI(n26531), .I0(n2096), .I1(n2126), .CO(n26532));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n26530), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n17772), 
            .D(n255[29]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_15 (.CI(n26530), .I0(n2097), .I1(n2126), .CO(n26531));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n25865), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n26529), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n25865), .I0(n1505), .I1(n1532), .CO(n25866));
    SB_CARRY mod_5_add_1473_14 (.CI(n26529), .I0(n2098), .I1(n2126), .CO(n26530));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n25864), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n25864), .I0(n1506), .I1(n1532), .CO(n25865));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n26528), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n25863), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n25863), .I0(n1507), .I1(n1532), .CO(n25864));
    SB_CARRY mod_5_add_1473_13 (.CI(n26528), .I0(n2099), .I1(n2126), .CO(n26529));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n25862), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n25862), .I0(n1508), .I1(n1532), .CO(n25863));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n35438), 
            .I3(n25861), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n26527), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n25520), .I0(bit_ctr[4]), .I1(GND_net), .CO(n25521));
    SB_LUT4 i3226_4_lut (.I0(n22737), .I1(n1039), .I2(\state[1] ), .I3(n16534), 
            .O(n4820));
    defparam i3226_4_lut.LUT_INIT = 16'h3f35;
    SB_CARRY mod_5_add_1473_12 (.CI(n26527), .I0(n2100), .I1(n2126), .CO(n26528));
    SB_CARRY mod_5_add_1071_3 (.CI(n25861), .I0(n1509), .I1(n35438), .CO(n25862));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n35438), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n35438), 
            .CO(n25861));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n25860), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n26526), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n26526), .I0(n2101), .I1(n2126), .CO(n26527));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n26525), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n26525), .I0(n2102), .I1(n2126), .CO(n26526));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n26524), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n26524), .I0(n2103), .I1(n2126), .CO(n26525));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n26523), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n26523), .I0(n2104), .I1(n2126), .CO(n26524));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n26522), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1461__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1461__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1473_7 (.CI(n26522), .I0(n2105), .I1(n2126), .CO(n26523));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n26521), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n26521), .I0(n2106), .I1(n2126), .CO(n26522));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n26520), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n26520), .I0(n2107), .I1(n2126), .CO(n26521));
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n25859), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n26519), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_6 (.CI(n25859), .I0(n906), .I1(VCC_net), .CO(n25860));
    SB_CARRY mod_5_add_1473_4 (.CI(n26519), .I0(n2108), .I1(n2126), .CO(n26520));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n35437), 
            .I3(n26518), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n26518), .I0(n2109), .I1(n35437), .CO(n26519));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n35437), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n35437), 
            .CO(n26518));
    SB_LUT4 i28415_4_lut (.I0(n27197), .I1(n31237), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n34387));
    defparam i28415_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n26517), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28208_2_lut (.I0(n31237), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n34056));
    defparam i28208_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n26516), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n26516), .I0(n2193), .I1(n2225), .CO(n26517));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n26515), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i53_4_lut (.I0(n34056), .I1(n22763), .I2(\state[1] ), .I3(n16468), 
            .O(n31350));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_CARRY mod_5_add_1540_18 (.CI(n26515), .I0(n2194), .I1(n2225), .CO(n26516));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n26514), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n26514), .I0(n2195), .I1(n2225), .CO(n26515));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n26513), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n26513), .I0(n2196), .I1(n2225), .CO(n26514));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n26512), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n26512), .I0(n2197), .I1(n2225), .CO(n26513));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n26511), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n31210), .I2(VCC_net), 
            .I3(n25858), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_14 (.CI(n26511), .I0(n2198), .I1(n2225), .CO(n26512));
    SB_CARRY mod_5_add_669_5 (.CI(n25858), .I0(n31210), .I1(VCC_net), 
            .CO(n25859));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n26510), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n26510), .I0(n2199), .I1(n2225), .CO(n26511));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n26509), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i52_4_lut (.I0(n31350), .I1(n34388), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n31384));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_533 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_12 (.CI(n26509), .I0(n2200), .I1(n2225), .CO(n26510));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n26508), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n26508), .I0(n2201), .I1(n2225), .CO(n26509));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n26507), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n26507), .I0(n2202), .I1(n2225), .CO(n26508));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n26506), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n26506), .I0(n2203), .I1(n2225), .CO(n26507));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n26505), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n26505), .I0(n2204), .I1(n2225), .CO(n26506));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n26504), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n26504), .I0(n2205), .I1(n2225), .CO(n26505));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n26503), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n26503), .I0(n2206), .I1(n2225), .CO(n26504));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n26502), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n26502), .I0(n2207), .I1(n2225), .CO(n26503));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17881), .I2(VCC_net), 
            .I3(n25857), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n26501), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n26501), .I0(n2208), .I1(n2225), .CO(n26502));
    SB_CARRY mod_5_add_669_4 (.CI(n25857), .I0(n17881), .I1(VCC_net), 
            .CO(n25858));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n15162), .I2(GND_net), 
            .I3(n25856), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n35439), 
            .I3(n26500), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n26500), .I0(n2209), .I1(n35439), .CO(n26501));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n35439), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n35439), 
            .CO(n26500));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n26499), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n26498), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n26498), .I0(n2292), .I1(n2324), .CO(n26499));
    SB_LUT4 i7_4_lut_adj_1592 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4760));
    defparam i7_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n26497), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n26497), .I0(n2293), .I1(n2324), .CO(n26498));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n26496), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n26496), .I0(n2294), .I1(n2324), .CO(n26497));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n26495), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n26495), .I0(n2295), .I1(n2324), .CO(n26496));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n26494), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n26494), .I0(n2296), .I1(n2324), .CO(n26495));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n26493), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n26493), .I0(n2297), .I1(n2324), .CO(n26494));
    SB_CARRY mod_5_add_669_3 (.CI(n25856), .I0(n15162), .I1(GND_net), 
            .CO(n25857));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n26492), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n26492), .I0(n2298), .I1(n2324), .CO(n26493));
    SB_LUT4 i9_4_lut_adj_1593 (.I0(n1504), .I1(n18_adj_4760), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4761));
    defparam i9_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n26491), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n26491), .I0(n2299), .I1(n2324), .CO(n26492));
    SB_LUT4 i4_3_lut_adj_1594 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4762));
    defparam i4_3_lut_adj_1594.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n26490), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n26490), .I0(n2300), .I1(n2324), .CO(n26491));
    SB_LUT4 i10_4_lut_adj_1595 (.I0(n15_adj_4762), .I1(n20_adj_4761), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n26489), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n26489), .I0(n2301), .I1(n2324), .CO(n26490));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n26488), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i29264_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35436));
    defparam i29264_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1607_10 (.CI(n26488), .I0(n2302), .I1(n2324), .CO(n26489));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n26487), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n26487), .I0(n2303), .I1(n2324), .CO(n26488));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n26486), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n26486), .I0(n2304), .I1(n2324), .CO(n26487));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n26485), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n26485), .I0(n2305), .I1(n2324), .CO(n26486));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n26484), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n26484), .I0(n2306), .I1(n2324), .CO(n26485));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n26483), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n26483), .I0(n2307), .I1(n2324), .CO(n26484));
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n25856));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n26482), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n26482), .I0(n2308), .I1(n2324), .CO(n26483));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n35440), 
            .I3(n26481), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n26481), .I0(n2309), .I1(n35440), .CO(n26482));
    SB_LUT4 i1_2_lut_adj_1596 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4763));
    defparam i1_2_lut_adj_1596.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n35440), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n35440), 
            .CO(n26481));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n26480), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18202_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n22779));
    defparam i18202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n26479), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n26479), .I0(n2391), .I1(n2423), .CO(n26480));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n26478), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i28781_4_lut (.I0(\state[1] ), .I1(n34034), .I2(n4820), .I3(state[0]), 
            .O(n17772));
    defparam i28781_4_lut.LUT_INIT = 16'h0f11;
    SB_CARRY mod_5_add_1674_20 (.CI(n26478), .I0(n2392), .I1(n2423), .CO(n26479));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n26477), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n26477), .I0(n2393), .I1(n2423), .CO(n26478));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n26476), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n26476), .I0(n2394), .I1(n2423), .CO(n26477));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n26475), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n26475), .I0(n2395), .I1(n2423), .CO(n26476));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n26474), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n26474), .I0(n2396), .I1(n2423), .CO(n26475));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n26473), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n26473), .I0(n2397), .I1(n2423), .CO(n26474));
    SB_LUT4 i13_4_lut_adj_1597 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4763), 
            .O(n30_adj_4764));
    defparam i13_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n26472), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n26472), .I0(n2398), .I1(n2423), .CO(n26473));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n26471), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n26471), .I0(n2399), .I1(n2423), .CO(n26472));
    SB_LUT4 i11_4_lut_adj_1598 (.I0(n2098), .I1(n22779), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4765));
    defparam i11_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n26470), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n26470), .I0(n2400), .I1(n2423), .CO(n26471));
    SB_LUT4 i12_4_lut_adj_1599 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4766));
    defparam i12_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n26469), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n26469), .I0(n2401), .I1(n2423), .CO(n26470));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n26468), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n26468), .I0(n2402), .I1(n2423), .CO(n26469));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n26467), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n26467), .I0(n2403), .I1(n2423), .CO(n26468));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n26466), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n26466), .I0(n2404), .I1(n2423), .CO(n26467));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n26465), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n26465), .I0(n2405), .I1(n2423), .CO(n26466));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n26464), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n26464), .I0(n2406), .I1(n2423), .CO(n26465));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n26463), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n26463), .I0(n2407), .I1(n2423), .CO(n26464));
    SB_LUT4 i10_4_lut_adj_1600 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4767));
    defparam i10_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n26462), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n26462), .I0(n2408), .I1(n2423), .CO(n26463));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n35441), 
            .I3(n26461), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n26461), .I0(n2409), .I1(n35441), .CO(n26462));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n35441), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i16_4_lut_adj_1601 (.I0(n27_adj_4767), .I1(n29_adj_4766), .I2(n28_adj_4765), 
            .I3(n30_adj_4764), .O(n2126));
    defparam i16_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n35441), 
            .CO(n26461));
    SB_LUT4 i29263_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35435));
    defparam i29263_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n26436), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n26435), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n26435), .I0(n2490), .I1(n2522), .CO(n26436));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n26434), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n26434), .I0(n2491), .I1(n2522), .CO(n26435));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n26433), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n26433), .I0(n2492), .I1(n2522), .CO(n26434));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n26432), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n26432), .I0(n2493), .I1(n2522), .CO(n26433));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n26431), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n26431), .I0(n2494), .I1(n2522), .CO(n26432));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n26430), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n26430), .I0(n2495), .I1(n2522), .CO(n26431));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n26429), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n26429), .I0(n2496), .I1(n2522), .CO(n26430));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n26428), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n26428), .I0(n2497), .I1(n2522), .CO(n26429));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n26427), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n26427), .I0(n2498), .I1(n2522), .CO(n26428));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n26426), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n26426), .I0(n2499), .I1(n2522), .CO(n26427));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n26425), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n26425), .I0(n2500), .I1(n2522), .CO(n26426));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n26424), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n26424), .I0(n2501), .I1(n2522), .CO(n26425));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n26423), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n26423), .I0(n2502), .I1(n2522), .CO(n26424));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n26422), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n26422), .I0(n2503), .I1(n2522), .CO(n26423));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n26421), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n26421), .I0(n2504), .I1(n2522), .CO(n26422));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n26420), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n26420), .I0(n2505), .I1(n2522), .CO(n26421));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n26419), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n26419), .I0(n2506), .I1(n2522), .CO(n26420));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n26418), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n26418), .I0(n2507), .I1(n2522), .CO(n26419));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n26417), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n26417), .I0(n2508), .I1(n2522), .CO(n26418));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n35442), 
            .I3(n26416), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n26416), .I0(n2509), .I1(n35442), .CO(n26417));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n35442), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n35442), 
            .CO(n26416));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n26415), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n26414), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n26414), .I0(n2589), .I1(n2621), .CO(n26415));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n26413), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n26413), .I0(n2590), .I1(n2621), .CO(n26414));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n26412), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n26412), .I0(n2591), .I1(n2621), .CO(n26413));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n26411), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n26411), .I0(n2592), .I1(n2621), .CO(n26412));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n26410), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n26410), .I0(n2593), .I1(n2621), .CO(n26411));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n26409), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n26409), .I0(n2594), .I1(n2621), .CO(n26410));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n26408), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n26408), .I0(n2595), .I1(n2621), .CO(n26409));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n26407), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n26407), .I0(n2596), .I1(n2621), .CO(n26408));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n26406), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n26406), .I0(n2597), .I1(n2621), .CO(n26407));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n26405), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n26405), .I0(n2598), .I1(n2621), .CO(n26406));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n26404), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n26404), .I0(n2599), .I1(n2621), .CO(n26405));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n26403), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n26403), .I0(n2600), .I1(n2621), .CO(n26404));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n26402), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n26402), .I0(n2601), .I1(n2621), .CO(n26403));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n26401), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n26401), .I0(n2602), .I1(n2621), .CO(n26402));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n26400), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n26400), .I0(n2603), .I1(n2621), .CO(n26401));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n26399), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n26399), .I0(n2604), .I1(n2621), .CO(n26400));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n26398), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n26398), .I0(n2605), .I1(n2621), .CO(n26399));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n26397), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n26397), .I0(n2606), .I1(n2621), .CO(n26398));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n26396), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n26396), .I0(n2607), .I1(n2621), .CO(n26397));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n26395), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n26395), .I0(n2608), .I1(n2621), .CO(n26396));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n35443), 
            .I3(n26394), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n26394), .I0(n2609), .I1(n35443), .CO(n26395));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n35443), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n35443), 
            .CO(n26394));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n26393), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n26392), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n26392), .I0(n1203), .I1(n1235), .CO(n26393));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n26391), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n26391), .I0(n1204), .I1(n1235), .CO(n26392));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n26390), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n26390), .I0(n1205), .I1(n1235), .CO(n26391));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n26389), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n26389), .I0(n1206), .I1(n1235), .CO(n26390));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n26388), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n26388), .I0(n1207), .I1(n1235), .CO(n26389));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n26387), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n26387), .I0(n1208), .I1(n1235), .CO(n26388));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n35444), 
            .I3(n26386), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n26386), .I0(n1209), .I1(n35444), .CO(n26387));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n35444), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n35444), 
            .CO(n26386));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n26385), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n26384), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n26384), .I0(n2688), .I1(n2720), .CO(n26385));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n26383), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n26383), .I0(n2689), .I1(n2720), .CO(n26384));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n26382), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n26382), .I0(n2690), .I1(n2720), .CO(n26383));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n26381), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n26381), .I0(n2691), .I1(n2720), .CO(n26382));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n26380), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n26380), .I0(n2692), .I1(n2720), .CO(n26381));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n26379), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n26379), .I0(n2693), .I1(n2720), .CO(n26380));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n26378), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n26378), .I0(n2694), .I1(n2720), .CO(n26379));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n26377), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n26377), .I0(n2695), .I1(n2720), .CO(n26378));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n26376), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n26376), .I0(n2696), .I1(n2720), .CO(n26377));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n26375), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n26375), .I0(n2697), .I1(n2720), .CO(n26376));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n26374), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n26374), .I0(n2698), .I1(n2720), .CO(n26375));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n26373), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n26373), .I0(n2699), .I1(n2720), .CO(n26374));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n26372), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n26372), .I0(n2700), .I1(n2720), .CO(n26373));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n26371), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n26371), .I0(n2701), .I1(n2720), .CO(n26372));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n26370), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n26370), .I0(n2702), .I1(n2720), .CO(n26371));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n26369), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n26369), .I0(n2703), .I1(n2720), .CO(n26370));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n26368), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n26368), .I0(n2704), .I1(n2720), .CO(n26369));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n26367), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n17772), 
            .D(n255[28]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1875_7 (.CI(n26367), .I0(n2705), .I1(n2720), .CO(n26368));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n26366), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n26366), .I0(n2706), .I1(n2720), .CO(n26367));
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n17772), 
            .D(n255[26]), .R(n17985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n26365), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n26365), .I0(n2707), .I1(n2720), .CO(n26366));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n26364), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n26364), .I0(n2708), .I1(n2720), .CO(n26365));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n35445), 
            .I3(n26363), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n26363), .I0(n2709), .I1(n35445), .CO(n26364));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n35445), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n35445), 
            .CO(n26363));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n26362), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n26361), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n26361), .I0(n2787), .I1(n2819), .CO(n26362));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n26360), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n26360), .I0(n2788), .I1(n2819), .CO(n26361));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n26359), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n26359), .I0(n2789), .I1(n2819), .CO(n26360));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n26358), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n26358), .I0(n2790), .I1(n2819), .CO(n26359));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n26357), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n26357), .I0(n2791), .I1(n2819), .CO(n26358));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n26356), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n26356), .I0(n2792), .I1(n2819), .CO(n26357));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n26355), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i18238_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n22815));
    defparam i18238_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1602 (.I0(n1403), .I1(n22815), .I2(n1404), .I3(n1405), 
            .O(n16_adj_4768));
    defparam i6_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1603 (.I0(n1402), .I1(n1400), .I2(n1401), .I3(n1406), 
            .O(n17_adj_4769));
    defparam i7_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1604 (.I0(n17_adj_4769), .I1(n1408), .I2(n16_adj_4768), 
            .I3(n1407), .O(n1433));
    defparam i9_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i29255_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35427));
    defparam i29255_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(n31372), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n14233));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i25055_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n22673), .I2(n608), 
            .I3(bit_ctr[29]), .O(n31212));
    defparam i25055_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 i18099_2_lut_3_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n22673));
    defparam i18099_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i28067_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17881));
    defparam i28067_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_LUT4 i3_4_lut_4_lut_adj_1605 (.I0(n807), .I1(n15144), .I2(n31167), 
            .I3(bit_ctr[27]), .O(n838));
    defparam i3_4_lut_4_lut_adj_1605.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n15144), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n31167), .O(n31210));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n33265), .I2(n33268), 
            .I3(n27729), .O(n35447));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i18186_4_lut (.I0(one_wire_N_470[9]), .I1(n16589), .I2(one_wire_N_470[11]), 
            .I3(one_wire_N_470[10]), .O(n22763));
    defparam i18186_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i25079_3_lut (.I0(one_wire_N_470[4]), .I1(n27418), .I2(one_wire_N_470[3]), 
            .I3(GND_net), .O(n31237));
    defparam i25079_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 n35447_bdd_4_lut (.I0(n35447), .I1(n34700), .I2(n33271), .I3(n27729), 
            .O(n35450));
    defparam n35447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1606 (.I0(one_wire_N_470[3]), .I1(one_wire_N_470[4]), 
            .I2(one_wire_N_470[2]), .I3(GND_net), .O(n27197));
    defparam i2_3_lut_adj_1606.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1607 (.I0(one_wire_N_470[5]), .I1(one_wire_N_470[11]), 
            .I2(one_wire_N_470[7]), .I3(n16589), .O(n14_adj_4770));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1608 (.I0(n9), .I1(n14_adj_4770), .I2(one_wire_N_470[10]), 
            .I3(one_wire_N_470[8]), .O(n16468));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i25206_4_lut (.I0(n16468), .I1(n27197), .I2(n31237), .I3(state[0]), 
            .O(n31372));
    defparam i25206_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i28220_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n33986));
    defparam i28220_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i25144_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n31372), .I3(GND_net), .O(n31304));
    defparam i25144_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1609 (.I0(n31304), .I1(n33986), .I2(\state[1] ), 
            .I3(n22763), .O(n7));
    defparam i15_4_lut_adj_1609.LUT_INIT = 16'h3a0a;
    SB_LUT4 i6_4_lut_adj_1610 (.I0(n11), .I1(n35), .I2(n33_adj_4682), 
            .I3(n29_adj_4685), .O(n14_adj_4771));
    defparam i6_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1611 (.I0(n49_adj_4666), .I1(n61), .I2(n15), 
            .I3(n51), .O(n13_adj_4772));
    defparam i5_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1612 (.I0(n41_adj_4671), .I1(n59), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4773));
    defparam i2_2_lut_adj_1612.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1613 (.I0(n31_adj_4684), .I1(n13_adj_4772), .I2(n14_adj_4771), 
            .I3(GND_net), .O(n19_adj_4774));
    defparam i1_3_lut_adj_1613.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_1614 (.I0(n21_adj_4693), .I1(n13_adj_4697), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4775));
    defparam i2_2_lut_adj_1614.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1615 (.I0(bit_ctr[3]), .I1(n6_adj_4775), .I2(n53), 
            .I3(n3209), .O(n32361));
    defparam i3_4_lut_adj_1615.LUT_INIT = 16'hfefc;
    SB_LUT4 i14_4_lut_adj_1616 (.I0(n39_adj_4673), .I1(n19_adj_4774), .I2(n19_adj_4695), 
            .I3(n20_adj_4773), .O(n32_adj_4776));
    defparam i14_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1617 (.I0(n63), .I1(n32361), .I2(n27_adj_4687), 
            .I3(n17_adj_4696), .O(n30_adj_4777));
    defparam i12_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1618 (.I0(n37_adj_4680), .I1(n55), .I2(n45_adj_4669), 
            .I3(n23_adj_4692), .O(n31_adj_4778));
    defparam i13_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1619 (.I0(n47_adj_4668), .I1(n43_adj_4670), .I2(n57), 
            .I3(n25_adj_4688), .O(n29_adj_4779));
    defparam i11_4_lut_adj_1619.LUT_INIT = 16'hfffe;
    SB_LUT4 i28895_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_518));   // verilog/neopixel.v(36[4] 116[11])
    defparam i28895_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i17_4_lut_adj_1620 (.I0(n29_adj_4779), .I1(n31_adj_4778), .I2(n30_adj_4777), 
            .I3(n32_adj_4776), .O(n27382));
    defparam i17_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1621 (.I0(n21_adj_4705), .I1(n23_adj_4730), .I2(n22_adj_4698), 
            .I3(n24_adj_4721), .O(n36_adj_4644));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i28306_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n27382), .I3(GND_net), 
            .O(color_bit_N_513[4]));
    defparam i28306_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i28221_4_lut (.I0(n35534), .I1(n27729), .I2(n35540), .I3(bit_ctr[2]), 
            .O(n34030));
    defparam i28221_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i17332_4_lut (.I0(n35450), .I1(\state_3__N_319[1] ), .I2(n34030), 
            .I3(color_bit_N_513[4]), .O(state_3__N_319[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i17332_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i2_2_lut_adj_1622 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4780));
    defparam i2_2_lut_adj_1622.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1623 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4781));
    defparam i12_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1624 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4782));
    defparam i10_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1625 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4783));
    defparam i11_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1626 (.I0(bit_ctr[15]), .I1(n18_adj_4780), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4784));
    defparam i9_4_lut_adj_1626.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1627 (.I0(n25_adj_4784), .I1(n27_adj_4783), .I2(n26_adj_4782), 
            .I3(n28_adj_4781), .O(n2027));
    defparam i15_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[2] , GND_net, \Kp[3] , \Kp[4] , IntegralLimit, 
            \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , \Kp[10] , 
            \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[1] , \Kp[0] , 
            PWMLimit, \Ki[0] , \Ki[14] , duty, clk32MHz, \Kp[15] , 
            VCC_net, \Ki[15] , \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , 
            \Ki[5] , \Ki[6] , \Ki[12] , setpoint, motor_state, \Ki[7] , 
            \Ki[8] , \Ki[9] , \Ki[10] , n35425, \Ki[11] , \Ki[13] ) /* synthesis syn_module_defined=1 */ ;
    input \Kp[2] ;
    input GND_net;
    input \Kp[3] ;
    input \Kp[4] ;
    input [23:0]IntegralLimit;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input [23:0]PWMLimit;
    input \Ki[0] ;
    input \Ki[14] ;
    output [23:0]duty;
    input clk32MHz;
    input \Kp[15] ;
    input VCC_net;
    input \Ki[15] ;
    input \Ki[1] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[12] ;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    output n35425;
    input \Ki[11] ;
    input \Ki[13] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n174, n247;
    wire [23:0]duty_23__N_3563;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n25615, n320;
    wire [23:0]n1_adj_4632;
    
    wire n393, n466, n27019;
    wire [12:0]n9454;
    
    wire n831, n27020;
    wire [13:0]n9438;
    
    wire n758, n27018, n539, n685, n27017, n612, n27016, n539_adj_4211, 
        n27015, n466_adj_4212, n27014, n393_adj_4213, n27013, n320_adj_4214, 
        n27012, n247_adj_4215, n27011, n612_adj_4216, n685_adj_4217, 
        n174_adj_4218, n27010, n32, n101;
    wire [14:0]n9421;
    
    wire n1120, n27009, n1047, n27008, n974, n27007, n901, n27006, 
        n828, n27005, n755, n27004, n682, n27003, n609, n27002, 
        n536, n27001, n463, n27000, n390, n26999, n317, n26998, 
        n244, n26997, n171, n26996, n29, n98;
    wire [15:0]n9403;
    
    wire n26995, n1117, n26994, n1044, n26993, n971, n26992, n898, 
        n26991, n825, n26990, n752, n26989, n679, n26988, n606, 
        n26987, n533, n26986, n460, n26985, n387, n26984, n314, 
        n26983, n241, n26982, n168, n26981, n26, n95;
    wire [16:0]n9384;
    
    wire n26980, n26979, n1114, n26978, n1041, n26977, n968, n26976, 
        n895, n26975, n822, n26974, n749, n26973, n676, n26972, 
        n603, n26971, n530, n26970, n457, n26969, n384, n26968, 
        n311, n26967, n238, n26966, n165, n26965, n23, n92;
    wire [17:0]n9364;
    
    wire n26964, n26963, n26962, n1111, n26961, n1038, n26960, 
        n965, n26959, n892, n26958, n819, n26957, n746, n26956, 
        n673, n26955, n600, n26954, n527, n26953, n454, n26952, 
        n381, n26951, n308, n26950, n235, n26949, n162, n26948, 
        n20, n89;
    wire [18:0]n9343;
    
    wire n26947, n26946, n26945, n26944, n1108, n26943, n1035, 
        n26942, n962, n26941, n889, n26940, n816, n26939, n743, 
        n26938, n670, n26937, n597, n26936, n524, n26935, n451, 
        n26934, n378, n26933, n305, n26932, n232, n26931, n159, 
        n26930, n17_adj_4219, n86;
    wire [19:0]n9321;
    
    wire n26929, n26928, n26927, n26926, n26925, n1105, n26924, 
        n1032, n26923, n959, n26922, n886, n26921, n813, n26920, 
        n740, n26919, n667, n26918, n594, n26917, n521, n26916, 
        n448, n26915, n375, n26914, n302, n26913, n229, n26912, 
        n156, n26911, n14_adj_4220, n83;
    wire [20:0]n9298;
    
    wire n26910, n26909, n26908, n26907, n26906, n26905, n1102, 
        n26904, n1029, n26903, n956, n26902, n883, n26901, n810, 
        n26900, n737, n26899, n664, n26898, n591, n26897, n518, 
        n26896, n445, n26895, n372, n26894, n299, n26893, n226, 
        n26892, n153, n26891, n11_adj_4221, n80;
    wire [0:0]n7409;
    wire [21:0]n9274;
    
    wire n26890;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3463 ;
    
    wire n26889, n26888, n26887, n26886, n26885, n26884, n26883, 
        n1096, n26882, n1023, n26881, n950, n26880, n877, n26879, 
        n804, n26878, n731, n26877, n658, n26876, n585, n26875, 
        n512, n26874, n439, n26873, n366, n26872, n293, n26871, 
        n220, n26870, n147, n26869, n5, n74, n26868, n26867, 
        n26866, n26865, n26864, n26863, n26862, n1099, n26861, 
        n1026, n26860, n953, n26859, n880, n26858, n807, n26857, 
        n734, n26856, n661, n26855, n588, n26854, n515, n26853, 
        n442, n26852, n369, n26851, n296, n26850, n223, n26849, 
        n150, n26848, n8, n77;
    wire [5:0]n9241;
    
    wire n32507, n490, n26847;
    wire [4:0]n9249;
    
    wire n417, n26846, n344, n26845, n271, n26844, n198_adj_4222, 
        n26843, n56, n125;
    wire [6:0]n9232;
    
    wire n560, n26842, n758_adj_4223, n831_adj_4224, n487, n26841, 
        n414, n26840, n904, n341, n26839, n977, n1050, n104, 
        n35, n177, \PID_CONTROLLER.integral_23__N_3511 ;
    wire [23:0]n3005;
    wire [23:0]n1_adj_4633;
    
    wire n250, n268, n26838, n195_adj_4231, n26837, n53, n122;
    wire [7:0]n9222;
    
    wire n630, n26836, n557, n26835, n484, n26834, n411, n26833, 
        n338, n26832, n34800, n29_adj_4232, n34801, n265, n26831, 
        n192_adj_4233, n26830, n50, n119;
    wire [8:0]n9211;
    
    wire n700, n26829, n627, n26828, n554, n26827, n481, n26826, 
        n408, n26825, n33, n31, n34207, n34201, n323, n30, n10_adj_4234, 
        n35_adj_4235, n34199, n34867, n694, n25616, n25750, n25751, 
        n335, n26824, n396, n469, n542, n615, n688, n761, n834, 
        n907, n980, n107, n38, n262, n26823, n180, n253, n767, 
        n326, n399, n840, n472, n545, n618, n691, n764, n837, 
        n910, n110, n41, n183_adj_4240, n256, n329, n402, n475, 
        n548, n189_adj_4241, n26822, n621, n113, n44, n47, n116;
    wire [23:0]n257;
    
    wire n256_adj_4245;
    wire [23:0]duty_23__N_3538;
    
    wire duty_23__N_3562;
    wire [23:0]duty_23__N_3439;
    wire [9:0]n9199;
    
    wire n770, n26821, n25749, n697, n26820, n34735, n624, n26819;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n25614, n551, n26818, n478, n26817, n405, n26816, n332, 
        n26815, n259_adj_4252, n26814, n186_adj_4253, n26813, n34914, 
        n77_adj_4254;
    wire [10:0]n9186;
    
    wire n26812, n26811, n37, n34915, n8_adj_4256, n150_adj_4257, 
        n223_adj_4258, n26810, n296_adj_4259, n369_adj_4260, n442_adj_4261, 
        n25748, n515_adj_4262, n588_adj_4263, n661_adj_4264, n26809, 
        n734_adj_4265, n807_adj_4266, n880_adj_4267, n953_adj_4268, 
        n1026_adj_4269, n1099_adj_4270, n26808, n39, n34898, n26807, 
        n74_adj_4271, n5_adj_4272, n147_adj_4273, n43, n41_adj_4274, 
        n34857, n34192, n34733, n34662, n45, n34190, n34816, n40, 
        n220_adj_4275, n293_adj_4276, n366_adj_4277, n34818, n26806, 
        n26805, n439_adj_4278, n26804, n26803, n512_adj_4279;
    wire [11:0]n9172;
    
    wire n26802, n26801, n585_adj_4281, n658_adj_4282, n731_adj_4284, 
        n804_adj_4285, n877_adj_4286, n950_adj_4287, n1023_adj_4289, 
        n1096_adj_4290, n26800, n26799, n80_adj_4291, n11_adj_4292, 
        n153_adj_4293, n26798, n41_adj_4294, n226_adj_4295, n26797, 
        n299_adj_4299, n26796;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3514 ;
    
    wire n25747, n372_adj_4300, n445_adj_4301, n518_adj_4302, n39_adj_4303, 
        n591_adj_4306, n664_adj_4307, n737_adj_4308, n810_adj_4309, 
        n883_adj_4310, n956_adj_4311, n1029_adj_4312, n1102_adj_4313, 
        n83_adj_4314, n14_adj_4315, n156_adj_4316, n229_adj_4317, n302_adj_4318, 
        n26795, n26794, n26793, n45_adj_4319, n25746, n26792, n43_adj_4320, 
        n25745, n375_adj_4321, n448_adj_4322, n521_adj_4323, n594_adj_4324, 
        n667_adj_4325, n740_adj_4326, n813_adj_4327, n886_adj_4328, 
        n959_adj_4329, n45_adj_4330;
    wire [12:0]n9157;
    
    wire n26791, n41_adj_4331, n25744, n26790, n43_adj_4332, n39_adj_4333, 
        n25743, n37_adj_4334, n29_adj_4335, n31_adj_4336, n23_adj_4337, 
        n25_adj_4338, n26789, n35_adj_4339, n9_adj_4340, n17_adj_4341, 
        n19_adj_4342, n21_adj_4343, n26788, n1032_adj_4344, n26787, 
        n26786, n26785, n26784, n37_adj_4345, n25742, n26783, n26782, 
        n35_adj_4346, n25741, n26781, n33_adj_4347, n25740, n31_adj_4348, 
        n25739, n26780;
    wire [13:0]n9141;
    
    wire n26779, n26778, n26777, n33_adj_4349, n26776, n26775, n26774, 
        n29_adj_4350, n25738, n27, n25737, n25_adj_4351, n25736, 
        n23_adj_4352, n25735, n26773, n26772, n21_adj_4353, n25734, 
        n26771, n26770, n19_adj_4354, n25733, n26769, n26768, n26767, 
        n32_adj_4355, n101_adj_4356;
    wire [14:0]n9124;
    
    wire n1120_adj_4357, n26766, n1047_adj_4358, n26765, n974_adj_4359, 
        n26764, n901_adj_4360, n26763, n828_adj_4361, n26762, n17_adj_4362, 
        n25732, n755_adj_4364, n26761, n682_adj_4365, n26760, n15_adj_4366, 
        n25731, n1105_adj_4368, n11_adj_4369, n13_adj_4370, n15_adj_4371, 
        n27_adj_4372, n34176, n34170, n12_adj_4373, n10_adj_4374, 
        n30_adj_4375, n86_adj_4376, n17_adj_4377, n34186, n34464, 
        n159_adj_4378, n232_adj_4379, n305_adj_4380, n378_adj_4381, 
        n609_adj_4382, n26759, n536_adj_4383, n26758, n451_adj_4384, 
        n34460, n34798, n34634, n34855, n16_adj_4385, n6_adj_4386, 
        n34780, n34781, n8_adj_4387, n524_adj_4388, n463_adj_4389, 
        n26757, n597_adj_4390, n670_adj_4391, n13_adj_4392, n25730, 
        n390_adj_4394, n26756, n743_adj_4395, n816_adj_4396, n889_adj_4397, 
        n317_adj_4398, n26755, n23_adj_4399, n25_adj_4400, n11_adj_4401, 
        n13_adj_4402, n15_adj_4403, n27_adj_4404, n9_adj_4405, n17_adj_4406, 
        n962_adj_4407, n904_adj_4408, n1035_adj_4409, n1108_adj_4410, 
        n244_adj_4411, n26754, n11_adj_4412, n25729, n9_adj_4414, 
        n25728, n25677, n19_adj_4416, n25676, n21_adj_4417, n171_adj_4418, 
        n26753, n7_adj_4419, n25727, n34214, n5_adj_4421, n25726, 
        n25675;
    wire [0:0]n7405;
    
    wire n25636, n24_adj_4423, n29_adj_4424, n98_adj_4425, n25635;
    wire [15:0]n9106;
    
    wire n26752, n12_adj_4426, n1117_adj_4427, n26751, n25674, n1044_adj_4428, 
        n26750, n89_adj_4429, n20_adj_4430, n971_adj_4431, n26749, 
        n162_adj_4432, n235_adj_4433, n25634, n898_adj_4434, n26748, 
        n825_adj_4435, n26747, n308_adj_4436, n381_adj_4437, n454_adj_4438, 
        n527_adj_4439, n752_adj_4440, n26746, n600_adj_4441, n673_adj_4442, 
        n25633, n3_adj_4443, n25725, n746_adj_4445, n819_adj_4446, 
        n892_adj_4447, n965_adj_4448, n25673, n25672, n25632, n25724, 
        n1038_adj_4451, n1111_adj_4452, n25671, n25631, n25723, n679_adj_4454, 
        n26745, n25670, n34156, n34154, n34664, n34739, n4_adj_4455, 
        n34778, n34779, n34166, n34164, n34869, n34741, n34916, 
        n34917, n34896, n34158, n34822, n40_adj_4456, n34824, n606_adj_4457, 
        n26744, n533_adj_4458, n26743, n460_adj_4459, n26742, n34227, 
        n6_adj_4460, n387_adj_4461, n26741, n92_adj_4462, n23_adj_4463, 
        n314_adj_4464, n26740, n165_adj_4465, n238_adj_4466, n311_adj_4467, 
        n384_adj_4468, n457_adj_4469, n530_adj_4470, n603_adj_4471, 
        n676_adj_4472, n241_adj_4473, n26739, n168_adj_4474, n26738, 
        n749_adj_4475, n26_adj_4476, n95_adj_4477;
    wire [16:0]n9087;
    
    wire n26737, n26736, n1114_adj_4478, n26735, n1041_adj_4479, n26734, 
        n822_adj_4480, n895_adj_4481, n968_adj_4483, n26733, n25669, 
        n26732, n25630, n26731, n25722, n26730, n26729, n25629, 
        n25668, n26728, n25667, n25721, n26727, n26726, n25666, 
        n26725, n26724, n26723, n26722, n25720;
    wire [17:0]n9067;
    
    wire n26721, n26720, n26719, n26718, n26717, n25719, n26716, 
        n26715, n26714, n25628, n26713, n26712, n26711, n26710, 
        n26709, n26708, n26707, n26706, n26705, n6_adj_4491;
    wire [3:0]n9256;
    wire [18:0]n9046;
    
    wire n26704, n26703, n26702, n25718, n25665;
    wire [1:0]n9267;
    
    wire n4_adj_4492;
    wire [2:0]n9262;
    
    wire n12_adj_4493, n8_adj_4494, n11_adj_4495, n26701, n6_adj_4496, 
        n25357, n18_adj_4497, n13_adj_4498, n25717, n34518, n26700, 
        n4_adj_4499, n26699, n26698, n26697, n26696, n26695, n25664, 
        n25716, n26694, n25627, n26693, n26692, n25715, n26691, 
        n25714, n26690, n26689, n26688, n26687, n25713, n25712, 
        n25663;
    wire [19:0]n9024;
    
    wire n26686, n26685, n26684, n26683, n26682, n26681, n25711, 
        n25710, n26680, n25662, n25626, n25625, n26679, n26678, 
        n26677, n26676, n26675, n26674, n26673, n26672, n25624, 
        n34493, n26671, n25709, n34806, n25661, n34650, n26670, 
        n26669, n26668;
    wire [20:0]n9001;
    
    wire n26667, n26666, n26665, n26664, n26663, n26662, n25623, 
        n26661, n26660, n26659, n26658, n26657, n26656, n26655, 
        n26654, n16_adj_4501, n25708, n25660, n25707, n25659, n25706, 
        n25658, n26653, n26652, n26651, n26650, n25770, n25769, 
        n25705, n25622, n25768, n26649, n26648;
    wire [21:0]n8977;
    
    wire n26647, n26646, n26645, n26644, n26643, n26642, n26641, 
        n26640, n26639, n26638, n25767, n26637, n26636, n26635, 
        n26634, n25657, n26633, n26632, n25621, n25766, n25704, 
        n26631, n34808, n25656, n26630, n26629, n26628, n8_adj_4504, 
        n26627, n26626, n26625, n26624, n26623, n26622, n26621, 
        n26620, n26619, n26618, n26617, n26616, n26615, n26614, 
        n26613, n26612, n26611, n26610, n26609, n26608, n26607, 
        n26606, n26605, n34809, n8_adj_4505, n24_adj_4506, n25765, 
        n25620, n25764, n34188, n4_adj_4507;
    wire [3:0]n9553;
    
    wire n6_adj_4508, n4_adj_4509;
    wire [4:0]n9546;
    wire [2:0]n9559;
    
    wire n25430, n4_adj_4510, n25763, n25703, n25655, n25762, n25702, 
        n25619, n25464;
    wire [1:0]n9564;
    
    wire n4_adj_4511, n25387;
    wire [5:0]n9538;
    
    wire n32845, n490_adj_4512, n27090, n417_adj_4513, n27089, n344_adj_4514, 
        n27088, n271_adj_4515, n27087, n198_adj_4516, n27086, n56_adj_4517, 
        n125_adj_4518;
    wire [6:0]n9529;
    
    wire n560_adj_4519, n27085, n487_adj_4520, n27084, n414_adj_4521, 
        n27083, n341_adj_4522, n27082, n268_adj_4523, n27081, n195_adj_4524, 
        n27080, n53_adj_4525, n122_adj_4526;
    wire [7:0]n9519;
    
    wire n630_adj_4527, n27079, n557_adj_4528, n27078, n484_adj_4529, 
        n27077, n411_adj_4530, n27076, n338_adj_4531, n27075, n265_adj_4532, 
        n27074, n192_adj_4533, n27073, n50_adj_4534, n119_adj_4535;
    wire [8:0]n9508;
    
    wire n700_adj_4536, n27072, n627_adj_4537, n27071, n554_adj_4538, 
        n27070, n481_adj_4539, n27069, n408_adj_4540, n27068, n335_adj_4541, 
        n27067, n262_adj_4542, n27066, n189_adj_4543, n27065, n47_adj_4544, 
        n116_adj_4545;
    wire [9:0]n9496;
    
    wire n770_adj_4546, n27064, n697_adj_4547, n27063, n624_adj_4548, 
        n27062, n551_adj_4549, n27061, n478_adj_4550, n27060, n17_adj_4551, 
        n405_adj_4552, n27059, n332_adj_4553, n27058, n259_adj_4554, 
        n27057, n186_adj_4555, n27056, n44_adj_4556, n113_adj_4557;
    wire [10:0]n9483;
    
    wire n840_adj_4558, n27055, n767_adj_4559, n27054, n694_adj_4560, 
        n27053, n621_adj_4561, n27052, n9_adj_4562, n548_adj_4563, 
        n27051, n11_adj_4564, n475_adj_4565, n27050, n34332, n402_adj_4566, 
        n27049, n34329, n329_adj_4567, n27048, n36254, n256_adj_4568, 
        n27047, n183_adj_4569, n27046, n41_adj_4570, n110_adj_4571, 
        n34698;
    wire [11:0]n9469;
    
    wire n910_adj_4572, n27045, n837_adj_4573, n27044, n34578, n764_adj_4574, 
        n27043, n691_adj_4575, n27042, n618_adj_4576, n27041, n36236, 
        n545_adj_4577, n27040, n472_adj_4578, n27039, n34576, n399_adj_4579, 
        n27038, n326_adj_4580, n27037, n34574, n253_adj_4581, n27036, 
        n180_adj_4582, n27035, n38_adj_4583, n107_adj_4584, n980_adj_4585, 
        n27034, n907_adj_4586, n27033, n834_adj_4587, n27032, n761_adj_4588, 
        n27031, n688_adj_4589, n27030, n615_adj_4590, n27029, n542_adj_4591, 
        n27028, n469_adj_4592, n27027, n396_adj_4593, n27026, n323_adj_4594, 
        n27025, n250_adj_4595, n27024, n177_adj_4596, n27023, n35_adj_4597, 
        n104_adj_4598, n1050_adj_4600, n27022, n977_adj_4601, n27021, 
        n36230, n34254, n34260, n25761, n16_adj_4605, n34229, n8_adj_4607, 
        n24_adj_4609, n34273, n25760, n34550, n25759, n25758, n34546, 
        n25757, n34832, n34676, n25756, n34863, n25755, n25618, 
        n25754, n25753, n34580, n36223, n34568, n36218, n12_adj_4613, 
        n34288, n36241, n10_adj_4614, n30_adj_4615, n34764, n34312, 
        n36221, n34692, n36247, n34837, n36212, n25617, n34891, 
        n36209, n16_adj_4616, n34275, n25752, n24_adj_4617, n6_adj_4618, 
        n34716, n34717, n34277, n36206, n34658, n34498, n4_adj_4619, 
        n34706, n34707, n12_adj_4620, n34240, n10_adj_4621, n30_adj_4622, 
        n34250, n34849, n34510, n34901, n34902, n34874, n6_adj_4623, 
        n34708, n34709, n34231, n34660, n34508, n34233, n34812, 
        n34516, n34861, n4_adj_4624, n34714, n34715, n34290, n34847, 
        n34500, n34899, n34900, n34878, n34279, n34810, n34506, 
        \PID_CONTROLLER.integral_23__N_3513 , n34859, n12_adj_4625, n8_adj_4626, 
        n11_adj_4627, n6_adj_4628, n25489, n18_adj_4629, n13_adj_4630, 
        n25332, n25298, n4_adj_4631, n25255;
    
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n25615), 
            .O(duty_23__N_3563[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5065_12 (.CI(n27019), .I0(n9454[9]), .I1(n831), .CO(n27020));
    SB_LUT4 add_5065_11_lut (.I0(GND_net), .I1(n9454[8]), .I2(n758), .I3(n27018), 
            .O(n9438[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5065_11 (.CI(n27018), .I0(n9454[8]), .I1(n758), .CO(n27019));
    SB_LUT4 add_5065_10_lut (.I0(GND_net), .I1(n9454[7]), .I2(n685), .I3(n27017), 
            .O(n9438[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_10 (.CI(n27017), .I0(n9454[7]), .I1(n685), .CO(n27018));
    SB_LUT4 add_5065_9_lut (.I0(GND_net), .I1(n9454[6]), .I2(n612), .I3(n27016), 
            .O(n9438[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_9 (.CI(n27016), .I0(n9454[6]), .I1(n612), .CO(n27017));
    SB_LUT4 add_5065_8_lut (.I0(GND_net), .I1(n9454[5]), .I2(n539_adj_4211), 
            .I3(n27015), .O(n9438[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_8 (.CI(n27015), .I0(n9454[5]), .I1(n539_adj_4211), 
            .CO(n27016));
    SB_LUT4 add_5065_7_lut (.I0(GND_net), .I1(n9454[4]), .I2(n466_adj_4212), 
            .I3(n27014), .O(n9438[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_7 (.CI(n27014), .I0(n9454[4]), .I1(n466_adj_4212), 
            .CO(n27015));
    SB_LUT4 add_5065_6_lut (.I0(GND_net), .I1(n9454[3]), .I2(n393_adj_4213), 
            .I3(n27013), .O(n9438[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_6 (.CI(n27013), .I0(n9454[3]), .I1(n393_adj_4213), 
            .CO(n27014));
    SB_LUT4 add_5065_5_lut (.I0(GND_net), .I1(n9454[2]), .I2(n320_adj_4214), 
            .I3(n27012), .O(n9438[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_5 (.CI(n27012), .I0(n9454[2]), .I1(n320_adj_4214), 
            .CO(n27013));
    SB_LUT4 add_5065_4_lut (.I0(GND_net), .I1(n9454[1]), .I2(n247_adj_4215), 
            .I3(n27011), .O(n9438[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4216));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4217));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5065_4 (.CI(n27011), .I0(n9454[1]), .I1(n247_adj_4215), 
            .CO(n27012));
    SB_LUT4 add_5065_3_lut (.I0(GND_net), .I1(n9454[0]), .I2(n174_adj_4218), 
            .I3(n27010), .O(n9438[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_3 (.CI(n27010), .I0(n9454[0]), .I1(n174_adj_4218), 
            .CO(n27011));
    SB_LUT4 add_5065_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n9438[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n27010));
    SB_LUT4 add_5064_16_lut (.I0(GND_net), .I1(n9438[13]), .I2(n1120), 
            .I3(n27009), .O(n9421[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5064_15_lut (.I0(GND_net), .I1(n9438[12]), .I2(n1047), 
            .I3(n27008), .O(n9421[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_15 (.CI(n27008), .I0(n9438[12]), .I1(n1047), .CO(n27009));
    SB_LUT4 add_5064_14_lut (.I0(GND_net), .I1(n9438[11]), .I2(n974), 
            .I3(n27007), .O(n9421[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_14 (.CI(n27007), .I0(n9438[11]), .I1(n974), .CO(n27008));
    SB_LUT4 add_5064_13_lut (.I0(GND_net), .I1(n9438[10]), .I2(n901), 
            .I3(n27006), .O(n9421[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_13 (.CI(n27006), .I0(n9438[10]), .I1(n901), .CO(n27007));
    SB_LUT4 add_5064_12_lut (.I0(GND_net), .I1(n9438[9]), .I2(n828), .I3(n27005), 
            .O(n9421[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_12 (.CI(n27005), .I0(n9438[9]), .I1(n828), .CO(n27006));
    SB_LUT4 add_5064_11_lut (.I0(GND_net), .I1(n9438[8]), .I2(n755), .I3(n27004), 
            .O(n9421[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_11 (.CI(n27004), .I0(n9438[8]), .I1(n755), .CO(n27005));
    SB_LUT4 add_5064_10_lut (.I0(GND_net), .I1(n9438[7]), .I2(n682), .I3(n27003), 
            .O(n9421[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_10 (.CI(n27003), .I0(n9438[7]), .I1(n682), .CO(n27004));
    SB_LUT4 add_5064_9_lut (.I0(GND_net), .I1(n9438[6]), .I2(n609), .I3(n27002), 
            .O(n9421[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_9 (.CI(n27002), .I0(n9438[6]), .I1(n609), .CO(n27003));
    SB_LUT4 add_5064_8_lut (.I0(GND_net), .I1(n9438[5]), .I2(n536), .I3(n27001), 
            .O(n9421[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_8 (.CI(n27001), .I0(n9438[5]), .I1(n536), .CO(n27002));
    SB_LUT4 add_5064_7_lut (.I0(GND_net), .I1(n9438[4]), .I2(n463), .I3(n27000), 
            .O(n9421[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_7 (.CI(n27000), .I0(n9438[4]), .I1(n463), .CO(n27001));
    SB_LUT4 add_5064_6_lut (.I0(GND_net), .I1(n9438[3]), .I2(n390), .I3(n26999), 
            .O(n9421[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_6 (.CI(n26999), .I0(n9438[3]), .I1(n390), .CO(n27000));
    SB_LUT4 add_5064_5_lut (.I0(GND_net), .I1(n9438[2]), .I2(n317), .I3(n26998), 
            .O(n9421[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_5 (.CI(n26998), .I0(n9438[2]), .I1(n317), .CO(n26999));
    SB_LUT4 add_5064_4_lut (.I0(GND_net), .I1(n9438[1]), .I2(n244), .I3(n26997), 
            .O(n9421[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_4 (.CI(n26997), .I0(n9438[1]), .I1(n244), .CO(n26998));
    SB_LUT4 add_5064_3_lut (.I0(GND_net), .I1(n9438[0]), .I2(n171), .I3(n26996), 
            .O(n9421[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_3 (.CI(n26996), .I0(n9438[0]), .I1(n171), .CO(n26997));
    SB_LUT4 add_5064_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n9421[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5064_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5064_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n26996));
    SB_LUT4 add_5063_17_lut (.I0(GND_net), .I1(n9421[14]), .I2(GND_net), 
            .I3(n26995), .O(n9403[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5063_16_lut (.I0(GND_net), .I1(n9421[13]), .I2(n1117), 
            .I3(n26994), .O(n9403[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_16 (.CI(n26994), .I0(n9421[13]), .I1(n1117), .CO(n26995));
    SB_LUT4 add_5063_15_lut (.I0(GND_net), .I1(n9421[12]), .I2(n1044), 
            .I3(n26993), .O(n9403[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_15 (.CI(n26993), .I0(n9421[12]), .I1(n1044), .CO(n26994));
    SB_LUT4 add_5063_14_lut (.I0(GND_net), .I1(n9421[11]), .I2(n971), 
            .I3(n26992), .O(n9403[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_14 (.CI(n26992), .I0(n9421[11]), .I1(n971), .CO(n26993));
    SB_LUT4 add_5063_13_lut (.I0(GND_net), .I1(n9421[10]), .I2(n898), 
            .I3(n26991), .O(n9403[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_13 (.CI(n26991), .I0(n9421[10]), .I1(n898), .CO(n26992));
    SB_LUT4 add_5063_12_lut (.I0(GND_net), .I1(n9421[9]), .I2(n825), .I3(n26990), 
            .O(n9403[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_12 (.CI(n26990), .I0(n9421[9]), .I1(n825), .CO(n26991));
    SB_LUT4 add_5063_11_lut (.I0(GND_net), .I1(n9421[8]), .I2(n752), .I3(n26989), 
            .O(n9403[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_11 (.CI(n26989), .I0(n9421[8]), .I1(n752), .CO(n26990));
    SB_LUT4 add_5063_10_lut (.I0(GND_net), .I1(n9421[7]), .I2(n679), .I3(n26988), 
            .O(n9403[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_10 (.CI(n26988), .I0(n9421[7]), .I1(n679), .CO(n26989));
    SB_LUT4 add_5063_9_lut (.I0(GND_net), .I1(n9421[6]), .I2(n606), .I3(n26987), 
            .O(n9403[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_9 (.CI(n26987), .I0(n9421[6]), .I1(n606), .CO(n26988));
    SB_LUT4 add_5063_8_lut (.I0(GND_net), .I1(n9421[5]), .I2(n533), .I3(n26986), 
            .O(n9403[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_8 (.CI(n26986), .I0(n9421[5]), .I1(n533), .CO(n26987));
    SB_LUT4 add_5063_7_lut (.I0(GND_net), .I1(n9421[4]), .I2(n460), .I3(n26985), 
            .O(n9403[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_7 (.CI(n26985), .I0(n9421[4]), .I1(n460), .CO(n26986));
    SB_LUT4 add_5063_6_lut (.I0(GND_net), .I1(n9421[3]), .I2(n387), .I3(n26984), 
            .O(n9403[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_6 (.CI(n26984), .I0(n9421[3]), .I1(n387), .CO(n26985));
    SB_LUT4 add_5063_5_lut (.I0(GND_net), .I1(n9421[2]), .I2(n314), .I3(n26983), 
            .O(n9403[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_5 (.CI(n26983), .I0(n9421[2]), .I1(n314), .CO(n26984));
    SB_LUT4 add_5063_4_lut (.I0(GND_net), .I1(n9421[1]), .I2(n241), .I3(n26982), 
            .O(n9403[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_4 (.CI(n26982), .I0(n9421[1]), .I1(n241), .CO(n26983));
    SB_LUT4 add_5063_3_lut (.I0(GND_net), .I1(n9421[0]), .I2(n168), .I3(n26981), 
            .O(n9403[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_3 (.CI(n26981), .I0(n9421[0]), .I1(n168), .CO(n26982));
    SB_LUT4 add_5063_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n9403[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5063_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5063_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n26981));
    SB_LUT4 add_5062_18_lut (.I0(GND_net), .I1(n9403[15]), .I2(GND_net), 
            .I3(n26980), .O(n9384[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5062_17_lut (.I0(GND_net), .I1(n9403[14]), .I2(GND_net), 
            .I3(n26979), .O(n9384[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_17 (.CI(n26979), .I0(n9403[14]), .I1(GND_net), .CO(n26980));
    SB_LUT4 add_5062_16_lut (.I0(GND_net), .I1(n9403[13]), .I2(n1114), 
            .I3(n26978), .O(n9384[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_16 (.CI(n26978), .I0(n9403[13]), .I1(n1114), .CO(n26979));
    SB_LUT4 add_5062_15_lut (.I0(GND_net), .I1(n9403[12]), .I2(n1041), 
            .I3(n26977), .O(n9384[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_15 (.CI(n26977), .I0(n9403[12]), .I1(n1041), .CO(n26978));
    SB_LUT4 add_5062_14_lut (.I0(GND_net), .I1(n9403[11]), .I2(n968), 
            .I3(n26976), .O(n9384[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_14 (.CI(n26976), .I0(n9403[11]), .I1(n968), .CO(n26977));
    SB_LUT4 add_5062_13_lut (.I0(GND_net), .I1(n9403[10]), .I2(n895), 
            .I3(n26975), .O(n9384[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_13 (.CI(n26975), .I0(n9403[10]), .I1(n895), .CO(n26976));
    SB_LUT4 add_5062_12_lut (.I0(GND_net), .I1(n9403[9]), .I2(n822), .I3(n26974), 
            .O(n9384[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_12 (.CI(n26974), .I0(n9403[9]), .I1(n822), .CO(n26975));
    SB_LUT4 add_5062_11_lut (.I0(GND_net), .I1(n9403[8]), .I2(n749), .I3(n26973), 
            .O(n9384[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_11 (.CI(n26973), .I0(n9403[8]), .I1(n749), .CO(n26974));
    SB_LUT4 add_5062_10_lut (.I0(GND_net), .I1(n9403[7]), .I2(n676), .I3(n26972), 
            .O(n9384[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_10 (.CI(n26972), .I0(n9403[7]), .I1(n676), .CO(n26973));
    SB_LUT4 add_5062_9_lut (.I0(GND_net), .I1(n9403[6]), .I2(n603), .I3(n26971), 
            .O(n9384[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_9 (.CI(n26971), .I0(n9403[6]), .I1(n603), .CO(n26972));
    SB_LUT4 add_5062_8_lut (.I0(GND_net), .I1(n9403[5]), .I2(n530), .I3(n26970), 
            .O(n9384[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_8 (.CI(n26970), .I0(n9403[5]), .I1(n530), .CO(n26971));
    SB_LUT4 add_5062_7_lut (.I0(GND_net), .I1(n9403[4]), .I2(n457), .I3(n26969), 
            .O(n9384[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_7 (.CI(n26969), .I0(n9403[4]), .I1(n457), .CO(n26970));
    SB_LUT4 add_5062_6_lut (.I0(GND_net), .I1(n9403[3]), .I2(n384), .I3(n26968), 
            .O(n9384[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_6 (.CI(n26968), .I0(n9403[3]), .I1(n384), .CO(n26969));
    SB_LUT4 add_5062_5_lut (.I0(GND_net), .I1(n9403[2]), .I2(n311), .I3(n26967), 
            .O(n9384[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_5 (.CI(n26967), .I0(n9403[2]), .I1(n311), .CO(n26968));
    SB_LUT4 add_5062_4_lut (.I0(GND_net), .I1(n9403[1]), .I2(n238), .I3(n26966), 
            .O(n9384[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_4 (.CI(n26966), .I0(n9403[1]), .I1(n238), .CO(n26967));
    SB_LUT4 add_5062_3_lut (.I0(GND_net), .I1(n9403[0]), .I2(n165), .I3(n26965), 
            .O(n9384[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_3 (.CI(n26965), .I0(n9403[0]), .I1(n165), .CO(n26966));
    SB_LUT4 add_5062_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n9384[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5062_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5062_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n26965));
    SB_LUT4 add_5061_19_lut (.I0(GND_net), .I1(n9384[16]), .I2(GND_net), 
            .I3(n26964), .O(n9364[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5061_18_lut (.I0(GND_net), .I1(n9384[15]), .I2(GND_net), 
            .I3(n26963), .O(n9364[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_18 (.CI(n26963), .I0(n9384[15]), .I1(GND_net), .CO(n26964));
    SB_LUT4 add_5061_17_lut (.I0(GND_net), .I1(n9384[14]), .I2(GND_net), 
            .I3(n26962), .O(n9364[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_17 (.CI(n26962), .I0(n9384[14]), .I1(GND_net), .CO(n26963));
    SB_LUT4 add_5061_16_lut (.I0(GND_net), .I1(n9384[13]), .I2(n1111), 
            .I3(n26961), .O(n9364[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_16 (.CI(n26961), .I0(n9384[13]), .I1(n1111), .CO(n26962));
    SB_LUT4 add_5061_15_lut (.I0(GND_net), .I1(n9384[12]), .I2(n1038), 
            .I3(n26960), .O(n9364[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_15 (.CI(n26960), .I0(n9384[12]), .I1(n1038), .CO(n26961));
    SB_LUT4 add_5061_14_lut (.I0(GND_net), .I1(n9384[11]), .I2(n965), 
            .I3(n26959), .O(n9364[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_14 (.CI(n26959), .I0(n9384[11]), .I1(n965), .CO(n26960));
    SB_LUT4 add_5061_13_lut (.I0(GND_net), .I1(n9384[10]), .I2(n892), 
            .I3(n26958), .O(n9364[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_13 (.CI(n26958), .I0(n9384[10]), .I1(n892), .CO(n26959));
    SB_LUT4 add_5061_12_lut (.I0(GND_net), .I1(n9384[9]), .I2(n819), .I3(n26957), 
            .O(n9364[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_12 (.CI(n26957), .I0(n9384[9]), .I1(n819), .CO(n26958));
    SB_LUT4 add_5061_11_lut (.I0(GND_net), .I1(n9384[8]), .I2(n746), .I3(n26956), 
            .O(n9364[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_11 (.CI(n26956), .I0(n9384[8]), .I1(n746), .CO(n26957));
    SB_LUT4 add_5061_10_lut (.I0(GND_net), .I1(n9384[7]), .I2(n673), .I3(n26955), 
            .O(n9364[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_10 (.CI(n26955), .I0(n9384[7]), .I1(n673), .CO(n26956));
    SB_LUT4 add_5061_9_lut (.I0(GND_net), .I1(n9384[6]), .I2(n600), .I3(n26954), 
            .O(n9364[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_9 (.CI(n26954), .I0(n9384[6]), .I1(n600), .CO(n26955));
    SB_LUT4 add_5061_8_lut (.I0(GND_net), .I1(n9384[5]), .I2(n527), .I3(n26953), 
            .O(n9364[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_8 (.CI(n26953), .I0(n9384[5]), .I1(n527), .CO(n26954));
    SB_LUT4 add_5061_7_lut (.I0(GND_net), .I1(n9384[4]), .I2(n454), .I3(n26952), 
            .O(n9364[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_7 (.CI(n26952), .I0(n9384[4]), .I1(n454), .CO(n26953));
    SB_LUT4 add_5061_6_lut (.I0(GND_net), .I1(n9384[3]), .I2(n381), .I3(n26951), 
            .O(n9364[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_6 (.CI(n26951), .I0(n9384[3]), .I1(n381), .CO(n26952));
    SB_LUT4 add_5061_5_lut (.I0(GND_net), .I1(n9384[2]), .I2(n308), .I3(n26950), 
            .O(n9364[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_5 (.CI(n26950), .I0(n9384[2]), .I1(n308), .CO(n26951));
    SB_LUT4 add_5061_4_lut (.I0(GND_net), .I1(n9384[1]), .I2(n235), .I3(n26949), 
            .O(n9364[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_4 (.CI(n26949), .I0(n9384[1]), .I1(n235), .CO(n26950));
    SB_LUT4 add_5061_3_lut (.I0(GND_net), .I1(n9384[0]), .I2(n162), .I3(n26948), 
            .O(n9364[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_3 (.CI(n26948), .I0(n9384[0]), .I1(n162), .CO(n26949));
    SB_LUT4 add_5061_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n9364[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5061_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5061_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n26948));
    SB_LUT4 add_5060_20_lut (.I0(GND_net), .I1(n9364[17]), .I2(GND_net), 
            .I3(n26947), .O(n9343[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5060_19_lut (.I0(GND_net), .I1(n9364[16]), .I2(GND_net), 
            .I3(n26946), .O(n9343[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_19 (.CI(n26946), .I0(n9364[16]), .I1(GND_net), .CO(n26947));
    SB_LUT4 add_5060_18_lut (.I0(GND_net), .I1(n9364[15]), .I2(GND_net), 
            .I3(n26945), .O(n9343[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_18 (.CI(n26945), .I0(n9364[15]), .I1(GND_net), .CO(n26946));
    SB_LUT4 add_5060_17_lut (.I0(GND_net), .I1(n9364[14]), .I2(GND_net), 
            .I3(n26944), .O(n9343[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_17 (.CI(n26944), .I0(n9364[14]), .I1(GND_net), .CO(n26945));
    SB_LUT4 add_5060_16_lut (.I0(GND_net), .I1(n9364[13]), .I2(n1108), 
            .I3(n26943), .O(n9343[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_16 (.CI(n26943), .I0(n9364[13]), .I1(n1108), .CO(n26944));
    SB_LUT4 add_5060_15_lut (.I0(GND_net), .I1(n9364[12]), .I2(n1035), 
            .I3(n26942), .O(n9343[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_15 (.CI(n26942), .I0(n9364[12]), .I1(n1035), .CO(n26943));
    SB_LUT4 add_5060_14_lut (.I0(GND_net), .I1(n9364[11]), .I2(n962), 
            .I3(n26941), .O(n9343[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_14 (.CI(n26941), .I0(n9364[11]), .I1(n962), .CO(n26942));
    SB_LUT4 add_5060_13_lut (.I0(GND_net), .I1(n9364[10]), .I2(n889), 
            .I3(n26940), .O(n9343[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_13 (.CI(n26940), .I0(n9364[10]), .I1(n889), .CO(n26941));
    SB_LUT4 add_5060_12_lut (.I0(GND_net), .I1(n9364[9]), .I2(n816), .I3(n26939), 
            .O(n9343[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_12 (.CI(n26939), .I0(n9364[9]), .I1(n816), .CO(n26940));
    SB_LUT4 add_5060_11_lut (.I0(GND_net), .I1(n9364[8]), .I2(n743), .I3(n26938), 
            .O(n9343[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_11 (.CI(n26938), .I0(n9364[8]), .I1(n743), .CO(n26939));
    SB_LUT4 add_5060_10_lut (.I0(GND_net), .I1(n9364[7]), .I2(n670), .I3(n26937), 
            .O(n9343[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_10 (.CI(n26937), .I0(n9364[7]), .I1(n670), .CO(n26938));
    SB_LUT4 add_5060_9_lut (.I0(GND_net), .I1(n9364[6]), .I2(n597), .I3(n26936), 
            .O(n9343[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_9 (.CI(n26936), .I0(n9364[6]), .I1(n597), .CO(n26937));
    SB_LUT4 add_5060_8_lut (.I0(GND_net), .I1(n9364[5]), .I2(n524), .I3(n26935), 
            .O(n9343[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_8 (.CI(n26935), .I0(n9364[5]), .I1(n524), .CO(n26936));
    SB_LUT4 add_5060_7_lut (.I0(GND_net), .I1(n9364[4]), .I2(n451), .I3(n26934), 
            .O(n9343[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_7 (.CI(n26934), .I0(n9364[4]), .I1(n451), .CO(n26935));
    SB_LUT4 add_5060_6_lut (.I0(GND_net), .I1(n9364[3]), .I2(n378), .I3(n26933), 
            .O(n9343[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_6 (.CI(n26933), .I0(n9364[3]), .I1(n378), .CO(n26934));
    SB_LUT4 add_5060_5_lut (.I0(GND_net), .I1(n9364[2]), .I2(n305), .I3(n26932), 
            .O(n9343[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_5 (.CI(n26932), .I0(n9364[2]), .I1(n305), .CO(n26933));
    SB_LUT4 add_5060_4_lut (.I0(GND_net), .I1(n9364[1]), .I2(n232), .I3(n26931), 
            .O(n9343[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_4 (.CI(n26931), .I0(n9364[1]), .I1(n232), .CO(n26932));
    SB_LUT4 add_5060_3_lut (.I0(GND_net), .I1(n9364[0]), .I2(n159), .I3(n26930), 
            .O(n9343[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_3 (.CI(n26930), .I0(n9364[0]), .I1(n159), .CO(n26931));
    SB_LUT4 add_5060_2_lut (.I0(GND_net), .I1(n17_adj_4219), .I2(n86), 
            .I3(GND_net), .O(n9343[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5060_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5060_2 (.CI(GND_net), .I0(n17_adj_4219), .I1(n86), .CO(n26930));
    SB_LUT4 add_5059_21_lut (.I0(GND_net), .I1(n9343[18]), .I2(GND_net), 
            .I3(n26929), .O(n9321[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5059_20_lut (.I0(GND_net), .I1(n9343[17]), .I2(GND_net), 
            .I3(n26928), .O(n9321[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_20 (.CI(n26928), .I0(n9343[17]), .I1(GND_net), .CO(n26929));
    SB_LUT4 add_5059_19_lut (.I0(GND_net), .I1(n9343[16]), .I2(GND_net), 
            .I3(n26927), .O(n9321[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_19 (.CI(n26927), .I0(n9343[16]), .I1(GND_net), .CO(n26928));
    SB_LUT4 add_5059_18_lut (.I0(GND_net), .I1(n9343[15]), .I2(GND_net), 
            .I3(n26926), .O(n9321[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_18 (.CI(n26926), .I0(n9343[15]), .I1(GND_net), .CO(n26927));
    SB_LUT4 add_5059_17_lut (.I0(GND_net), .I1(n9343[14]), .I2(GND_net), 
            .I3(n26925), .O(n9321[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_17 (.CI(n26925), .I0(n9343[14]), .I1(GND_net), .CO(n26926));
    SB_LUT4 add_5059_16_lut (.I0(GND_net), .I1(n9343[13]), .I2(n1105), 
            .I3(n26924), .O(n9321[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_16 (.CI(n26924), .I0(n9343[13]), .I1(n1105), .CO(n26925));
    SB_LUT4 add_5059_15_lut (.I0(GND_net), .I1(n9343[12]), .I2(n1032), 
            .I3(n26923), .O(n9321[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_15 (.CI(n26923), .I0(n9343[12]), .I1(n1032), .CO(n26924));
    SB_LUT4 add_5059_14_lut (.I0(GND_net), .I1(n9343[11]), .I2(n959), 
            .I3(n26922), .O(n9321[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_14 (.CI(n26922), .I0(n9343[11]), .I1(n959), .CO(n26923));
    SB_LUT4 add_5059_13_lut (.I0(GND_net), .I1(n9343[10]), .I2(n886), 
            .I3(n26921), .O(n9321[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_13 (.CI(n26921), .I0(n9343[10]), .I1(n886), .CO(n26922));
    SB_LUT4 add_5059_12_lut (.I0(GND_net), .I1(n9343[9]), .I2(n813), .I3(n26920), 
            .O(n9321[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_12 (.CI(n26920), .I0(n9343[9]), .I1(n813), .CO(n26921));
    SB_LUT4 add_5059_11_lut (.I0(GND_net), .I1(n9343[8]), .I2(n740), .I3(n26919), 
            .O(n9321[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_11 (.CI(n26919), .I0(n9343[8]), .I1(n740), .CO(n26920));
    SB_LUT4 add_5059_10_lut (.I0(GND_net), .I1(n9343[7]), .I2(n667), .I3(n26918), 
            .O(n9321[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_10 (.CI(n26918), .I0(n9343[7]), .I1(n667), .CO(n26919));
    SB_LUT4 add_5059_9_lut (.I0(GND_net), .I1(n9343[6]), .I2(n594), .I3(n26917), 
            .O(n9321[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_9 (.CI(n26917), .I0(n9343[6]), .I1(n594), .CO(n26918));
    SB_LUT4 add_5059_8_lut (.I0(GND_net), .I1(n9343[5]), .I2(n521), .I3(n26916), 
            .O(n9321[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_8 (.CI(n26916), .I0(n9343[5]), .I1(n521), .CO(n26917));
    SB_LUT4 add_5059_7_lut (.I0(GND_net), .I1(n9343[4]), .I2(n448), .I3(n26915), 
            .O(n9321[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_7 (.CI(n26915), .I0(n9343[4]), .I1(n448), .CO(n26916));
    SB_LUT4 add_5059_6_lut (.I0(GND_net), .I1(n9343[3]), .I2(n375), .I3(n26914), 
            .O(n9321[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_6 (.CI(n26914), .I0(n9343[3]), .I1(n375), .CO(n26915));
    SB_LUT4 add_5059_5_lut (.I0(GND_net), .I1(n9343[2]), .I2(n302), .I3(n26913), 
            .O(n9321[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_5 (.CI(n26913), .I0(n9343[2]), .I1(n302), .CO(n26914));
    SB_LUT4 add_5059_4_lut (.I0(GND_net), .I1(n9343[1]), .I2(n229), .I3(n26912), 
            .O(n9321[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_4 (.CI(n26912), .I0(n9343[1]), .I1(n229), .CO(n26913));
    SB_LUT4 add_5059_3_lut (.I0(GND_net), .I1(n9343[0]), .I2(n156), .I3(n26911), 
            .O(n9321[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_3 (.CI(n26911), .I0(n9343[0]), .I1(n156), .CO(n26912));
    SB_LUT4 add_5059_2_lut (.I0(GND_net), .I1(n14_adj_4220), .I2(n83), 
            .I3(GND_net), .O(n9321[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5059_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5059_2 (.CI(GND_net), .I0(n14_adj_4220), .I1(n83), .CO(n26911));
    SB_LUT4 add_5058_22_lut (.I0(GND_net), .I1(n9321[19]), .I2(GND_net), 
            .I3(n26910), .O(n9298[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5058_21_lut (.I0(GND_net), .I1(n9321[18]), .I2(GND_net), 
            .I3(n26909), .O(n9298[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_21 (.CI(n26909), .I0(n9321[18]), .I1(GND_net), .CO(n26910));
    SB_LUT4 add_5058_20_lut (.I0(GND_net), .I1(n9321[17]), .I2(GND_net), 
            .I3(n26908), .O(n9298[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_20 (.CI(n26908), .I0(n9321[17]), .I1(GND_net), .CO(n26909));
    SB_LUT4 add_5058_19_lut (.I0(GND_net), .I1(n9321[16]), .I2(GND_net), 
            .I3(n26907), .O(n9298[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_19 (.CI(n26907), .I0(n9321[16]), .I1(GND_net), .CO(n26908));
    SB_LUT4 add_5058_18_lut (.I0(GND_net), .I1(n9321[15]), .I2(GND_net), 
            .I3(n26906), .O(n9298[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_18 (.CI(n26906), .I0(n9321[15]), .I1(GND_net), .CO(n26907));
    SB_LUT4 add_5058_17_lut (.I0(GND_net), .I1(n9321[14]), .I2(GND_net), 
            .I3(n26905), .O(n9298[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_17 (.CI(n26905), .I0(n9321[14]), .I1(GND_net), .CO(n26906));
    SB_LUT4 add_5058_16_lut (.I0(GND_net), .I1(n9321[13]), .I2(n1102), 
            .I3(n26904), .O(n9298[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_16 (.CI(n26904), .I0(n9321[13]), .I1(n1102), .CO(n26905));
    SB_LUT4 add_5058_15_lut (.I0(GND_net), .I1(n9321[12]), .I2(n1029), 
            .I3(n26903), .O(n9298[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_15 (.CI(n26903), .I0(n9321[12]), .I1(n1029), .CO(n26904));
    SB_LUT4 add_5058_14_lut (.I0(GND_net), .I1(n9321[11]), .I2(n956), 
            .I3(n26902), .O(n9298[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_14 (.CI(n26902), .I0(n9321[11]), .I1(n956), .CO(n26903));
    SB_LUT4 add_5058_13_lut (.I0(GND_net), .I1(n9321[10]), .I2(n883), 
            .I3(n26901), .O(n9298[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_13 (.CI(n26901), .I0(n9321[10]), .I1(n883), .CO(n26902));
    SB_LUT4 add_5058_12_lut (.I0(GND_net), .I1(n9321[9]), .I2(n810), .I3(n26900), 
            .O(n9298[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_12 (.CI(n26900), .I0(n9321[9]), .I1(n810), .CO(n26901));
    SB_LUT4 add_5058_11_lut (.I0(GND_net), .I1(n9321[8]), .I2(n737), .I3(n26899), 
            .O(n9298[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_11 (.CI(n26899), .I0(n9321[8]), .I1(n737), .CO(n26900));
    SB_LUT4 add_5058_10_lut (.I0(GND_net), .I1(n9321[7]), .I2(n664), .I3(n26898), 
            .O(n9298[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_10 (.CI(n26898), .I0(n9321[7]), .I1(n664), .CO(n26899));
    SB_LUT4 add_5058_9_lut (.I0(GND_net), .I1(n9321[6]), .I2(n591), .I3(n26897), 
            .O(n9298[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_9 (.CI(n26897), .I0(n9321[6]), .I1(n591), .CO(n26898));
    SB_LUT4 add_5058_8_lut (.I0(GND_net), .I1(n9321[5]), .I2(n518), .I3(n26896), 
            .O(n9298[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_8 (.CI(n26896), .I0(n9321[5]), .I1(n518), .CO(n26897));
    SB_LUT4 add_5058_7_lut (.I0(GND_net), .I1(n9321[4]), .I2(n445), .I3(n26895), 
            .O(n9298[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_7 (.CI(n26895), .I0(n9321[4]), .I1(n445), .CO(n26896));
    SB_LUT4 add_5058_6_lut (.I0(GND_net), .I1(n9321[3]), .I2(n372), .I3(n26894), 
            .O(n9298[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_6 (.CI(n26894), .I0(n9321[3]), .I1(n372), .CO(n26895));
    SB_LUT4 add_5058_5_lut (.I0(GND_net), .I1(n9321[2]), .I2(n299), .I3(n26893), 
            .O(n9298[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_5 (.CI(n26893), .I0(n9321[2]), .I1(n299), .CO(n26894));
    SB_LUT4 add_5058_4_lut (.I0(GND_net), .I1(n9321[1]), .I2(n226), .I3(n26892), 
            .O(n9298[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_4 (.CI(n26892), .I0(n9321[1]), .I1(n226), .CO(n26893));
    SB_LUT4 add_5058_3_lut (.I0(GND_net), .I1(n9321[0]), .I2(n153), .I3(n26891), 
            .O(n9298[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_3 (.CI(n26891), .I0(n9321[0]), .I1(n153), .CO(n26892));
    SB_LUT4 add_5058_2_lut (.I0(GND_net), .I1(n11_adj_4221), .I2(n80), 
            .I3(GND_net), .O(n9298[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5058_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5058_2 (.CI(GND_net), .I0(n11_adj_4221), .I1(n80), .CO(n26891));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3463 [23]), 
            .I1(n9274[21]), .I2(GND_net), .I3(n26890), .O(n7409[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9274[20]), .I2(GND_net), 
            .I3(n26889), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n26889), .I0(n9274[20]), .I1(GND_net), 
            .CO(n26890));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9274[19]), .I2(GND_net), 
            .I3(n26888), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n26888), .I0(n9274[19]), .I1(GND_net), 
            .CO(n26889));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9274[18]), .I2(GND_net), 
            .I3(n26887), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n26887), .I0(n9274[18]), .I1(GND_net), 
            .CO(n26888));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9274[17]), .I2(GND_net), 
            .I3(n26886), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n26886), .I0(n9274[17]), .I1(GND_net), 
            .CO(n26887));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9274[16]), .I2(GND_net), 
            .I3(n26885), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n26885), .I0(n9274[16]), .I1(GND_net), 
            .CO(n26886));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9274[15]), .I2(GND_net), 
            .I3(n26884), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n26884), .I0(n9274[15]), .I1(GND_net), 
            .CO(n26885));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9274[14]), .I2(GND_net), 
            .I3(n26883), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n26883), .I0(n9274[14]), .I1(GND_net), 
            .CO(n26884));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9274[13]), .I2(n1096), 
            .I3(n26882), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n26882), .I0(n9274[13]), .I1(n1096), 
            .CO(n26883));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9274[12]), .I2(n1023), 
            .I3(n26881), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n26881), .I0(n9274[12]), .I1(n1023), 
            .CO(n26882));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9274[11]), .I2(n950), 
            .I3(n26880), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n26880), .I0(n9274[11]), .I1(n950), 
            .CO(n26881));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9274[10]), .I2(n877), 
            .I3(n26879), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n26879), .I0(n9274[10]), .I1(n877), 
            .CO(n26880));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9274[9]), .I2(n804), 
            .I3(n26878), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n26878), .I0(n9274[9]), .I1(n804), 
            .CO(n26879));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9274[8]), .I2(n731), 
            .I3(n26877), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n26877), .I0(n9274[8]), .I1(n731), 
            .CO(n26878));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9274[7]), .I2(n658), 
            .I3(n26876), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n26876), .I0(n9274[7]), .I1(n658), 
            .CO(n26877));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9274[6]), .I2(n585), 
            .I3(n26875), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n26875), .I0(n9274[6]), .I1(n585), 
            .CO(n26876));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9274[5]), .I2(n512), 
            .I3(n26874), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n26874), .I0(n9274[5]), .I1(n512), 
            .CO(n26875));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9274[4]), .I2(n439), 
            .I3(n26873), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n26873), .I0(n9274[4]), .I1(n439), 
            .CO(n26874));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9274[3]), .I2(n366), 
            .I3(n26872), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n26872), .I0(n9274[3]), .I1(n366), 
            .CO(n26873));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9274[2]), .I2(n293), 
            .I3(n26871), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n26871), .I0(n9274[2]), .I1(n293), 
            .CO(n26872));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9274[1]), .I2(n220), 
            .I3(n26870), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n26870), .I0(n9274[1]), .I1(n220), 
            .CO(n26871));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9274[0]), .I2(n147), 
            .I3(n26869), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n26869), .I0(n9274[0]), .I1(n147), 
            .CO(n26870));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n26869));
    SB_LUT4 add_5057_23_lut (.I0(GND_net), .I1(n9298[20]), .I2(GND_net), 
            .I3(n26868), .O(n9274[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5057_22_lut (.I0(GND_net), .I1(n9298[19]), .I2(GND_net), 
            .I3(n26867), .O(n9274[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_22 (.CI(n26867), .I0(n9298[19]), .I1(GND_net), .CO(n26868));
    SB_LUT4 add_5057_21_lut (.I0(GND_net), .I1(n9298[18]), .I2(GND_net), 
            .I3(n26866), .O(n9274[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_21 (.CI(n26866), .I0(n9298[18]), .I1(GND_net), .CO(n26867));
    SB_LUT4 add_5057_20_lut (.I0(GND_net), .I1(n9298[17]), .I2(GND_net), 
            .I3(n26865), .O(n9274[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_20 (.CI(n26865), .I0(n9298[17]), .I1(GND_net), .CO(n26866));
    SB_LUT4 add_5057_19_lut (.I0(GND_net), .I1(n9298[16]), .I2(GND_net), 
            .I3(n26864), .O(n9274[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_19 (.CI(n26864), .I0(n9298[16]), .I1(GND_net), .CO(n26865));
    SB_LUT4 add_5057_18_lut (.I0(GND_net), .I1(n9298[15]), .I2(GND_net), 
            .I3(n26863), .O(n9274[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_18 (.CI(n26863), .I0(n9298[15]), .I1(GND_net), .CO(n26864));
    SB_LUT4 add_5057_17_lut (.I0(GND_net), .I1(n9298[14]), .I2(GND_net), 
            .I3(n26862), .O(n9274[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_17 (.CI(n26862), .I0(n9298[14]), .I1(GND_net), .CO(n26863));
    SB_LUT4 add_5057_16_lut (.I0(GND_net), .I1(n9298[13]), .I2(n1099), 
            .I3(n26861), .O(n9274[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_16 (.CI(n26861), .I0(n9298[13]), .I1(n1099), .CO(n26862));
    SB_LUT4 add_5057_15_lut (.I0(GND_net), .I1(n9298[12]), .I2(n1026), 
            .I3(n26860), .O(n9274[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_15 (.CI(n26860), .I0(n9298[12]), .I1(n1026), .CO(n26861));
    SB_LUT4 add_5057_14_lut (.I0(GND_net), .I1(n9298[11]), .I2(n953), 
            .I3(n26859), .O(n9274[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_14 (.CI(n26859), .I0(n9298[11]), .I1(n953), .CO(n26860));
    SB_LUT4 add_5057_13_lut (.I0(GND_net), .I1(n9298[10]), .I2(n880), 
            .I3(n26858), .O(n9274[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_13 (.CI(n26858), .I0(n9298[10]), .I1(n880), .CO(n26859));
    SB_LUT4 add_5057_12_lut (.I0(GND_net), .I1(n9298[9]), .I2(n807), .I3(n26857), 
            .O(n9274[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_12 (.CI(n26857), .I0(n9298[9]), .I1(n807), .CO(n26858));
    SB_LUT4 add_5057_11_lut (.I0(GND_net), .I1(n9298[8]), .I2(n734), .I3(n26856), 
            .O(n9274[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_11 (.CI(n26856), .I0(n9298[8]), .I1(n734), .CO(n26857));
    SB_LUT4 add_5057_10_lut (.I0(GND_net), .I1(n9298[7]), .I2(n661), .I3(n26855), 
            .O(n9274[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_10 (.CI(n26855), .I0(n9298[7]), .I1(n661), .CO(n26856));
    SB_LUT4 add_5057_9_lut (.I0(GND_net), .I1(n9298[6]), .I2(n588), .I3(n26854), 
            .O(n9274[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_9 (.CI(n26854), .I0(n9298[6]), .I1(n588), .CO(n26855));
    SB_LUT4 add_5057_8_lut (.I0(GND_net), .I1(n9298[5]), .I2(n515), .I3(n26853), 
            .O(n9274[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_8 (.CI(n26853), .I0(n9298[5]), .I1(n515), .CO(n26854));
    SB_LUT4 add_5057_7_lut (.I0(GND_net), .I1(n9298[4]), .I2(n442), .I3(n26852), 
            .O(n9274[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_7 (.CI(n26852), .I0(n9298[4]), .I1(n442), .CO(n26853));
    SB_LUT4 add_5057_6_lut (.I0(GND_net), .I1(n9298[3]), .I2(n369), .I3(n26851), 
            .O(n9274[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_6 (.CI(n26851), .I0(n9298[3]), .I1(n369), .CO(n26852));
    SB_LUT4 add_5057_5_lut (.I0(GND_net), .I1(n9298[2]), .I2(n296), .I3(n26850), 
            .O(n9274[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_5 (.CI(n26850), .I0(n9298[2]), .I1(n296), .CO(n26851));
    SB_LUT4 add_5057_4_lut (.I0(GND_net), .I1(n9298[1]), .I2(n223), .I3(n26849), 
            .O(n9274[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_4 (.CI(n26849), .I0(n9298[1]), .I1(n223), .CO(n26850));
    SB_LUT4 add_5057_3_lut (.I0(GND_net), .I1(n9298[0]), .I2(n150), .I3(n26848), 
            .O(n9274[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_3 (.CI(n26848), .I0(n9298[0]), .I1(n150), .CO(n26849));
    SB_LUT4 add_5057_2_lut (.I0(GND_net), .I1(n8), .I2(n77), .I3(GND_net), 
            .O(n9274[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5057_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5057_2 (.CI(GND_net), .I0(n8), .I1(n77), .CO(n26848));
    SB_LUT4 add_5051_7_lut (.I0(GND_net), .I1(n32507), .I2(n490), .I3(n26847), 
            .O(n9241[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5051_6_lut (.I0(GND_net), .I1(n9249[3]), .I2(n417), .I3(n26846), 
            .O(n9241[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5051_6 (.CI(n26846), .I0(n9249[3]), .I1(n417), .CO(n26847));
    SB_LUT4 add_5051_5_lut (.I0(GND_net), .I1(n9249[2]), .I2(n344), .I3(n26845), 
            .O(n9241[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5051_5 (.CI(n26845), .I0(n9249[2]), .I1(n344), .CO(n26846));
    SB_LUT4 add_5051_4_lut (.I0(GND_net), .I1(n9249[1]), .I2(n271), .I3(n26844), 
            .O(n9241[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5051_4 (.CI(n26844), .I0(n9249[1]), .I1(n271), .CO(n26845));
    SB_LUT4 add_5051_3_lut (.I0(GND_net), .I1(n9249[0]), .I2(n198_adj_4222), 
            .I3(n26843), .O(n9241[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5051_3 (.CI(n26843), .I0(n9249[0]), .I1(n198_adj_4222), 
            .CO(n26844));
    SB_LUT4 add_5051_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n9241[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5051_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5051_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n26843));
    SB_LUT4 add_5050_8_lut (.I0(GND_net), .I1(n9241[5]), .I2(n560), .I3(n26842), 
            .O(n9232[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4224));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5050_7_lut (.I0(GND_net), .I1(n9241[4]), .I2(n487), .I3(n26841), 
            .O(n9232[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_7 (.CI(n26841), .I0(n9241[4]), .I1(n487), .CO(n26842));
    SB_LUT4 add_5050_6_lut (.I0(GND_net), .I1(n9241[3]), .I2(n414), .I3(n26840), 
            .O(n9232[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_6 (.CI(n26840), .I0(n9241[3]), .I1(n414), .CO(n26841));
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5050_5_lut (.I0(GND_net), .I1(n9241[2]), .I2(n341), .I3(n26839), 
            .O(n9232[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17345_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17815_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17815_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5050_5 (.CI(n26839), .I0(n9241[2]), .I1(n341), .CO(n26840));
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5050_4_lut (.I0(GND_net), .I1(n9241[1]), .I2(n268), .I3(n26838), 
            .O(n9232[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_4 (.CI(n26838), .I0(n9241[1]), .I1(n268), .CO(n26839));
    SB_LUT4 add_5050_3_lut (.I0(GND_net), .I1(n9241[0]), .I2(n195_adj_4231), 
            .I3(n26837), .O(n9232[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_3 (.CI(n26837), .I0(n9241[0]), .I1(n195_adj_4231), 
            .CO(n26838));
    SB_LUT4 add_5050_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n9232[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n26837));
    SB_LUT4 add_5049_9_lut (.I0(GND_net), .I1(n9232[6]), .I2(n630), .I3(n26836), 
            .O(n9222[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5049_8_lut (.I0(GND_net), .I1(n9232[5]), .I2(n557), .I3(n26835), 
            .O(n9222[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_8 (.CI(n26835), .I0(n9232[5]), .I1(n557), .CO(n26836));
    SB_LUT4 add_5049_7_lut (.I0(GND_net), .I1(n9232[4]), .I2(n484), .I3(n26834), 
            .O(n9222[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_7 (.CI(n26834), .I0(n9232[4]), .I1(n484), .CO(n26835));
    SB_LUT4 add_5049_6_lut (.I0(GND_net), .I1(n9232[3]), .I2(n411), .I3(n26833), 
            .O(n9222[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_6 (.CI(n26833), .I0(n9232[3]), .I1(n411), .CO(n26834));
    SB_LUT4 add_5049_5_lut (.I0(GND_net), .I1(n9232[2]), .I2(n338), .I3(n26832), 
            .O(n9222[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28627_3_lut (.I0(n34800), .I1(duty_23__N_3563[14]), .I2(n29_adj_4232), 
            .I3(GND_net), .O(n34801));   // verilog/motorControl.v(36[10:25])
    defparam i28627_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5049_5 (.CI(n26832), .I0(n9232[2]), .I1(n338), .CO(n26833));
    SB_LUT4 add_5049_4_lut (.I0(GND_net), .I1(n9232[1]), .I2(n265), .I3(n26831), 
            .O(n9222[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_4 (.CI(n26831), .I0(n9232[1]), .I1(n265), .CO(n26832));
    SB_LUT4 add_5049_3_lut (.I0(GND_net), .I1(n9232[0]), .I2(n192_adj_4233), 
            .I3(n26830), .O(n9222[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_3 (.CI(n26830), .I0(n9232[0]), .I1(n192_adj_4233), 
            .CO(n26831));
    SB_LUT4 add_5049_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n9222[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5049_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5049_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n26830));
    SB_LUT4 add_5048_10_lut (.I0(GND_net), .I1(n9222[7]), .I2(n700), .I3(n26829), 
            .O(n9211[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5048_9_lut (.I0(GND_net), .I1(n9222[6]), .I2(n627), .I3(n26828), 
            .O(n9211[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5048_9 (.CI(n26828), .I0(n9222[6]), .I1(n627), .CO(n26829));
    SB_LUT4 add_5048_8_lut (.I0(GND_net), .I1(n9222[5]), .I2(n554), .I3(n26827), 
            .O(n9211[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5048_8 (.CI(n26827), .I0(n9222[5]), .I1(n554), .CO(n26828));
    SB_LUT4 add_5048_7_lut (.I0(GND_net), .I1(n9222[4]), .I2(n481), .I3(n26826), 
            .O(n9211[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5048_7 (.CI(n26826), .I0(n9222[4]), .I1(n481), .CO(n26827));
    SB_LUT4 add_5048_6_lut (.I0(GND_net), .I1(n9222[3]), .I2(n408), .I3(n26825), 
            .O(n9211[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28029_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4232), .I3(n34207), 
            .O(n34201));
    defparam i28029_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5048_6 (.CI(n26825), .I0(n9222[3]), .I1(n408), .CO(n26826));
    SB_LUT4 i28693_4_lut (.I0(n30), .I1(n10_adj_4234), .I2(n35_adj_4235), 
            .I3(n34199), .O(n34867));   // verilog/motorControl.v(36[10:25])
    defparam i28693_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_4 (.CI(n25615), .I0(n106[2]), .I1(n155[2]), .CO(n25616));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n25750), .I0(GND_net), .I1(n1_adj_4633[3]), 
            .CO(n25751));
    SB_LUT4 add_5048_5_lut (.I0(GND_net), .I1(n9222[2]), .I2(n335), .I3(n26824), 
            .O(n9211[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5048_5 (.CI(n26824), .I0(n9222[2]), .I1(n335), .CO(n26825));
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5048_4_lut (.I0(GND_net), .I1(n9222[1]), .I2(n262), .I3(n26823), 
            .O(n9211[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5048_4 (.CI(n26823), .I0(n9222[1]), .I1(n262), .CO(n26824));
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4240));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5048_3_lut (.I0(GND_net), .I1(n9222[0]), .I2(n189_adj_4241), 
            .I3(n26822), .O(n9211[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5048_3 (.CI(n26822), .I0(n9222[0]), .I1(n189_adj_4241), 
            .CO(n26823));
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5048_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n9211[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5048_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5048_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n26822));
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3563[23]), .I1(n257[23]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3538[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3563[22]), .I1(n257[22]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3538[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3563[21]), .I1(n257[21]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3538[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_11_lut (.I0(GND_net), .I1(n9211[8]), .I2(n770), .I3(n26821), 
            .O(n9199[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3563[20]), .I1(n257[20]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[2]), 
            .I3(n25749), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3538[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_10_lut (.I0(GND_net), .I1(n9211[7]), .I2(n697), .I3(n26820), 
            .O(n9199[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5047_10 (.CI(n26820), .I0(n9211[7]), .I1(n697), .CO(n26821));
    SB_LUT4 i28561_3_lut (.I0(n34801), .I1(duty_23__N_3563[15]), .I2(n31), 
            .I3(GND_net), .O(n34735));   // verilog/motorControl.v(36[10:25])
    defparam i28561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_9_lut (.I0(GND_net), .I1(n9211[6]), .I2(n624), .I3(n26819), 
            .O(n9199[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3439[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3563[19]), .I1(n257[19]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3538[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5047_9 (.CI(n26819), .I0(n9211[6]), .I1(n624), .CO(n26820));
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3563[18]), .I1(n257[18]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n25614), 
            .O(duty_23__N_3563[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5047_8_lut (.I0(GND_net), .I1(n9211[5]), .I2(n551), .I3(n26818), 
            .O(n9199[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_3 (.CI(n25614), .I0(n106[1]), .I1(n155[1]), .CO(n25615));
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3538[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n25749), .I0(GND_net), .I1(n1_adj_4633[2]), 
            .CO(n25750));
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3563[17]), .I1(n257[17]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3538[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5047_8 (.CI(n26818), .I0(n9211[5]), .I1(n551), .CO(n26819));
    SB_LUT4 add_5047_7_lut (.I0(GND_net), .I1(n9211[4]), .I2(n478), .I3(n26817), 
            .O(n9199[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3563[16]), .I1(n257[16]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3538[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3563[15]), .I1(n257[15]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3538[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3563[14]), .I1(n257[14]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5047_7 (.CI(n26817), .I0(n9211[4]), .I1(n478), .CO(n26818));
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3538[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3563[13]), .I1(n257[13]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3538[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_6_lut (.I0(GND_net), .I1(n9211[3]), .I2(n405), .I3(n26816), 
            .O(n9199[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5047_6 (.CI(n26816), .I0(n9211[3]), .I1(n405), .CO(n26817));
    SB_LUT4 add_5047_5_lut (.I0(GND_net), .I1(n9211[2]), .I2(n332), .I3(n26815), 
            .O(n9199[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3563[12]), .I1(n257[12]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3538[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5047_5 (.CI(n26815), .I0(n9211[2]), .I1(n332), .CO(n26816));
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3563[11]), .I1(n257[11]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3538[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3563[10]), .I1(n257[10]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3538[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3563[9]), .I1(n257[9]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3538[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3563[8]), .I1(n257[8]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3538[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_4_lut (.I0(GND_net), .I1(n9211[1]), .I2(n259_adj_4252), 
            .I3(n26814), .O(n9199[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5047_4 (.CI(n26814), .I0(n9211[1]), .I1(n259_adj_4252), 
            .CO(n26815));
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3563[7]), .I1(n257[7]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_3_lut (.I0(GND_net), .I1(n9211[0]), .I2(n186_adj_4253), 
            .I3(n26813), .O(n9199[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3538[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3563[6]), .I1(n257[6]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3538[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3563[5]), .I1(n257[5]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3538[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3563[4]), .I1(n257[4]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5047_3 (.CI(n26813), .I0(n9211[0]), .I1(n186_adj_4253), 
            .CO(n26814));
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3538[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3563[3]), .I1(n257[3]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3538[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5047_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n9199[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5047_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5047_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n26813));
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4252));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28740_4_lut (.I0(n34735), .I1(n34867), .I2(n35_adj_4235), 
            .I3(n34201), .O(n34914));   // verilog/motorControl.v(36[10:25])
    defparam i28740_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4254));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5046_12_lut (.I0(GND_net), .I1(n9199[9]), .I2(n840), .I3(n26812), 
            .O(n9186[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5046_11_lut (.I0(GND_net), .I1(n9199[8]), .I2(n767), .I3(n26811), 
            .O(n9186[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_11 (.CI(n26811), .I0(n9199[8]), .I1(n767), .CO(n26812));
    SB_LUT4 i28741_3_lut (.I0(n34914), .I1(duty_23__N_3563[18]), .I2(n37), 
            .I3(GND_net), .O(n34915));   // verilog/motorControl.v(36[10:25])
    defparam i28741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4257));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4258));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5046_10_lut (.I0(GND_net), .I1(n9199[7]), .I2(n694), .I3(n26810), 
            .O(n9186[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4259));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4260));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5046_10 (.CI(n26810), .I0(n9199[7]), .I1(n694), .CO(n26811));
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4261));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[1]), 
            .I3(n25748), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4263));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4264));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3563[2]), .I1(n257[2]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3538[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5046_9_lut (.I0(GND_net), .I1(n9199[6]), .I2(n621), .I3(n26809), 
            .O(n9186[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4266));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5046_9 (.CI(n26809), .I0(n9199[6]), .I1(n621), .CO(n26810));
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4267));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4269));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4270));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5046_8_lut (.I0(GND_net), .I1(n9199[5]), .I2(n548), .I3(n26808), 
            .O(n9186[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28724_3_lut (.I0(n34915), .I1(duty_23__N_3563[19]), .I2(n39), 
            .I3(GND_net), .O(n34898));   // verilog/motorControl.v(36[10:25])
    defparam i28724_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5046_8 (.CI(n26808), .I0(n9199[5]), .I1(n548), .CO(n26809));
    SB_LUT4 add_5046_7_lut (.I0(GND_net), .I1(n9199[4]), .I2(n475), .I3(n26807), 
            .O(n9186[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4272));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4273));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28020_4_lut (.I0(n43), .I1(n41_adj_4274), .I2(n39), .I3(n34857), 
            .O(n34192));
    defparam i28020_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28642_4_lut (.I0(n34733), .I1(n34662), .I2(n45), .I3(n34190), 
            .O(n34816));   // verilog/motorControl.v(36[10:25])
    defparam i28642_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28710_3_lut (.I0(n34898), .I1(duty_23__N_3563[20]), .I2(n41_adj_4274), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i28710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4275));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4276));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4277));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28644_4_lut (.I0(n40), .I1(n34816), .I2(n45), .I3(n34192), 
            .O(n34818));   // verilog/motorControl.v(36[10:25])
    defparam i28644_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5046_7 (.CI(n26807), .I0(n9199[4]), .I1(n475), .CO(n26808));
    SB_LUT4 i28645_3_lut (.I0(n34818), .I1(PWMLimit[23]), .I2(duty_23__N_3563[23]), 
            .I3(GND_net), .O(duty_23__N_3562));   // verilog/motorControl.v(36[10:25])
    defparam i28645_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5046_6_lut (.I0(GND_net), .I1(n9199[3]), .I2(n402), .I3(n26806), 
            .O(n9186[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_6 (.CI(n26806), .I0(n9199[3]), .I1(n402), .CO(n26807));
    SB_LUT4 add_5046_5_lut (.I0(GND_net), .I1(n9199[2]), .I2(n329), .I3(n26805), 
            .O(n9186[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4278));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17816_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17816_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5046_5 (.CI(n26805), .I0(n9199[2]), .I1(n329), .CO(n26806));
    SB_LUT4 add_5046_4_lut (.I0(GND_net), .I1(n9199[1]), .I2(n256), .I3(n26804), 
            .O(n9186[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_4 (.CI(n26804), .I0(n9199[1]), .I1(n256), .CO(n26805));
    SB_LUT4 add_5046_3_lut (.I0(GND_net), .I1(n9199[0]), .I2(n183_adj_4240), 
            .I3(n26803), .O(n9186[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_3 (.CI(n26803), .I0(n9199[0]), .I1(n183_adj_4240), 
            .CO(n26804));
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4279));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5046_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n9186[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5046_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5046_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n26803));
    SB_LUT4 add_5045_13_lut (.I0(GND_net), .I1(n9186[10]), .I2(n910), 
            .I3(n26802), .O(n9172[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5045_12_lut (.I0(GND_net), .I1(n9186[9]), .I2(n837), .I3(n26801), 
            .O(n9172[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4281));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5045_12 (.CI(n26801), .I0(n9186[9]), .I1(n837), .CO(n26802));
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4282));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17817_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17817_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4284));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4285));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4286));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4287));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4289));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4290));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5045_11_lut (.I0(GND_net), .I1(n9186[8]), .I2(n764), .I3(n26800), 
            .O(n9172[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_11 (.CI(n26800), .I0(n9186[8]), .I1(n764), .CO(n26801));
    SB_LUT4 add_5045_10_lut (.I0(GND_net), .I1(n9186[7]), .I2(n691), .I3(n26799), 
            .O(n9172[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n25748), .I0(GND_net), .I1(n1_adj_4633[1]), 
            .CO(n25749));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3563[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_10 (.CI(n26799), .I0(n9186[7]), .I1(n691), .CO(n26800));
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4291));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4292));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5045_9_lut (.I0(GND_net), .I1(n9186[6]), .I2(n618), .I3(n26798), 
            .O(n9172[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4633[0]), 
            .CO(n25748));
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3563[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4294));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4295));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5045_9 (.CI(n26798), .I0(n9186[6]), .I1(n618), .CO(n26799));
    SB_LUT4 add_5045_8_lut (.I0(GND_net), .I1(n9186[5]), .I2(n545), .I3(n26797), 
            .O(n9172[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_8 (.CI(n26797), .I0(n9186[5]), .I1(n545), .CO(n26798));
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5045_7_lut (.I0(GND_net), .I1(n9186[4]), .I2(n472), .I3(n26796), 
            .O(n9172[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4632[23]), 
            .I3(n25747), .O(\PID_CONTROLLER.integral_23__N_3514 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n25614));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4300));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4301));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3563[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4303));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17818_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17818_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17819_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17819_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17820_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17820_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4306));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4307));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4309));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4310));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4312));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4313));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4315));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4316));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4318));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5045_7 (.CI(n26796), .I0(n9186[4]), .I1(n472), .CO(n26797));
    SB_LUT4 add_5045_6_lut (.I0(GND_net), .I1(n9186[3]), .I2(n399), .I3(n26795), 
            .O(n9172[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_6 (.CI(n26795), .I0(n9186[3]), .I1(n399), .CO(n26796));
    SB_LUT4 add_5045_5_lut (.I0(GND_net), .I1(n9186[2]), .I2(n326), .I3(n26794), 
            .O(n9172[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_5 (.CI(n26794), .I0(n9186[2]), .I1(n326), .CO(n26795));
    SB_LUT4 add_5045_4_lut (.I0(GND_net), .I1(n9186[1]), .I2(n253), .I3(n26793), 
            .O(n9172[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5045_4 (.CI(n26793), .I0(n9186[1]), .I1(n253), .CO(n26794));
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4632[22]), .I3(n25746), .O(n45_adj_4319)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5045_3_lut (.I0(GND_net), .I1(n9186[0]), .I2(n180), .I3(n26792), 
            .O(n9172[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17821_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17821_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n25746), .I0(GND_net), .I1(n1_adj_4632[22]), 
            .CO(n25747));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4632[21]), .I3(n25745), .O(n43_adj_4320)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4321));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4322));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4324));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4325));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4327));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5045_3 (.CI(n26792), .I0(n9186[0]), .I1(n180), .CO(n26793));
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4328));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3563[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4330));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5045_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n9172[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5045_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n25745), .I0(GND_net), .I1(n1_adj_4632[21]), 
            .CO(n25746));
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4214));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5045_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n26792));
    SB_LUT4 add_5044_14_lut (.I0(GND_net), .I1(n9172[11]), .I2(n980), 
            .I3(n26791), .O(n9157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4632[20]), .I3(n25744), .O(n41_adj_4331)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n25744), .I0(GND_net), .I1(n1_adj_4632[20]), 
            .CO(n25745));
    SB_LUT4 add_5044_13_lut (.I0(GND_net), .I1(n9172[10]), .I2(n907), 
            .I3(n26790), .O(n9157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_13 (.CI(n26790), .I0(n9172[10]), .I1(n907), .CO(n26791));
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3563[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4332));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4632[19]), .I3(n25743), .O(n39_adj_4333)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3563[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4334));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3563[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4335));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3563[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4336));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3563[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4337));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3563[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4338));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5044_12_lut (.I0(GND_net), .I1(n9172[9]), .I2(n834), .I3(n26789), 
            .O(n9157[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3563[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4339));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3563[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4340));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3563[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4341));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3563[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4342));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3563[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4343));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5044_12 (.CI(n26789), .I0(n9172[9]), .I1(n834), .CO(n26790));
    SB_LUT4 add_5044_11_lut (.I0(GND_net), .I1(n9172[8]), .I2(n761), .I3(n26788), 
            .O(n9157[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n25743), .I0(GND_net), .I1(n1_adj_4632[19]), 
            .CO(n25744));
    SB_CARRY add_5044_11 (.CI(n26788), .I0(n9172[8]), .I1(n761), .CO(n26789));
    SB_LUT4 i17822_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17822_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5044_10_lut (.I0(GND_net), .I1(n9172[7]), .I2(n688), .I3(n26787), 
            .O(n9157[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_10 (.CI(n26787), .I0(n9172[7]), .I1(n688), .CO(n26788));
    SB_LUT4 add_5044_9_lut (.I0(GND_net), .I1(n9172[6]), .I2(n615), .I3(n26786), 
            .O(n9157[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_9 (.CI(n26786), .I0(n9172[6]), .I1(n615), .CO(n26787));
    SB_LUT4 add_5044_8_lut (.I0(GND_net), .I1(n9172[5]), .I2(n542), .I3(n26785), 
            .O(n9157[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_8 (.CI(n26785), .I0(n9172[5]), .I1(n542), .CO(n26786));
    SB_LUT4 add_5044_7_lut (.I0(GND_net), .I1(n9172[4]), .I2(n469), .I3(n26784), 
            .O(n9157[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4632[18]), .I3(n25742), .O(n37_adj_4345)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5044_7 (.CI(n26784), .I0(n9172[4]), .I1(n469), .CO(n26785));
    SB_LUT4 add_5044_6_lut (.I0(GND_net), .I1(n9172[3]), .I2(n396), .I3(n26783), 
            .O(n9157[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_6 (.CI(n26783), .I0(n9172[3]), .I1(n396), .CO(n26784));
    SB_LUT4 add_5044_5_lut (.I0(GND_net), .I1(n9172[2]), .I2(n323), .I3(n26782), 
            .O(n9157[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_5 (.CI(n26782), .I0(n9172[2]), .I1(n323), .CO(n26783));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n25742), .I0(GND_net), .I1(n1_adj_4632[18]), 
            .CO(n25743));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4632[17]), .I3(n25741), .O(n35_adj_4346)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5044_4_lut (.I0(GND_net), .I1(n9172[1]), .I2(n250), .I3(n26781), 
            .O(n9157[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n25741), .I0(GND_net), .I1(n1_adj_4632[17]), 
            .CO(n25742));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4632[16]), .I3(n25740), .O(n33_adj_4347)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n25740), .I0(GND_net), .I1(n1_adj_4632[16]), 
            .CO(n25741));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4632[15]), .I3(n25739), .O(n31_adj_4348)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5044_4 (.CI(n26781), .I0(n9172[1]), .I1(n250), .CO(n26782));
    SB_LUT4 add_5044_3_lut (.I0(GND_net), .I1(n9172[0]), .I2(n177), .I3(n26780), 
            .O(n9157[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_3 (.CI(n26780), .I0(n9172[0]), .I1(n177), .CO(n26781));
    SB_LUT4 add_5044_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n9157[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5044_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5044_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n26780));
    SB_LUT4 add_5043_15_lut (.I0(GND_net), .I1(n9157[12]), .I2(n1050), 
            .I3(n26779), .O(n9141[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_14_lut (.I0(GND_net), .I1(n9157[11]), .I2(n977), 
            .I3(n26778), .O(n9141[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_14 (.CI(n26778), .I0(n9157[11]), .I1(n977), .CO(n26779));
    SB_LUT4 add_5043_13_lut (.I0(GND_net), .I1(n9157[10]), .I2(n904), 
            .I3(n26777), .O(n9141[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3563[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4349));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n25739), .I0(GND_net), .I1(n1_adj_4632[15]), 
            .CO(n25740));
    SB_CARRY add_5043_13 (.CI(n26777), .I0(n9157[10]), .I1(n904), .CO(n26778));
    SB_LUT4 add_5043_12_lut (.I0(GND_net), .I1(n9157[9]), .I2(n831_adj_4224), 
            .I3(n26776), .O(n9141[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_12 (.CI(n26776), .I0(n9157[9]), .I1(n831_adj_4224), 
            .CO(n26777));
    SB_LUT4 add_5043_11_lut (.I0(GND_net), .I1(n9157[8]), .I2(n758_adj_4223), 
            .I3(n26775), .O(n9141[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_11 (.CI(n26775), .I0(n9157[8]), .I1(n758_adj_4223), 
            .CO(n26776));
    SB_LUT4 add_5043_10_lut (.I0(GND_net), .I1(n9157[7]), .I2(n685_adj_4217), 
            .I3(n26774), .O(n9141[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4632[14]), .I3(n25738), .O(n29_adj_4350)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n25738), .I0(GND_net), .I1(n1_adj_4632[14]), 
            .CO(n25739));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4632[13]), .I3(n25737), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n25737), .I0(GND_net), .I1(n1_adj_4632[13]), 
            .CO(n25738));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4632[12]), .I3(n25736), .O(n25_adj_4351)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n25736), .I0(GND_net), .I1(n1_adj_4632[12]), 
            .CO(n25737));
    SB_CARRY add_5043_10 (.CI(n26774), .I0(n9157[7]), .I1(n685_adj_4217), 
            .CO(n26775));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4632[11]), .I3(n25735), .O(n23_adj_4352)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5043_9_lut (.I0(GND_net), .I1(n9157[6]), .I2(n612_adj_4216), 
            .I3(n26773), .O(n9141[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_9 (.CI(n26773), .I0(n9157[6]), .I1(n612_adj_4216), 
            .CO(n26774));
    SB_LUT4 add_5043_8_lut (.I0(GND_net), .I1(n9157[5]), .I2(n539), .I3(n26772), 
            .O(n9141[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_8 (.CI(n26772), .I0(n9157[5]), .I1(n539), .CO(n26773));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n25735), .I0(GND_net), .I1(n1_adj_4632[11]), 
            .CO(n25736));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4632[10]), .I3(n25734), .O(n21_adj_4353)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5043_7_lut (.I0(GND_net), .I1(n9157[4]), .I2(n466), .I3(n26771), 
            .O(n9141[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_7 (.CI(n26771), .I0(n9157[4]), .I1(n466), .CO(n26772));
    SB_LUT4 add_5043_6_lut (.I0(GND_net), .I1(n9157[3]), .I2(n393), .I3(n26770), 
            .O(n9141[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n25734), .I0(GND_net), .I1(n1_adj_4632[10]), 
            .CO(n25735));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4632[9]), .I3(n25733), .O(n19_adj_4354)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5043_6 (.CI(n26770), .I0(n9157[3]), .I1(n393), .CO(n26771));
    SB_LUT4 add_5043_5_lut (.I0(GND_net), .I1(n9157[2]), .I2(n320), .I3(n26769), 
            .O(n9141[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_5 (.CI(n26769), .I0(n9157[2]), .I1(n320), .CO(n26770));
    SB_LUT4 add_5043_4_lut (.I0(GND_net), .I1(n9157[1]), .I2(n247), .I3(n26768), 
            .O(n9141[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_4 (.CI(n26768), .I0(n9157[1]), .I1(n247), .CO(n26769));
    SB_LUT4 add_5043_3_lut (.I0(GND_net), .I1(n9157[0]), .I2(n174), .I3(n26767), 
            .O(n9141[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_3 (.CI(n26767), .I0(n9157[0]), .I1(n174), .CO(n26768));
    SB_LUT4 add_5043_2_lut (.I0(GND_net), .I1(n32_adj_4355), .I2(n101_adj_4356), 
            .I3(GND_net), .O(n9141[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_2 (.CI(GND_net), .I0(n32_adj_4355), .I1(n101_adj_4356), 
            .CO(n26767));
    SB_LUT4 add_5042_16_lut (.I0(GND_net), .I1(n9141[13]), .I2(n1120_adj_4357), 
            .I3(n26766), .O(n9124[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5042_15_lut (.I0(GND_net), .I1(n9141[12]), .I2(n1047_adj_4358), 
            .I3(n26765), .O(n9124[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_15 (.CI(n26765), .I0(n9141[12]), .I1(n1047_adj_4358), 
            .CO(n26766));
    SB_LUT4 add_5042_14_lut (.I0(GND_net), .I1(n9141[11]), .I2(n974_adj_4359), 
            .I3(n26764), .O(n9124[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_14 (.CI(n26764), .I0(n9141[11]), .I1(n974_adj_4359), 
            .CO(n26765));
    SB_LUT4 add_5042_13_lut (.I0(GND_net), .I1(n9141[10]), .I2(n901_adj_4360), 
            .I3(n26763), .O(n9124[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_13 (.CI(n26763), .I0(n9141[10]), .I1(n901_adj_4360), 
            .CO(n26764));
    SB_LUT4 add_5042_12_lut (.I0(GND_net), .I1(n9141[9]), .I2(n828_adj_4361), 
            .I3(n26762), .O(n9124[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_12 (.CI(n26762), .I0(n9141[9]), .I1(n828_adj_4361), 
            .CO(n26763));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n25733), .I0(GND_net), .I1(n1_adj_4632[9]), 
            .CO(n25734));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4632[8]), .I3(n25732), .O(n17_adj_4362)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5042_11_lut (.I0(GND_net), .I1(n9141[8]), .I2(n755_adj_4364), 
            .I3(n26761), .O(n9124[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n25732), .I0(GND_net), .I1(n1_adj_4632[8]), 
            .CO(n25733));
    SB_CARRY add_5042_11 (.CI(n26761), .I0(n9141[8]), .I1(n755_adj_4364), 
            .CO(n26762));
    SB_LUT4 add_5042_10_lut (.I0(GND_net), .I1(n9141[7]), .I2(n682_adj_4365), 
            .I3(n26760), .O(n9124[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4632[7]), .I3(n25731), .O(n15_adj_4366)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4368));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3563[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4369));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3563[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4370));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3563[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4371));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3563[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4372));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28004_4_lut (.I0(n21_adj_4343), .I1(n19_adj_4342), .I2(n17_adj_4341), 
            .I3(n9_adj_4340), .O(n34176));
    defparam i28004_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i27998_4_lut (.I0(n27_adj_4372), .I1(n15_adj_4371), .I2(n13_adj_4370), 
            .I3(n11_adj_4369), .O(n34170));
    defparam i27998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4349), 
            .I3(GND_net), .O(n12_adj_4373));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4370), 
            .I3(GND_net), .O(n10_adj_4374));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4373), .I1(n257[17]), .I2(n35_adj_4339), 
            .I3(GND_net), .O(n30_adj_4375));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4376));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4377));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17823_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17823_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28290_4_lut (.I0(n13_adj_4370), .I1(n11_adj_4369), .I2(n9_adj_4340), 
            .I3(n34186), .O(n34464));
    defparam i28290_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5042_10 (.CI(n26760), .I0(n9141[7]), .I1(n682_adj_4365), 
            .CO(n26761));
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4379));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4380));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5042_9_lut (.I0(GND_net), .I1(n9141[6]), .I2(n609_adj_4382), 
            .I3(n26759), .O(n9124[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_9 (.CI(n26759), .I0(n9141[6]), .I1(n609_adj_4382), 
            .CO(n26760));
    SB_LUT4 add_5042_8_lut (.I0(GND_net), .I1(n9141[5]), .I2(n536_adj_4383), 
            .I3(n26758), .O(n9124[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28286_4_lut (.I0(n19_adj_4342), .I1(n17_adj_4341), .I2(n15_adj_4371), 
            .I3(n34464), .O(n34460));
    defparam i28286_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i28624_4_lut (.I0(n25_adj_4338), .I1(n23_adj_4337), .I2(n21_adj_4343), 
            .I3(n34460), .O(n34798));
    defparam i28624_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28460_4_lut (.I0(n31_adj_4336), .I1(n29_adj_4335), .I2(n27_adj_4372), 
            .I3(n34798), .O(n34634));
    defparam i28460_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i28681_4_lut (.I0(n37_adj_4334), .I1(n35_adj_4339), .I2(n33_adj_4349), 
            .I3(n34634), .O(n34855));
    defparam i28681_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4332), 
            .I3(GND_net), .O(n16_adj_4385));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28606_3_lut (.I0(n6_adj_4386), .I1(n257[10]), .I2(n21_adj_4343), 
            .I3(GND_net), .O(n34780));   // verilog/motorControl.v(38[19:35])
    defparam i28606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28607_3_lut (.I0(n34780), .I1(n257[11]), .I2(n23_adj_4337), 
            .I3(GND_net), .O(n34781));   // verilog/motorControl.v(38[19:35])
    defparam i28607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4341), 
            .I3(GND_net), .O(n8_adj_4387));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4388));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5042_8 (.CI(n26758), .I0(n9141[5]), .I1(n536_adj_4383), 
            .CO(n26759));
    SB_LUT4 add_5042_7_lut (.I0(GND_net), .I1(n9141[4]), .I2(n463_adj_4389), 
            .I3(n26757), .O(n9124[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4390));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4391));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n25731), .I0(GND_net), .I1(n1_adj_4632[7]), 
            .CO(n25732));
    SB_CARRY add_5042_7 (.CI(n26757), .I0(n9141[4]), .I1(n463_adj_4389), 
            .CO(n26758));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4632[6]), .I3(n25730), .O(n13_adj_4392)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5042_6_lut (.I0(GND_net), .I1(n9141[3]), .I2(n390_adj_4394), 
            .I3(n26756), .O(n9124[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_6 (.CI(n26756), .I0(n9141[3]), .I1(n390_adj_4394), 
            .CO(n26757));
    SB_LUT4 i17824_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17824_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4395));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4397));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5042_5_lut (.I0(GND_net), .I1(n9141[2]), .I2(n317_adj_4398), 
            .I3(n26755), .O(n9124[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_5 (.CI(n26755), .I0(n9141[2]), .I1(n317_adj_4398), 
            .CO(n26756));
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_832_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3563[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3563[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4274));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3563[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3563[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3563[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4232));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3563[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3563[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3563[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4399));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3563[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4400));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3563[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4235));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3563[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3563[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4401));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3563[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4402));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3563[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4403));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3563[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4404));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3563[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4405));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3563[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4406));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4407));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4409));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4410));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17825_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17825_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5042_4_lut (.I0(GND_net), .I1(n9141[1]), .I2(n244_adj_4411), 
            .I3(n26754), .O(n9124[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n25730), .I0(GND_net), .I1(n1_adj_4632[6]), 
            .CO(n25731));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4632[5]), .I3(n25729), .O(n11_adj_4412)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n25729), .I0(GND_net), .I1(n1_adj_4632[5]), 
            .CO(n25730));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4632[4]), .I3(n25728), .O(n9_adj_4414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n25728), .I0(GND_net), .I1(n1_adj_4632[4]), 
            .CO(n25729));
    SB_LUT4 add_694_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3005[23]), .I3(n25677), .O(\PID_CONTROLLER.integral_23__N_3463 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_832_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3563[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4416));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_694_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3005[22]), .I3(n25676), .O(\PID_CONTROLLER.integral_23__N_3463 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_4 (.CI(n26754), .I0(n9141[1]), .I1(n244_adj_4411), 
            .CO(n26755));
    SB_LUT4 duty_23__I_832_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3563[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4417));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5042_3_lut (.I0(GND_net), .I1(n9141[0]), .I2(n171_adj_4418), 
            .I3(n26753), .O(n9124[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_3 (.CI(n26753), .I0(n9141[0]), .I1(n171_adj_4418), 
            .CO(n26754));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4632[3]), .I3(n25727), .O(n7_adj_4419)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_694_24 (.CI(n25676), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3005[22]), .CO(n25677));
    SB_LUT4 i28042_4_lut (.I0(n21_adj_4417), .I1(n19_adj_4416), .I2(n17_adj_4406), 
            .I3(n9_adj_4405), .O(n34214));
    defparam i28042_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3563[1]), .I1(n257[1]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3538[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n25727), .I0(GND_net), .I1(n1_adj_4632[3]), 
            .CO(n25728));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4632[2]), .I3(n25726), .O(n5_adj_4421)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_694_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3005[21]), .I3(n25675), .O(\PID_CONTROLLER.integral_23__N_3463 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_23 (.CI(n25675), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3005[21]), .CO(n25676));
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n7405[0]), .I2(n7409[0]), 
            .I3(n25636), .O(duty_23__N_3563[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4385), .I1(n257[22]), .I2(n45_adj_4330), 
            .I3(GND_net), .O(n24_adj_4423));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5042_2_lut (.I0(GND_net), .I1(n29_adj_4424), .I2(n98_adj_4425), 
            .I3(GND_net), .O(n9124[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5042_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n25635), .O(duty_23__N_3563[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5042_2 (.CI(GND_net), .I0(n29_adj_4424), .I1(n98_adj_4425), 
            .CO(n26753));
    SB_LUT4 i28035_4_lut (.I0(n27_adj_4404), .I1(n15_adj_4403), .I2(n13_adj_4402), 
            .I3(n11_adj_4401), .O(n34207));
    defparam i28035_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5041_17_lut (.I0(GND_net), .I1(n9124[14]), .I2(GND_net), 
            .I3(n26752), .O(n9106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_832_i12_3_lut (.I0(duty_23__N_3563[7]), .I1(duty_23__N_3563[16]), 
            .I2(n33), .I3(GND_net), .O(n12_adj_4426));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5041_16_lut (.I0(GND_net), .I1(n9124[13]), .I2(n1117_adj_4427), 
            .I3(n26751), .O(n9106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_16 (.CI(n26751), .I0(n9124[13]), .I1(n1117_adj_4427), 
            .CO(n26752));
    SB_LUT4 add_694_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3005[20]), .I3(n25674), .O(\PID_CONTROLLER.integral_23__N_3463 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_15_lut (.I0(GND_net), .I1(n9124[12]), .I2(n1044_adj_4428), 
            .I3(n26750), .O(n9106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4429));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4430));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_15 (.CI(n26750), .I0(n9124[12]), .I1(n1044_adj_4428), 
            .CO(n26751));
    SB_LUT4 add_5041_14_lut (.I0(GND_net), .I1(n9124[11]), .I2(n971_adj_4431), 
            .I3(n26749), .O(n9106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_14 (.CI(n26749), .I0(n9124[11]), .I1(n971_adj_4431), 
            .CO(n26750));
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4432));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_24 (.CI(n25635), .I0(n106[22]), .I1(n155[22]), .CO(n25636));
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4433));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n25634), .O(duty_23__N_3563[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n25634), .I0(n106[21]), .I1(n155[21]), .CO(n25635));
    SB_LUT4 add_5041_13_lut (.I0(GND_net), .I1(n9124[10]), .I2(n898_adj_4434), 
            .I3(n26748), .O(n9106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_13 (.CI(n26748), .I0(n9124[10]), .I1(n898_adj_4434), 
            .CO(n26749));
    SB_LUT4 add_5041_12_lut (.I0(GND_net), .I1(n9124[9]), .I2(n825_adj_4435), 
            .I3(n26747), .O(n9106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4436));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4437));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4438));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_12 (.CI(n26747), .I0(n9124[9]), .I1(n825_adj_4435), 
            .CO(n26748));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n25726), .I0(GND_net), .I1(n1_adj_4632[2]), 
            .CO(n25727));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5041_11_lut (.I0(GND_net), .I1(n9124[8]), .I2(n752_adj_4440), 
            .I3(n26746), .O(n9106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4441));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_694_22 (.CI(n25674), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3005[20]), .CO(n25675));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n25633), .O(duty_23__N_3563[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4632[1]), .I3(n25725), .O(n3_adj_4443)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n25725), .I0(GND_net), .I1(n1_adj_4632[1]), 
            .CO(n25726));
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4446));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4447));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4632[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3514 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4632[0]), 
            .CO(n25725));
    SB_CARRY add_5041_11 (.CI(n26746), .I0(n9124[8]), .I1(n752_adj_4440), 
            .CO(n26747));
    SB_LUT4 add_694_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3005[19]), .I3(n25673), .O(\PID_CONTROLLER.integral_23__N_3463 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_21 (.CI(n25673), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3005[19]), .CO(n25674));
    SB_LUT4 add_694_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3005[18]), .I3(n25672), .O(\PID_CONTROLLER.integral_23__N_3463 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n25633), .I0(n106[20]), .I1(n155[20]), .CO(n25634));
    SB_CARRY add_694_20 (.CI(n25672), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3005[18]), .CO(n25673));
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n25632), .O(duty_23__N_3563[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n25632), .I0(n106[19]), .I1(n155[19]), .CO(n25633));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n25724), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4452));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_694_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3005[17]), .I3(n25671), .O(\PID_CONTROLLER.integral_23__N_3463 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_19 (.CI(n25671), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3005[17]), .CO(n25672));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n25631), .O(duty_23__N_3563[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n25723), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5041_10_lut (.I0(GND_net), .I1(n9124[7]), .I2(n679_adj_4454), 
            .I3(n26745), .O(n9106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n25723), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n25724));
    SB_LUT4 add_694_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3005[16]), .I3(n25670), .O(\PID_CONTROLLER.integral_23__N_3463 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_18 (.CI(n25670), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3005[16]), .CO(n25671));
    SB_LUT4 i27984_4_lut (.I0(n43_adj_4332), .I1(n25_adj_4338), .I2(n23_adj_4337), 
            .I3(n34176), .O(n34156));
    defparam i27984_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28490_4_lut (.I0(n24_adj_4423), .I1(n8_adj_4387), .I2(n45_adj_4330), 
            .I3(n34154), .O(n34664));   // verilog/motorControl.v(38[19:35])
    defparam i28490_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28565_3_lut (.I0(n34781), .I1(n257[12]), .I2(n25_adj_4338), 
            .I3(GND_net), .O(n34739));   // verilog/motorControl.v(38[19:35])
    defparam i28565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3563[0]), .I1(n257[1]), 
            .I2(duty_23__N_3563[1]), .I3(n257[0]), .O(n4_adj_4455));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i28604_3_lut (.I0(n4_adj_4455), .I1(n257[13]), .I2(n27_adj_4372), 
            .I3(GND_net), .O(n34778));   // verilog/motorControl.v(38[19:35])
    defparam i28604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28605_3_lut (.I0(n34778), .I1(n257[14]), .I2(n29_adj_4335), 
            .I3(GND_net), .O(n34779));   // verilog/motorControl.v(38[19:35])
    defparam i28605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27994_4_lut (.I0(n33_adj_4349), .I1(n31_adj_4336), .I2(n29_adj_4335), 
            .I3(n34170), .O(n34166));
    defparam i27994_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28695_4_lut (.I0(n30_adj_4375), .I1(n10_adj_4374), .I2(n35_adj_4339), 
            .I3(n34164), .O(n34869));   // verilog/motorControl.v(38[19:35])
    defparam i28695_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28567_3_lut (.I0(n34779), .I1(n257[15]), .I2(n31_adj_4336), 
            .I3(GND_net), .O(n34741));   // verilog/motorControl.v(38[19:35])
    defparam i28567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28742_4_lut (.I0(n34741), .I1(n34869), .I2(n35_adj_4339), 
            .I3(n34166), .O(n34916));   // verilog/motorControl.v(38[19:35])
    defparam i28742_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28743_3_lut (.I0(n34916), .I1(n257[18]), .I2(n37_adj_4334), 
            .I3(GND_net), .O(n34917));   // verilog/motorControl.v(38[19:35])
    defparam i28743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28722_3_lut (.I0(n34917), .I1(n257[19]), .I2(n39_adj_4303), 
            .I3(GND_net), .O(n34896));   // verilog/motorControl.v(38[19:35])
    defparam i28722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27986_4_lut (.I0(n43_adj_4332), .I1(n41_adj_4294), .I2(n39_adj_4303), 
            .I3(n34855), .O(n34158));
    defparam i27986_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28648_4_lut (.I0(n34739), .I1(n34664), .I2(n45_adj_4330), 
            .I3(n34156), .O(n34822));   // verilog/motorControl.v(38[19:35])
    defparam i28648_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28712_3_lut (.I0(n34896), .I1(n257[20]), .I2(n41_adj_4294), 
            .I3(GND_net), .O(n40_adj_4456));   // verilog/motorControl.v(38[19:35])
    defparam i28712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28650_4_lut (.I0(n40_adj_4456), .I1(n34822), .I2(n45_adj_4330), 
            .I3(n34158), .O(n34824));   // verilog/motorControl.v(38[19:35])
    defparam i28650_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28651_3_lut (.I0(n34824), .I1(duty_23__N_3563[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4245));   // verilog/motorControl.v(38[19:35])
    defparam i28651_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3563[0]), .I1(n257[0]), .I2(n256_adj_4245), 
            .I3(GND_net), .O(duty_23__N_3538[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3538[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3562), .I3(GND_net), .O(duty_23__N_3439[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_10 (.CI(n26745), .I0(n9124[7]), .I1(n679_adj_4454), 
            .CO(n26746));
    SB_LUT4 add_5041_9_lut (.I0(GND_net), .I1(n9124[6]), .I2(n606_adj_4457), 
            .I3(n26744), .O(n9106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_9 (.CI(n26744), .I0(n9124[6]), .I1(n606_adj_4457), 
            .CO(n26745));
    SB_LUT4 add_5041_8_lut (.I0(GND_net), .I1(n9124[5]), .I2(n533_adj_4458), 
            .I3(n26743), .O(n9106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_8 (.CI(n26743), .I0(n9124[5]), .I1(n533_adj_4458), 
            .CO(n26744));
    SB_LUT4 add_5041_7_lut (.I0(GND_net), .I1(n9124[4]), .I2(n460_adj_4459), 
            .I3(n26742), .O(n9106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28055_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3563[3]), 
            .I2(duty_23__N_3563[2]), .I3(PWMLimit[2]), .O(n34227));   // verilog/motorControl.v(36[10:25])
    defparam i28055_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_832_i10_3_lut (.I0(duty_23__N_3563[5]), .I1(duty_23__N_3563[6]), 
            .I2(n13_adj_4402), .I3(GND_net), .O(n10_adj_4234));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3563[3]), 
            .I2(duty_23__N_3563[2]), .I3(GND_net), .O(n6_adj_4460));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_5041_7 (.CI(n26742), .I0(n9124[4]), .I1(n460_adj_4459), 
            .CO(n26743));
    SB_LUT4 add_5041_6_lut (.I0(GND_net), .I1(n9124[3]), .I2(n387_adj_4461), 
            .I3(n26741), .O(n9106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4462));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_6 (.CI(n26741), .I0(n9124[3]), .I1(n387_adj_4461), 
            .CO(n26742));
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5041_5_lut (.I0(GND_net), .I1(n9124[2]), .I2(n314_adj_4464), 
            .I3(n26740), .O(n9106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4465));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4467));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4468));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17826_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17826_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4470));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17827_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17827_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4471));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17828_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17828_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5041_5 (.CI(n26740), .I0(n9124[2]), .I1(n314_adj_4464), 
            .CO(n26741));
    SB_LUT4 add_5041_4_lut (.I0(GND_net), .I1(n9124[1]), .I2(n241_adj_4473), 
            .I3(n26739), .O(n9106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_4 (.CI(n26739), .I0(n9124[1]), .I1(n241_adj_4473), 
            .CO(n26740));
    SB_LUT4 add_5041_3_lut (.I0(GND_net), .I1(n9124[0]), .I2(n168_adj_4474), 
            .I3(n26738), .O(n9106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_3 (.CI(n26738), .I0(n9124[0]), .I1(n168_adj_4474), 
            .CO(n26739));
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5041_2_lut (.I0(GND_net), .I1(n26_adj_4476), .I2(n95_adj_4477), 
            .I3(GND_net), .O(n9106[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5041_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5041_2 (.CI(GND_net), .I0(n26_adj_4476), .I1(n95_adj_4477), 
            .CO(n26738));
    SB_LUT4 add_5040_18_lut (.I0(GND_net), .I1(n9106[15]), .I2(GND_net), 
            .I3(n26737), .O(n9087[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_17_lut (.I0(GND_net), .I1(n9106[14]), .I2(GND_net), 
            .I3(n26736), .O(n9087[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_17 (.CI(n26736), .I0(n9106[14]), .I1(GND_net), .CO(n26737));
    SB_LUT4 add_5040_16_lut (.I0(GND_net), .I1(n9106[13]), .I2(n1114_adj_4478), 
            .I3(n26735), .O(n9087[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_16 (.CI(n26735), .I0(n9106[13]), .I1(n1114_adj_4478), 
            .CO(n26736));
    SB_LUT4 add_5040_15_lut (.I0(GND_net), .I1(n9106[12]), .I2(n1041_adj_4479), 
            .I3(n26734), .O(n9087[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4480));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17829_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17829_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4483));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4213));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4212));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4211));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5040_15 (.CI(n26734), .I0(n9106[12]), .I1(n1041_adj_4479), 
            .CO(n26735));
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5040_14_lut (.I0(GND_net), .I1(n9106[11]), .I2(n968_adj_4483), 
            .I3(n26733), .O(n9087[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_14 (.CI(n26733), .I0(n9106[11]), .I1(n968_adj_4483), 
            .CO(n26734));
    SB_CARRY add_12_20 (.CI(n25631), .I0(n106[18]), .I1(n155[18]), .CO(n25632));
    SB_LUT4 add_694_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3005[15]), .I3(n25669), .O(\PID_CONTROLLER.integral_23__N_3463 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_13_lut (.I0(GND_net), .I1(n9106[10]), .I2(n895_adj_4481), 
            .I3(n26732), .O(n9087[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_832_i30_3_lut (.I0(n12_adj_4426), .I1(duty_23__N_3563[17]), 
            .I2(n35_adj_4235), .I3(GND_net), .O(n30));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n25630), .O(duty_23__N_3563[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_13 (.CI(n26732), .I0(n9106[10]), .I1(n895_adj_4481), 
            .CO(n26733));
    SB_LUT4 add_5040_12_lut (.I0(GND_net), .I1(n9106[9]), .I2(n822_adj_4480), 
            .I3(n26731), .O(n9087[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_12 (.CI(n26731), .I0(n9106[9]), .I1(n822_adj_4480), 
            .CO(n26732));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n25722), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_11_lut (.I0(GND_net), .I1(n9106[8]), .I2(n749_adj_4475), 
            .I3(n26730), .O(n9087[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_17 (.CI(n25669), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3005[15]), .CO(n25670));
    SB_CARRY add_5040_11 (.CI(n26730), .I0(n9106[8]), .I1(n749_adj_4475), 
            .CO(n26731));
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4479));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5040_10_lut (.I0(GND_net), .I1(n9106[7]), .I2(n676_adj_4472), 
            .I3(n26729), .O(n9087[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n25630), .I0(n106[17]), .I1(n155[17]), .CO(n25631));
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_23 (.CI(n25722), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n25723));
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4477));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4476));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5040_10 (.CI(n26729), .I0(n9106[7]), .I1(n676_adj_4472), 
            .CO(n26730));
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n25629), .O(duty_23__N_3563[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4474));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4473));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_694_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3005[14]), .I3(n25668), .O(\PID_CONTROLLER.integral_23__N_3463 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4464));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_18 (.CI(n25629), .I0(n106[16]), .I1(n155[16]), .CO(n25630));
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4461));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4459));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4458));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_694_16 (.CI(n25668), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3005[14]), .CO(n25669));
    SB_LUT4 add_5040_9_lut (.I0(GND_net), .I1(n9106[6]), .I2(n603_adj_4471), 
            .I3(n26728), .O(n9087[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17830_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17830_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_694_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3005[13]), .I3(n25667), .O(\PID_CONTROLLER.integral_23__N_3463 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_9 (.CI(n26728), .I0(n9106[6]), .I1(n603_adj_4471), 
            .CO(n26729));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n25721), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_15 (.CI(n25667), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3005[13]), .CO(n25668));
    SB_LUT4 add_5040_8_lut (.I0(GND_net), .I1(n9106[5]), .I2(n530_adj_4470), 
            .I3(n26727), .O(n9087[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_8 (.CI(n26727), .I0(n9106[5]), .I1(n530_adj_4470), 
            .CO(n26728));
    SB_LUT4 add_5040_7_lut (.I0(GND_net), .I1(n9106[4]), .I2(n457_adj_4469), 
            .I3(n26726), .O(n9087[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_7 (.CI(n26726), .I0(n9106[4]), .I1(n457_adj_4469), 
            .CO(n26727));
    SB_LUT4 add_694_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3005[12]), .I3(n25666), .O(\PID_CONTROLLER.integral_23__N_3463 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_6_lut (.I0(GND_net), .I1(n9106[3]), .I2(n384_adj_4468), 
            .I3(n26725), .O(n9087[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_6 (.CI(n26725), .I0(n9106[3]), .I1(n384_adj_4468), 
            .CO(n26726));
    SB_LUT4 add_5040_5_lut (.I0(GND_net), .I1(n9106[2]), .I2(n311_adj_4467), 
            .I3(n26724), .O(n9087[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_5 (.CI(n26724), .I0(n9106[2]), .I1(n311_adj_4467), 
            .CO(n26725));
    SB_LUT4 add_5040_4_lut (.I0(GND_net), .I1(n9106[1]), .I2(n238_adj_4466), 
            .I3(n26723), .O(n9087[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n25721), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n25722));
    SB_CARRY add_5040_4 (.CI(n26723), .I0(n9106[1]), .I1(n238_adj_4466), 
            .CO(n26724));
    SB_LUT4 add_5040_3_lut (.I0(GND_net), .I1(n9106[0]), .I2(n165_adj_4465), 
            .I3(n26722), .O(n9087[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_3 (.CI(n26722), .I0(n9106[0]), .I1(n165_adj_4465), 
            .CO(n26723));
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n25720), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_2_lut (.I0(GND_net), .I1(n23_adj_4463), .I2(n92_adj_4462), 
            .I3(GND_net), .O(n9087[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n25720), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n25721));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5040_2 (.CI(GND_net), .I0(n23_adj_4463), .I1(n92_adj_4462), 
            .CO(n26722));
    SB_LUT4 add_5039_19_lut (.I0(GND_net), .I1(n9087[16]), .I2(GND_net), 
            .I3(n26721), .O(n9067[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_14 (.CI(n25666), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3005[12]), .CO(n25667));
    SB_LUT4 add_5039_18_lut (.I0(GND_net), .I1(n9087[15]), .I2(GND_net), 
            .I3(n26720), .O(n9067[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_18 (.CI(n26720), .I0(n9087[15]), .I1(GND_net), .CO(n26721));
    SB_LUT4 add_5039_17_lut (.I0(GND_net), .I1(n9087[14]), .I2(GND_net), 
            .I3(n26719), .O(n9067[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_17 (.CI(n26719), .I0(n9087[14]), .I1(GND_net), .CO(n26720));
    SB_LUT4 add_5039_16_lut (.I0(GND_net), .I1(n9087[13]), .I2(n1111_adj_4452), 
            .I3(n26718), .O(n9067[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_16 (.CI(n26718), .I0(n9087[13]), .I1(n1111_adj_4452), 
            .CO(n26719));
    SB_LUT4 add_5039_15_lut (.I0(GND_net), .I1(n9087[12]), .I2(n1038_adj_4451), 
            .I3(n26717), .O(n9067[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n25719), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_15 (.CI(n26717), .I0(n9087[12]), .I1(n1038_adj_4451), 
            .CO(n26718));
    SB_LUT4 add_5039_14_lut (.I0(GND_net), .I1(n9087[11]), .I2(n965_adj_4448), 
            .I3(n26716), .O(n9067[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_14 (.CI(n26716), .I0(n9087[11]), .I1(n965_adj_4448), 
            .CO(n26717));
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_13_lut (.I0(GND_net), .I1(n9087[10]), .I2(n892_adj_4447), 
            .I3(n26715), .O(n9067[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_13 (.CI(n26715), .I0(n9087[10]), .I1(n892_adj_4447), 
            .CO(n26716));
    SB_CARRY sub_3_add_2_20 (.CI(n25719), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n25720));
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_12_lut (.I0(GND_net), .I1(n9087[9]), .I2(n819_adj_4446), 
            .I3(n26714), .O(n9067[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_12 (.CI(n26714), .I0(n9087[9]), .I1(n819_adj_4446), 
            .CO(n26715));
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n25628), .O(duty_23__N_3563[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_11_lut (.I0(GND_net), .I1(n9087[8]), .I2(n746_adj_4445), 
            .I3(n26713), .O(n9067[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4233));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_11 (.CI(n26713), .I0(n9087[8]), .I1(n746_adj_4445), 
            .CO(n26714));
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_10_lut (.I0(GND_net), .I1(n9087[7]), .I2(n673_adj_4442), 
            .I3(n26712), .O(n9067[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_10 (.CI(n26712), .I0(n9087[7]), .I1(n673_adj_4442), 
            .CO(n26713));
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_9_lut (.I0(GND_net), .I1(n9087[6]), .I2(n600_adj_4441), 
            .I3(n26711), .O(n9067[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_9 (.CI(n26711), .I0(n9087[6]), .I1(n600_adj_4441), 
            .CO(n26712));
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4231));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_8_lut (.I0(GND_net), .I1(n9087[5]), .I2(n527_adj_4439), 
            .I3(n26710), .O(n9067[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_8 (.CI(n26710), .I0(n9087[5]), .I1(n527_adj_4439), 
            .CO(n26711));
    SB_LUT4 add_5039_7_lut (.I0(GND_net), .I1(n9087[4]), .I2(n454_adj_4438), 
            .I3(n26709), .O(n9067[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29253_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n35425));   // verilog/motorControl.v(29[14] 48[8])
    defparam i29253_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_7 (.CI(n26709), .I0(n9087[4]), .I1(n454_adj_4438), 
            .CO(n26710));
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_6_lut (.I0(GND_net), .I1(n9087[3]), .I2(n381_adj_4437), 
            .I3(n26708), .O(n9067[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_6 (.CI(n26708), .I0(n9087[3]), .I1(n381_adj_4437), 
            .CO(n26709));
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5039_5_lut (.I0(GND_net), .I1(n9087[2]), .I2(n308_adj_4436), 
            .I3(n26707), .O(n9067[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_5 (.CI(n26707), .I0(n9087[2]), .I1(n308_adj_4436), 
            .CO(n26708));
    SB_LUT4 add_5039_4_lut (.I0(GND_net), .I1(n9087[1]), .I2(n235_adj_4433), 
            .I3(n26706), .O(n9067[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_4 (.CI(n26706), .I0(n9087[1]), .I1(n235_adj_4433), 
            .CO(n26707));
    SB_LUT4 add_5039_3_lut (.I0(GND_net), .I1(n9087[0]), .I2(n162_adj_4432), 
            .I3(n26705), .O(n9067[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4222));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5039_3 (.CI(n26705), .I0(n9087[0]), .I1(n162_adj_4432), 
            .CO(n26706));
    SB_LUT4 i2_4_lut (.I0(n6_adj_4491), .I1(\Kp[4] ), .I2(n9256[2]), .I3(n1[18]), 
            .O(n9249[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 add_5039_2_lut (.I0(GND_net), .I1(n20_adj_4430), .I2(n89_adj_4429), 
            .I3(GND_net), .O(n9067[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5039_2 (.CI(GND_net), .I0(n20_adj_4430), .I1(n89_adj_4429), 
            .CO(n26705));
    SB_LUT4 add_5038_20_lut (.I0(GND_net), .I1(n9067[17]), .I2(GND_net), 
            .I3(n26704), .O(n9046[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5038_19_lut (.I0(GND_net), .I1(n9067[16]), .I2(GND_net), 
            .I3(n26703), .O(n9046[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_19 (.CI(n26703), .I0(n9067[16]), .I1(GND_net), .CO(n26704));
    SB_LUT4 add_5038_18_lut (.I0(GND_net), .I1(n9067[15]), .I2(GND_net), 
            .I3(n26702), .O(n9046[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3439[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5038_18 (.CI(n26702), .I0(n9067[15]), .I1(GND_net), .CO(n26703));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n25718), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_694_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3005[11]), .I3(n25665), .O(\PID_CONTROLLER.integral_23__N_3463 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20790_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n9267[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20790_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1478 (.I0(n4_adj_4492), .I1(\Kp[3] ), .I2(n9262[1]), 
            .I3(n1[19]), .O(n9256[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1478.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1479 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4493));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1479.LUT_INIT = 16'h9c50;
    SB_LUT4 i20726_4_lut (.I0(n9256[2]), .I1(\Kp[4] ), .I2(n6_adj_4491), 
            .I3(n1[18]), .O(n8_adj_4494));   // verilog/motorControl.v(34[16:22])
    defparam i20726_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), .I3(n1[21]), 
            .O(n11_adj_4495));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i17831_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17831_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5038_17_lut (.I0(GND_net), .I1(n9067[14]), .I2(GND_net), 
            .I3(n26701), .O(n9046[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20757_4_lut (.I0(n9262[1]), .I1(\Kp[3] ), .I2(n4_adj_4492), 
            .I3(n1[19]), .O(n6_adj_4496));   // verilog/motorControl.v(34[16:22])
    defparam i20757_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i20792_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n25357));   // verilog/motorControl.v(34[16:22])
    defparam i20792_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4496), .I1(n11_adj_4495), .I2(n8_adj_4494), 
            .I3(n12_adj_4493), .O(n18_adj_4497));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), .I3(n1[22]), 
            .O(n13_adj_4498));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_12_17 (.CI(n25628), .I0(n106[15]), .I1(n155[15]), .CO(n25629));
    SB_LUT4 i28014_3_lut_4_lut (.I0(duty_23__N_3563[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3563[2]), .O(n34186));   // verilog/motorControl.v(38[19:35])
    defparam i28014_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY sub_3_add_2_19 (.CI(n25718), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n25719));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n25717), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_17 (.CI(n26701), .I0(n9067[14]), .I1(GND_net), .CO(n26702));
    SB_LUT4 i28344_4_lut (.I0(n13_adj_4402), .I1(n11_adj_4401), .I2(n9_adj_4405), 
            .I3(n34227), .O(n34518));
    defparam i28344_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_5038_16_lut (.I0(GND_net), .I1(n9067[13]), .I2(n1108_adj_4410), 
            .I3(n26700), .O(n9046[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4498), .I1(n18_adj_4497), .I2(n25357), 
            .I3(n4_adj_4499), .O(n32507));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3563[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4386));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5038_16 (.CI(n26700), .I0(n9067[13]), .I1(n1108_adj_4410), 
            .CO(n26701));
    SB_LUT4 add_5038_15_lut (.I0(GND_net), .I1(n9067[12]), .I2(n1035_adj_4409), 
            .I3(n26699), .O(n9046[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_15 (.CI(n26699), .I0(n9067[12]), .I1(n1035_adj_4409), 
            .CO(n26700));
    SB_LUT4 add_5038_14_lut (.I0(GND_net), .I1(n9067[11]), .I2(n962_adj_4407), 
            .I3(n26698), .O(n9046[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_14 (.CI(n26698), .I0(n9067[11]), .I1(n962_adj_4407), 
            .CO(n26699));
    SB_CARRY add_694_13 (.CI(n25665), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3005[11]), .CO(n25666));
    SB_LUT4 add_5038_13_lut (.I0(GND_net), .I1(n9067[10]), .I2(n889_adj_4397), 
            .I3(n26697), .O(n9046[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_13 (.CI(n26697), .I0(n9067[10]), .I1(n889_adj_4397), 
            .CO(n26698));
    SB_LUT4 add_5038_12_lut (.I0(GND_net), .I1(n9067[9]), .I2(n816_adj_4396), 
            .I3(n26696), .O(n9046[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_12 (.CI(n26696), .I0(n9067[9]), .I1(n816_adj_4396), 
            .CO(n26697));
    SB_LUT4 add_5038_11_lut (.I0(GND_net), .I1(n9067[8]), .I2(n743_adj_4395), 
            .I3(n26695), .O(n9046[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n25717), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n25718));
    SB_CARRY add_5038_11 (.CI(n26695), .I0(n9067[8]), .I1(n743_adj_4395), 
            .CO(n26696));
    SB_LUT4 add_694_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3005[10]), .I3(n25664), .O(\PID_CONTROLLER.integral_23__N_3463 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n25716), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5038_10_lut (.I0(GND_net), .I1(n9067[7]), .I2(n670_adj_4391), 
            .I3(n26694), .O(n9046[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n25627), .O(duty_23__N_3563[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_10 (.CI(n26694), .I0(n9067[7]), .I1(n670_adj_4391), 
            .CO(n26695));
    SB_LUT4 i17832_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17832_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17833_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17833_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_17 (.CI(n25716), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n25717));
    SB_LUT4 add_5038_9_lut (.I0(GND_net), .I1(n9067[6]), .I2(n597_adj_4390), 
            .I3(n26693), .O(n9046[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5038_9 (.CI(n26693), .I0(n9067[6]), .I1(n597_adj_4390), 
            .CO(n26694));
    SB_LUT4 add_5038_8_lut (.I0(GND_net), .I1(n9067[5]), .I2(n524_adj_4388), 
            .I3(n26692), .O(n9046[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_8 (.CI(n26692), .I0(n9067[5]), .I1(n524_adj_4388), 
            .CO(n26693));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n25715), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4221));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_16 (.CI(n25715), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n25716));
    SB_LUT4 add_5038_7_lut (.I0(GND_net), .I1(n9067[4]), .I2(n451_adj_4384), 
            .I3(n26691), .O(n9046[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_7 (.CI(n26691), .I0(n9067[4]), .I1(n451_adj_4384), 
            .CO(n26692));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n25714), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4440));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_15 (.CI(n25714), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n25715));
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4435));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4434));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5038_6_lut (.I0(GND_net), .I1(n9067[3]), .I2(n378_adj_4381), 
            .I3(n26690), .O(n9046[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_6 (.CI(n26690), .I0(n9067[3]), .I1(n378_adj_4381), 
            .CO(n26691));
    SB_LUT4 add_5038_5_lut (.I0(GND_net), .I1(n9067[2]), .I2(n305_adj_4380), 
            .I3(n26689), .O(n9046[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_5 (.CI(n26689), .I0(n9067[2]), .I1(n305_adj_4380), 
            .CO(n26690));
    SB_LUT4 add_5038_4_lut (.I0(GND_net), .I1(n9067[1]), .I2(n232_adj_4379), 
            .I3(n26688), .O(n9046[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_4 (.CI(n26688), .I0(n9067[1]), .I1(n232_adj_4379), 
            .CO(n26689));
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4220));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4431));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5038_3_lut (.I0(GND_net), .I1(n9067[0]), .I2(n159_adj_4378), 
            .I3(n26687), .O(n9046[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n25713), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4428));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_14 (.CI(n25713), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n25714));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n25712), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_12 (.CI(n25664), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3005[10]), .CO(n25665));
    SB_CARRY add_5038_3 (.CI(n26687), .I0(n9067[0]), .I1(n159_adj_4378), 
            .CO(n26688));
    SB_CARRY add_12_16 (.CI(n25627), .I0(n106[14]), .I1(n155[14]), .CO(n25628));
    SB_CARRY sub_3_add_2_13 (.CI(n25712), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n25713));
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4219));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17834_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17834_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4427));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_694_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3005[9]), .I3(n25663), .O(\PID_CONTROLLER.integral_23__N_3463 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5038_2_lut (.I0(GND_net), .I1(n17_adj_4377), .I2(n86_adj_4376), 
            .I3(GND_net), .O(n9046[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5038_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5038_2 (.CI(GND_net), .I0(n17_adj_4377), .I1(n86_adj_4376), 
            .CO(n26687));
    SB_LUT4 add_5037_21_lut (.I0(GND_net), .I1(n9046[18]), .I2(GND_net), 
            .I3(n26686), .O(n9024[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_20_lut (.I0(GND_net), .I1(n9046[17]), .I2(GND_net), 
            .I3(n26685), .O(n9024[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_20 (.CI(n26685), .I0(n9046[17]), .I1(GND_net), .CO(n26686));
    SB_LUT4 add_5037_19_lut (.I0(GND_net), .I1(n9046[16]), .I2(GND_net), 
            .I3(n26684), .O(n9024[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_19 (.CI(n26684), .I0(n9046[16]), .I1(GND_net), .CO(n26685));
    SB_LUT4 add_5037_18_lut (.I0(GND_net), .I1(n9046[15]), .I2(GND_net), 
            .I3(n26683), .O(n9024[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_18 (.CI(n26683), .I0(n9046[15]), .I1(GND_net), .CO(n26684));
    SB_LUT4 add_5037_17_lut (.I0(GND_net), .I1(n9046[14]), .I2(GND_net), 
            .I3(n26682), .O(n9024[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_17 (.CI(n26682), .I0(n9046[14]), .I1(GND_net), .CO(n26683));
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4425));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5037_16_lut (.I0(GND_net), .I1(n9046[13]), .I2(n1105_adj_4368), 
            .I3(n26681), .O(n9024[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4424));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_694_11 (.CI(n25663), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3005[9]), .CO(n25664));
    SB_CARRY add_5037_16 (.CI(n26681), .I0(n9046[13]), .I1(n1105_adj_4368), 
            .CO(n26682));
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17835_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17835_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n25711), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_12 (.CI(n25711), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n25712));
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n25710), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_15_lut (.I0(GND_net), .I1(n9046[12]), .I2(n1032_adj_4344), 
            .I3(n26680), .O(n9024[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_694_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3005[8]), .I3(n25662), .O(\PID_CONTROLLER.integral_23__N_3463 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n25626), .O(duty_23__N_3563[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n25626), .I0(n106[13]), .I1(n155[13]), .CO(n25627));
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n25625), .O(duty_23__N_3563[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_14 (.CI(n25625), .I0(n106[12]), .I1(n155[12]), .CO(n25626));
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5037_15 (.CI(n26680), .I0(n9046[12]), .I1(n1032_adj_4344), 
            .CO(n26681));
    SB_LUT4 add_5037_14_lut (.I0(GND_net), .I1(n9046[11]), .I2(n959_adj_4329), 
            .I3(n26679), .O(n9024[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5037_14 (.CI(n26679), .I0(n9046[11]), .I1(n959_adj_4329), 
            .CO(n26680));
    SB_LUT4 add_5037_13_lut (.I0(GND_net), .I1(n9046[10]), .I2(n886_adj_4328), 
            .I3(n26678), .O(n9024[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_13 (.CI(n26678), .I0(n9046[10]), .I1(n886_adj_4328), 
            .CO(n26679));
    SB_LUT4 add_5037_12_lut (.I0(GND_net), .I1(n9046[9]), .I2(n813_adj_4327), 
            .I3(n26677), .O(n9024[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_12 (.CI(n26677), .I0(n9046[9]), .I1(n813_adj_4327), 
            .CO(n26678));
    SB_LUT4 add_5037_11_lut (.I0(GND_net), .I1(n9046[8]), .I2(n740_adj_4326), 
            .I3(n26676), .O(n9024[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_11 (.CI(n26676), .I0(n9046[8]), .I1(n740_adj_4326), 
            .CO(n26677));
    SB_LUT4 add_5037_10_lut (.I0(GND_net), .I1(n9046[7]), .I2(n667_adj_4325), 
            .I3(n26675), .O(n9024[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_10 (.CI(n26675), .I0(n9046[7]), .I1(n667_adj_4325), 
            .CO(n26676));
    SB_LUT4 add_5037_9_lut (.I0(GND_net), .I1(n9046[6]), .I2(n594_adj_4324), 
            .I3(n26674), .O(n9024[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_9 (.CI(n26674), .I0(n9046[6]), .I1(n594_adj_4324), 
            .CO(n26675));
    SB_LUT4 add_5037_8_lut (.I0(GND_net), .I1(n9046[5]), .I2(n521_adj_4323), 
            .I3(n26673), .O(n9024[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_8 (.CI(n26673), .I0(n9046[5]), .I1(n521_adj_4323), 
            .CO(n26674));
    SB_LUT4 add_5037_7_lut (.I0(GND_net), .I1(n9046[4]), .I2(n448_adj_4322), 
            .I3(n26672), .O(n9024[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_7 (.CI(n26672), .I0(n9046[4]), .I1(n448_adj_4322), 
            .CO(n26673));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n25624), .O(duty_23__N_3563[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28319_4_lut (.I0(n19_adj_4416), .I1(n17_adj_4406), .I2(n15_adj_4403), 
            .I3(n34518), .O(n34493));
    defparam i28319_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5037_6_lut (.I0(GND_net), .I1(n9046[3]), .I2(n375_adj_4321), 
            .I3(n26671), .O(n9024[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n25710), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n25711));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n25709), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n25709), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n25710));
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_694_10 (.CI(n25662), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3005[8]), .CO(n25663));
    SB_CARRY add_12_13 (.CI(n25624), .I0(n106[11]), .I1(n155[11]), .CO(n25625));
    SB_LUT4 i28632_4_lut (.I0(n25_adj_4400), .I1(n23_adj_4399), .I2(n21_adj_4417), 
            .I3(n34493), .O(n34806));
    defparam i28632_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_694_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3005[7]), .I3(n25661), .O(\PID_CONTROLLER.integral_23__N_3463 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28476_4_lut (.I0(n31), .I1(n29_adj_4232), .I2(n27_adj_4404), 
            .I3(n34806), .O(n34650));
    defparam i28476_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_5037_6 (.CI(n26671), .I0(n9046[3]), .I1(n375_adj_4321), 
            .CO(n26672));
    SB_LUT4 add_5037_5_lut (.I0(GND_net), .I1(n9046[2]), .I2(n302_adj_4318), 
            .I3(n26670), .O(n9024[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_5 (.CI(n26670), .I0(n9046[2]), .I1(n302_adj_4318), 
            .CO(n26671));
    SB_LUT4 add_5037_4_lut (.I0(GND_net), .I1(n9046[1]), .I2(n229_adj_4317), 
            .I3(n26669), .O(n9024[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_4 (.CI(n26669), .I0(n9046[1]), .I1(n229_adj_4317), 
            .CO(n26670));
    SB_LUT4 add_5037_3_lut (.I0(GND_net), .I1(n9046[0]), .I2(n156_adj_4316), 
            .I3(n26668), .O(n9024[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_3 (.CI(n26668), .I0(n9046[0]), .I1(n156_adj_4316), 
            .CO(n26669));
    SB_LUT4 add_5037_2_lut (.I0(GND_net), .I1(n14_adj_4315), .I2(n83_adj_4314), 
            .I3(GND_net), .O(n9024[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_2 (.CI(GND_net), .I0(n14_adj_4315), .I1(n83_adj_4314), 
            .CO(n26668));
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_694_9 (.CI(n25661), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3005[7]), .CO(n25662));
    SB_LUT4 i28683_4_lut (.I0(n37), .I1(n35_adj_4235), .I2(n33), .I3(n34650), 
            .O(n34857));
    defparam i28683_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5036_22_lut (.I0(GND_net), .I1(n9024[19]), .I2(GND_net), 
            .I3(n26667), .O(n9001[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5036_21_lut (.I0(GND_net), .I1(n9024[18]), .I2(GND_net), 
            .I3(n26666), .O(n9001[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_21 (.CI(n26666), .I0(n9024[18]), .I1(GND_net), .CO(n26667));
    SB_LUT4 add_5036_20_lut (.I0(GND_net), .I1(n9024[17]), .I2(GND_net), 
            .I3(n26665), .O(n9001[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_20 (.CI(n26665), .I0(n9024[17]), .I1(GND_net), .CO(n26666));
    SB_LUT4 add_5036_19_lut (.I0(GND_net), .I1(n9024[16]), .I2(GND_net), 
            .I3(n26664), .O(n9001[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_19 (.CI(n26664), .I0(n9024[16]), .I1(GND_net), .CO(n26665));
    SB_LUT4 add_5036_18_lut (.I0(GND_net), .I1(n9024[15]), .I2(GND_net), 
            .I3(n26663), .O(n9001[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_18 (.CI(n26663), .I0(n9024[15]), .I1(GND_net), .CO(n26664));
    SB_LUT4 add_5036_17_lut (.I0(GND_net), .I1(n9024[14]), .I2(GND_net), 
            .I3(n26662), .O(n9001[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n25623), .O(duty_23__N_3563[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4218));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5036_17 (.CI(n26662), .I0(n9024[14]), .I1(GND_net), .CO(n26663));
    SB_LUT4 add_5036_16_lut (.I0(GND_net), .I1(n9024[13]), .I2(n1102_adj_4313), 
            .I3(n26661), .O(n9001[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_16 (.CI(n26661), .I0(n9024[13]), .I1(n1102_adj_4313), 
            .CO(n26662));
    SB_LUT4 add_5036_15_lut (.I0(GND_net), .I1(n9024[12]), .I2(n1029_adj_4312), 
            .I3(n26660), .O(n9001[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_15 (.CI(n26660), .I0(n9024[12]), .I1(n1029_adj_4312), 
            .CO(n26661));
    SB_LUT4 add_5036_14_lut (.I0(GND_net), .I1(n9024[11]), .I2(n956_adj_4311), 
            .I3(n26659), .O(n9001[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_14 (.CI(n26659), .I0(n9024[11]), .I1(n956_adj_4311), 
            .CO(n26660));
    SB_LUT4 add_5036_13_lut (.I0(GND_net), .I1(n9024[10]), .I2(n883_adj_4310), 
            .I3(n26658), .O(n9001[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_13 (.CI(n26658), .I0(n9024[10]), .I1(n883_adj_4310), 
            .CO(n26659));
    SB_LUT4 add_5036_12_lut (.I0(GND_net), .I1(n9024[9]), .I2(n810_adj_4309), 
            .I3(n26657), .O(n9001[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_12 (.CI(n26657), .I0(n9024[9]), .I1(n810_adj_4309), 
            .CO(n26658));
    SB_LUT4 add_5036_11_lut (.I0(GND_net), .I1(n9024[8]), .I2(n737_adj_4308), 
            .I3(n26656), .O(n9001[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_11 (.CI(n26656), .I0(n9024[8]), .I1(n737_adj_4308), 
            .CO(n26657));
    SB_LUT4 add_5036_10_lut (.I0(GND_net), .I1(n9024[7]), .I2(n664_adj_4307), 
            .I3(n26655), .O(n9001[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_10 (.CI(n26655), .I0(n9024[7]), .I1(n664_adj_4307), 
            .CO(n26656));
    SB_LUT4 add_5036_9_lut (.I0(GND_net), .I1(n9024[6]), .I2(n591_adj_4306), 
            .I3(n26654), .O(n9001[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_832_i16_3_lut (.I0(duty_23__N_3563[9]), .I1(duty_23__N_3563[21]), 
            .I2(n43), .I3(GND_net), .O(n16_adj_4501));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n25708), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_694_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3005[6]), .I3(n25660), .O(\PID_CONTROLLER.integral_23__N_3463 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n25708), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n25709));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n25707), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_8 (.CI(n25660), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3005[6]), .CO(n25661));
    SB_CARRY sub_3_add_2_8 (.CI(n25707), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n25708));
    SB_LUT4 add_694_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3005[5]), .I3(n25659), .O(\PID_CONTROLLER.integral_23__N_3463 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_7 (.CI(n25659), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3005[5]), .CO(n25660));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n25706), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_694_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3005[4]), .I3(n25658), .O(\PID_CONTROLLER.integral_23__N_3463 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_9 (.CI(n26654), .I0(n9024[6]), .I1(n591_adj_4306), 
            .CO(n26655));
    SB_LUT4 add_5036_8_lut (.I0(GND_net), .I1(n9024[5]), .I2(n518_adj_4302), 
            .I3(n26653), .O(n9001[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_8 (.CI(n26653), .I0(n9024[5]), .I1(n518_adj_4302), 
            .CO(n26654));
    SB_LUT4 add_5036_7_lut (.I0(GND_net), .I1(n9024[4]), .I2(n445_adj_4301), 
            .I3(n26652), .O(n9001[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_7 (.CI(n26652), .I0(n9024[4]), .I1(n445_adj_4301), 
            .CO(n26653));
    SB_LUT4 add_5036_6_lut (.I0(GND_net), .I1(n9024[3]), .I2(n372_adj_4300), 
            .I3(n26651), .O(n9001[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_6 (.CI(n26651), .I0(n9024[3]), .I1(n372_adj_4300), 
            .CO(n26652));
    SB_CARRY add_12_12 (.CI(n25623), .I0(n106[10]), .I1(n155[10]), .CO(n25624));
    SB_LUT4 add_5036_5_lut (.I0(GND_net), .I1(n9024[2]), .I2(n299_adj_4299), 
            .I3(n26650), .O(n9001[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_5 (.CI(n26650), .I0(n9024[2]), .I1(n299_adj_4299), 
            .CO(n26651));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[23]), 
            .I3(n25770), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n25706), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n25707));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[22]), 
            .I3(n25769), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n25705), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n25769), .I0(GND_net), .I1(n1_adj_4633[22]), 
            .CO(n25770));
    SB_CARRY sub_3_add_2_6 (.CI(n25705), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n25706));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n25622), 
            .O(duty_23__N_3563[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[21]), 
            .I3(n25768), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5036_4_lut (.I0(GND_net), .I1(n9024[1]), .I2(n226_adj_4295), 
            .I3(n26649), .O(n9001[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_4 (.CI(n26649), .I0(n9024[1]), .I1(n226_adj_4295), 
            .CO(n26650));
    SB_LUT4 add_5036_3_lut (.I0(GND_net), .I1(n9024[0]), .I2(n153_adj_4293), 
            .I3(n26648), .O(n9001[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_3 (.CI(n26648), .I0(n9024[0]), .I1(n153_adj_4293), 
            .CO(n26649));
    SB_LUT4 add_5036_2_lut (.I0(GND_net), .I1(n11_adj_4292), .I2(n80_adj_4291), 
            .I3(GND_net), .O(n9001[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n25768), .I0(GND_net), .I1(n1_adj_4633[21]), 
            .CO(n25769));
    SB_CARRY add_694_6 (.CI(n25658), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3005[4]), .CO(n25659));
    SB_CARRY add_12_11 (.CI(n25622), .I0(n106[9]), .I1(n155[9]), .CO(n25623));
    SB_CARRY add_5036_2 (.CI(GND_net), .I0(n11_adj_4292), .I1(n80_adj_4291), 
            .CO(n26648));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n8977[21]), .I2(GND_net), 
            .I3(n26647), .O(n7405[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n8977[20]), .I2(GND_net), 
            .I3(n26646), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n26646), .I0(n8977[20]), .I1(GND_net), 
            .CO(n26647));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n8977[19]), .I2(GND_net), 
            .I3(n26645), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n26645), .I0(n8977[19]), .I1(GND_net), 
            .CO(n26646));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n8977[18]), .I2(GND_net), 
            .I3(n26644), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n26644), .I0(n8977[18]), .I1(GND_net), 
            .CO(n26645));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n8977[17]), .I2(GND_net), 
            .I3(n26643), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n26643), .I0(n8977[17]), .I1(GND_net), 
            .CO(n26644));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n8977[16]), .I2(GND_net), 
            .I3(n26642), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n26642), .I0(n8977[16]), .I1(GND_net), 
            .CO(n26643));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n8977[15]), .I2(GND_net), 
            .I3(n26641), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n26641), .I0(n8977[15]), .I1(GND_net), 
            .CO(n26642));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n8977[14]), .I2(GND_net), 
            .I3(n26640), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n26640), .I0(n8977[14]), .I1(GND_net), 
            .CO(n26641));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n8977[13]), .I2(n1096_adj_4290), 
            .I3(n26639), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n26639), .I0(n8977[13]), .I1(n1096_adj_4290), 
            .CO(n26640));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n8977[12]), .I2(n1023_adj_4289), 
            .I3(n26638), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n26638), .I0(n8977[12]), .I1(n1023_adj_4289), 
            .CO(n26639));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[20]), 
            .I3(n25767), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n8977[11]), .I2(n950_adj_4287), 
            .I3(n26637), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n26637), .I0(n8977[11]), .I1(n950_adj_4287), 
            .CO(n26638));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n8977[10]), .I2(n877_adj_4286), 
            .I3(n26636), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n26636), .I0(n8977[10]), .I1(n877_adj_4286), 
            .CO(n26637));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n25767), .I0(GND_net), .I1(n1_adj_4633[20]), 
            .CO(n25768));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n8977[9]), .I2(n804_adj_4285), 
            .I3(n26635), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n26635), .I0(n8977[9]), .I1(n804_adj_4285), 
            .CO(n26636));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n8977[8]), .I2(n731_adj_4284), 
            .I3(n26634), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_694_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3005[3]), .I3(n25657), .O(\PID_CONTROLLER.integral_23__N_3463 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n26634), .I0(n8977[8]), .I1(n731_adj_4284), 
            .CO(n26635));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n8977[7]), .I2(n658_adj_4282), 
            .I3(n26633), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n26633), .I0(n8977[7]), .I1(n658_adj_4282), 
            .CO(n26634));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n8977[6]), .I2(n585_adj_4281), 
            .I3(n26632), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n25621), 
            .O(duty_23__N_3563[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n26632), .I0(n8977[6]), .I1(n585_adj_4281), 
            .CO(n26633));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[19]), 
            .I3(n25766), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n25704), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n8977[5]), .I2(n512_adj_4279), 
            .I3(n26631), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28634_3_lut (.I0(n6_adj_4460), .I1(duty_23__N_3563[10]), .I2(n21_adj_4417), 
            .I3(GND_net), .O(n34808));   // verilog/motorControl.v(36[10:25])
    defparam i28634_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_694_5 (.CI(n25657), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3005[3]), .CO(n25658));
    SB_LUT4 add_694_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3005[2]), .I3(n25656), .O(\PID_CONTROLLER.integral_23__N_3463 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n25766), .I0(GND_net), .I1(n1_adj_4633[19]), 
            .CO(n25767));
    SB_CARRY mult_10_add_1225_8 (.CI(n26631), .I0(n8977[5]), .I1(n512_adj_4279), 
            .CO(n26632));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n8977[4]), .I2(n439_adj_4278), 
            .I3(n26630), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n26630), .I0(n8977[4]), .I1(n439_adj_4278), 
            .CO(n26631));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n8977[3]), .I2(n366_adj_4277), 
            .I3(n26629), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n26629), .I0(n8977[3]), .I1(n366_adj_4277), 
            .CO(n26630));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n8977[2]), .I2(n293_adj_4276), 
            .I3(n26628), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n26628), .I0(n8977[2]), .I1(n293_adj_4276), 
            .CO(n26629));
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4504));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n8977[1]), .I2(n220_adj_4275), 
            .I3(n26627), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n26627), .I0(n8977[1]), .I1(n220_adj_4275), 
            .CO(n26628));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n8977[0]), .I2(n147_adj_4273), 
            .I3(n26626), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n26626), .I0(n8977[0]), .I1(n147_adj_4273), 
            .CO(n26627));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4272), .I2(n74_adj_4271), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4272), .I1(n74_adj_4271), 
            .CO(n26626));
    SB_LUT4 add_5035_23_lut (.I0(GND_net), .I1(n9001[20]), .I2(GND_net), 
            .I3(n26625), .O(n8977[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5035_22_lut (.I0(GND_net), .I1(n9001[19]), .I2(GND_net), 
            .I3(n26624), .O(n8977[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_22 (.CI(n26624), .I0(n9001[19]), .I1(GND_net), .CO(n26625));
    SB_LUT4 add_5035_21_lut (.I0(GND_net), .I1(n9001[18]), .I2(GND_net), 
            .I3(n26623), .O(n8977[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_21 (.CI(n26623), .I0(n9001[18]), .I1(GND_net), .CO(n26624));
    SB_LUT4 add_5035_20_lut (.I0(GND_net), .I1(n9001[17]), .I2(GND_net), 
            .I3(n26622), .O(n8977[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_20 (.CI(n26622), .I0(n9001[17]), .I1(GND_net), .CO(n26623));
    SB_LUT4 add_5035_19_lut (.I0(GND_net), .I1(n9001[16]), .I2(GND_net), 
            .I3(n26621), .O(n8977[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_19 (.CI(n26621), .I0(n9001[16]), .I1(GND_net), .CO(n26622));
    SB_LUT4 add_5035_18_lut (.I0(GND_net), .I1(n9001[15]), .I2(GND_net), 
            .I3(n26620), .O(n8977[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_18 (.CI(n26620), .I0(n9001[15]), .I1(GND_net), .CO(n26621));
    SB_LUT4 add_5035_17_lut (.I0(GND_net), .I1(n9001[14]), .I2(GND_net), 
            .I3(n26619), .O(n8977[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_17 (.CI(n26619), .I0(n9001[14]), .I1(GND_net), .CO(n26620));
    SB_LUT4 add_5035_16_lut (.I0(GND_net), .I1(n9001[13]), .I2(n1099_adj_4270), 
            .I3(n26618), .O(n8977[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_16 (.CI(n26618), .I0(n9001[13]), .I1(n1099_adj_4270), 
            .CO(n26619));
    SB_LUT4 add_5035_15_lut (.I0(GND_net), .I1(n9001[12]), .I2(n1026_adj_4269), 
            .I3(n26617), .O(n8977[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_15 (.CI(n26617), .I0(n9001[12]), .I1(n1026_adj_4269), 
            .CO(n26618));
    SB_LUT4 add_5035_14_lut (.I0(GND_net), .I1(n9001[11]), .I2(n953_adj_4268), 
            .I3(n26616), .O(n8977[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_14 (.CI(n26616), .I0(n9001[11]), .I1(n953_adj_4268), 
            .CO(n26617));
    SB_LUT4 add_5035_13_lut (.I0(GND_net), .I1(n9001[10]), .I2(n880_adj_4267), 
            .I3(n26615), .O(n8977[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_13 (.CI(n26615), .I0(n9001[10]), .I1(n880_adj_4267), 
            .CO(n26616));
    SB_LUT4 add_5035_12_lut (.I0(GND_net), .I1(n9001[9]), .I2(n807_adj_4266), 
            .I3(n26614), .O(n8977[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_12 (.CI(n26614), .I0(n9001[9]), .I1(n807_adj_4266), 
            .CO(n26615));
    SB_LUT4 add_5035_11_lut (.I0(GND_net), .I1(n9001[8]), .I2(n734_adj_4265), 
            .I3(n26613), .O(n8977[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3439[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5035_11 (.CI(n26613), .I0(n9001[8]), .I1(n734_adj_4265), 
            .CO(n26614));
    SB_LUT4 add_5035_10_lut (.I0(GND_net), .I1(n9001[7]), .I2(n661_adj_4264), 
            .I3(n26612), .O(n8977[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_10 (.CI(n26612), .I0(n9001[7]), .I1(n661_adj_4264), 
            .CO(n26613));
    SB_LUT4 add_5035_9_lut (.I0(GND_net), .I1(n9001[6]), .I2(n588_adj_4263), 
            .I3(n26611), .O(n8977[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_9 (.CI(n26611), .I0(n9001[6]), .I1(n588_adj_4263), 
            .CO(n26612));
    SB_LUT4 add_5035_8_lut (.I0(GND_net), .I1(n9001[5]), .I2(n515_adj_4262), 
            .I3(n26610), .O(n8977[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_8 (.CI(n26610), .I0(n9001[5]), .I1(n515_adj_4262), 
            .CO(n26611));
    SB_LUT4 add_5035_7_lut (.I0(GND_net), .I1(n9001[4]), .I2(n442_adj_4261), 
            .I3(n26609), .O(n8977[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_7 (.CI(n26609), .I0(n9001[4]), .I1(n442_adj_4261), 
            .CO(n26610));
    SB_LUT4 add_5035_6_lut (.I0(GND_net), .I1(n9001[3]), .I2(n369_adj_4260), 
            .I3(n26608), .O(n8977[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_6 (.CI(n26608), .I0(n9001[3]), .I1(n369_adj_4260), 
            .CO(n26609));
    SB_CARRY add_12_10 (.CI(n25621), .I0(n106[8]), .I1(n155[8]), .CO(n25622));
    SB_LUT4 add_5035_5_lut (.I0(GND_net), .I1(n9001[2]), .I2(n296_adj_4259), 
            .I3(n26607), .O(n8977[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_5 (.CI(n26607), .I0(n9001[2]), .I1(n296_adj_4259), 
            .CO(n26608));
    SB_LUT4 add_5035_4_lut (.I0(GND_net), .I1(n9001[1]), .I2(n223_adj_4258), 
            .I3(n26606), .O(n8977[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_4 (.CI(n26606), .I0(n9001[1]), .I1(n223_adj_4258), 
            .CO(n26607));
    SB_LUT4 add_5035_3_lut (.I0(GND_net), .I1(n9001[0]), .I2(n150_adj_4257), 
            .I3(n26605), .O(n8977[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_3 (.CI(n26605), .I0(n9001[0]), .I1(n150_adj_4257), 
            .CO(n26606));
    SB_LUT4 i28635_3_lut (.I0(n34808), .I1(duty_23__N_3563[11]), .I2(n23_adj_4399), 
            .I3(GND_net), .O(n34809));   // verilog/motorControl.v(36[10:25])
    defparam i28635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5035_2_lut (.I0(GND_net), .I1(n8_adj_4256), .I2(n77_adj_4254), 
            .I3(GND_net), .O(n8977[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5035_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5035_2 (.CI(GND_net), .I0(n8_adj_4256), .I1(n77_adj_4254), 
            .CO(n26605));
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3439[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3439[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3439[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3439[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3439[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3439[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3439[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3439[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3439[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3439[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3439[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3439[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3439[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3439[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3439[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3439[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3439[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3439[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3439[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3439[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3439[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3463 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 duty_23__I_832_i8_3_lut (.I0(duty_23__N_3563[4]), .I1(duty_23__N_3563[8]), 
            .I2(n17_adj_4406), .I3(GND_net), .O(n8_adj_4505));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i24_3_lut (.I0(n16_adj_4501), .I1(duty_23__N_3563[22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_4506));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[18]), 
            .I3(n25765), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n25765), .I0(GND_net), .I1(n1_adj_4633[18]), 
            .CO(n25766));
    SB_LUT4 i28018_4_lut (.I0(n43), .I1(n25_adj_4400), .I2(n23_adj_4399), 
            .I3(n34214), .O(n34190));
    defparam i28018_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n25620), 
            .O(duty_23__N_3563[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[17]), 
            .I3(n25764), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_4 (.CI(n25656), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3005[2]), .CO(n25657));
    SB_LUT4 i28488_4_lut (.I0(n24_adj_4506), .I1(n8_adj_4505), .I2(n45), 
            .I3(n34188), .O(n34662));   // verilog/motorControl.v(36[10:25])
    defparam i28488_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n25764), .I0(GND_net), .I1(n1_adj_4633[17]), 
            .CO(n25765));
    SB_CARRY sub_3_add_2_5 (.CI(n25704), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n25705));
    SB_LUT4 i28016_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3563[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3563[9]), .O(n34188));
    defparam i28016_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i28559_3_lut (.I0(n34809), .I1(duty_23__N_3563[12]), .I2(n25_adj_4400), 
            .I3(GND_net), .O(n34733));   // verilog/motorControl.v(36[10:25])
    defparam i28559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20840_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I2(n4_adj_4507), .I3(n9553[1]), .O(n6_adj_4508));   // verilog/motorControl.v(34[25:36])
    defparam i20840_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 duty_23__I_832_i4_4_lut (.I0(duty_23__N_3563[0]), .I1(duty_23__N_3563[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4509));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i28626_3_lut (.I0(n4_adj_4509), .I1(duty_23__N_3563[13]), .I2(n27_adj_4404), 
            .I3(GND_net), .O(n34800));   // verilog/motorControl.v(36[10:25])
    defparam i28626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I2(n9553[1]), .I3(n4_adj_4507), .O(n9546[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1480 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [19]), 
            .I2(n9559[0]), .I3(n25430), .O(n9553[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1480.LUT_INIT = 16'h8778;
    SB_LUT4 i20871_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [19]), 
            .I2(n25430), .I3(n9559[0]), .O(n4_adj_4510));   // verilog/motorControl.v(34[25:36])
    defparam i20871_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20858_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [19]), .I3(\Ki[1] ), 
            .O(n9553[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20858_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[16]), 
            .I3(n25763), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n25763), .I0(GND_net), .I1(n1_adj_4633[16]), 
            .CO(n25764));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n25703), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20860_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [19]), .I3(\Ki[1] ), 
            .O(n25430));   // verilog/motorControl.v(34[25:36])
    defparam i20860_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_694_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3005[1]), .I3(n25655), .O(\PID_CONTROLLER.integral_23__N_3463 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_3 (.CI(n25655), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3005[1]), .CO(n25656));
    SB_CARRY sub_3_add_2_4 (.CI(n25703), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n25704));
    SB_CARRY add_12_9 (.CI(n25620), .I0(n106[7]), .I1(n155[7]), .CO(n25621));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[15]), 
            .I3(n25762), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_694_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3005[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3463 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_694_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_694_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3005[0]), .CO(n25655));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n25702), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n25619), 
            .O(duty_23__N_3563[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20902_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [20]), 
            .I2(n25464), .I3(n9564[0]), .O(n4_adj_4511));   // verilog/motorControl.v(34[25:36])
    defparam i20902_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [20]), 
            .I2(n9564[0]), .I3(n25464), .O(n9559[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h8778;
    SB_LUT4 i20889_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [20]), .I3(\Ki[1] ), 
            .O(n9559[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20889_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20891_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [20]), .I3(\Ki[1] ), 
            .O(n25464));   // verilog/motorControl.v(34[25:36])
    defparam i20891_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_3_lut_4_lut_adj_1482 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I2(n9553[0]), .I3(n25387), .O(n9546[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1482.LUT_INIT = 16'h8778;
    SB_LUT4 i20832_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I2(n25387), .I3(n9553[0]), .O(n4_adj_4507));   // verilog/motorControl.v(34[25:36])
    defparam i20832_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20821_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [18]), .I3(\Ki[1] ), 
            .O(n25387));   // verilog/motorControl.v(34[25:36])
    defparam i20821_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20819_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3463 [18]), .I3(\Ki[1] ), 
            .O(n9546[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20819_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28027_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3563[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3563[7]), .O(n34199));
    defparam i28027_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i27982_2_lut_4_lut (.I0(duty_23__N_3563[21]), .I1(n257[21]), 
            .I2(duty_23__N_3563[9]), .I3(n257[9]), .O(n34154));
    defparam i27982_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i27992_2_lut_4_lut (.I0(duty_23__N_3563[16]), .I1(n257[16]), 
            .I2(duty_23__N_3563[7]), .I3(n257[7]), .O(n34164));
    defparam i27992_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4418));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5073_7_lut (.I0(GND_net), .I1(n32845), .I2(n490_adj_4512), 
            .I3(n27090), .O(n9538[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5073_6_lut (.I0(GND_net), .I1(n9546[3]), .I2(n417_adj_4513), 
            .I3(n27089), .O(n9538[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_6 (.CI(n27089), .I0(n9546[3]), .I1(n417_adj_4513), 
            .CO(n27090));
    SB_LUT4 add_5073_5_lut (.I0(GND_net), .I1(n9546[2]), .I2(n344_adj_4514), 
            .I3(n27088), .O(n9538[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_5 (.CI(n27088), .I0(n9546[2]), .I1(n344_adj_4514), 
            .CO(n27089));
    SB_LUT4 i17836_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17836_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5073_4_lut (.I0(GND_net), .I1(n9546[1]), .I2(n271_adj_4515), 
            .I3(n27087), .O(n9538[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_4 (.CI(n27087), .I0(n9546[1]), .I1(n271_adj_4515), 
            .CO(n27088));
    SB_LUT4 add_5073_3_lut (.I0(GND_net), .I1(n9546[0]), .I2(n198_adj_4516), 
            .I3(n27086), .O(n9538[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_3 (.CI(n27086), .I0(n9546[0]), .I1(n198_adj_4516), 
            .CO(n27087));
    SB_LUT4 add_5073_2_lut (.I0(GND_net), .I1(n56_adj_4517), .I2(n125_adj_4518), 
            .I3(GND_net), .O(n9538[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5073_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5073_2 (.CI(GND_net), .I0(n56_adj_4517), .I1(n125_adj_4518), 
            .CO(n27086));
    SB_LUT4 add_5072_8_lut (.I0(GND_net), .I1(n9538[5]), .I2(n560_adj_4519), 
            .I3(n27085), .O(n9529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5072_7_lut (.I0(GND_net), .I1(n9538[4]), .I2(n487_adj_4520), 
            .I3(n27084), .O(n9529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_7 (.CI(n27084), .I0(n9538[4]), .I1(n487_adj_4520), 
            .CO(n27085));
    SB_LUT4 add_5072_6_lut (.I0(GND_net), .I1(n9538[3]), .I2(n414_adj_4521), 
            .I3(n27083), .O(n9529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_6 (.CI(n27083), .I0(n9538[3]), .I1(n414_adj_4521), 
            .CO(n27084));
    SB_LUT4 add_5072_5_lut (.I0(GND_net), .I1(n9538[2]), .I2(n341_adj_4522), 
            .I3(n27082), .O(n9529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_5 (.CI(n27082), .I0(n9538[2]), .I1(n341_adj_4522), 
            .CO(n27083));
    SB_LUT4 add_5072_4_lut (.I0(GND_net), .I1(n9538[1]), .I2(n268_adj_4523), 
            .I3(n27081), .O(n9529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_4 (.CI(n27081), .I0(n9538[1]), .I1(n268_adj_4523), 
            .CO(n27082));
    SB_LUT4 add_5072_3_lut (.I0(GND_net), .I1(n9538[0]), .I2(n195_adj_4524), 
            .I3(n27080), .O(n9529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_3 (.CI(n27080), .I0(n9538[0]), .I1(n195_adj_4524), 
            .CO(n27081));
    SB_LUT4 add_5072_2_lut (.I0(GND_net), .I1(n53_adj_4525), .I2(n122_adj_4526), 
            .I3(GND_net), .O(n9529[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5072_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5072_2 (.CI(GND_net), .I0(n53_adj_4525), .I1(n122_adj_4526), 
            .CO(n27080));
    SB_LUT4 add_5071_9_lut (.I0(GND_net), .I1(n9529[6]), .I2(n630_adj_4527), 
            .I3(n27079), .O(n9519[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5071_8_lut (.I0(GND_net), .I1(n9529[5]), .I2(n557_adj_4528), 
            .I3(n27078), .O(n9519[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_8 (.CI(n27078), .I0(n9529[5]), .I1(n557_adj_4528), 
            .CO(n27079));
    SB_LUT4 add_5071_7_lut (.I0(GND_net), .I1(n9529[4]), .I2(n484_adj_4529), 
            .I3(n27077), .O(n9519[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_7 (.CI(n27077), .I0(n9529[4]), .I1(n484_adj_4529), 
            .CO(n27078));
    SB_LUT4 add_5071_6_lut (.I0(GND_net), .I1(n9529[3]), .I2(n411_adj_4530), 
            .I3(n27076), .O(n9519[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_6 (.CI(n27076), .I0(n9529[3]), .I1(n411_adj_4530), 
            .CO(n27077));
    SB_LUT4 add_5071_5_lut (.I0(GND_net), .I1(n9529[2]), .I2(n338_adj_4531), 
            .I3(n27075), .O(n9519[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_5 (.CI(n27075), .I0(n9529[2]), .I1(n338_adj_4531), 
            .CO(n27076));
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5071_4_lut (.I0(GND_net), .I1(n9529[1]), .I2(n265_adj_4532), 
            .I3(n27074), .O(n9519[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_4 (.CI(n27074), .I0(n9529[1]), .I1(n265_adj_4532), 
            .CO(n27075));
    SB_LUT4 add_5071_3_lut (.I0(GND_net), .I1(n9529[0]), .I2(n192_adj_4533), 
            .I3(n27073), .O(n9519[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_3 (.CI(n27073), .I0(n9529[0]), .I1(n192_adj_4533), 
            .CO(n27074));
    SB_LUT4 add_5071_2_lut (.I0(GND_net), .I1(n50_adj_4534), .I2(n119_adj_4535), 
            .I3(GND_net), .O(n9519[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5071_2 (.CI(GND_net), .I0(n50_adj_4534), .I1(n119_adj_4535), 
            .CO(n27073));
    SB_LUT4 add_5070_10_lut (.I0(GND_net), .I1(n9519[7]), .I2(n700_adj_4536), 
            .I3(n27072), .O(n9508[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_9_lut (.I0(GND_net), .I1(n9519[6]), .I2(n627_adj_4537), 
            .I3(n27071), .O(n9508[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_9 (.CI(n27071), .I0(n9519[6]), .I1(n627_adj_4537), 
            .CO(n27072));
    SB_LUT4 add_5070_8_lut (.I0(GND_net), .I1(n9519[5]), .I2(n554_adj_4538), 
            .I3(n27070), .O(n9508[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_8 (.CI(n27070), .I0(n9519[5]), .I1(n554_adj_4538), 
            .CO(n27071));
    SB_LUT4 add_5070_7_lut (.I0(GND_net), .I1(n9519[4]), .I2(n481_adj_4539), 
            .I3(n27069), .O(n9508[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_7 (.CI(n27069), .I0(n9519[4]), .I1(n481_adj_4539), 
            .CO(n27070));
    SB_LUT4 add_5070_6_lut (.I0(GND_net), .I1(n9519[3]), .I2(n408_adj_4540), 
            .I3(n27068), .O(n9508[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_6 (.CI(n27068), .I0(n9519[3]), .I1(n408_adj_4540), 
            .CO(n27069));
    SB_LUT4 add_5070_5_lut (.I0(GND_net), .I1(n9519[2]), .I2(n335_adj_4541), 
            .I3(n27067), .O(n9508[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_5 (.CI(n27067), .I0(n9519[2]), .I1(n335_adj_4541), 
            .CO(n27068));
    SB_LUT4 add_5070_4_lut (.I0(GND_net), .I1(n9519[1]), .I2(n262_adj_4542), 
            .I3(n27066), .O(n9508[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_4 (.CI(n27066), .I0(n9519[1]), .I1(n262_adj_4542), 
            .CO(n27067));
    SB_LUT4 add_5070_3_lut (.I0(GND_net), .I1(n9519[0]), .I2(n189_adj_4543), 
            .I3(n27065), .O(n9508[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_3 (.CI(n27065), .I0(n9519[0]), .I1(n189_adj_4543), 
            .CO(n27066));
    SB_LUT4 add_5070_2_lut (.I0(GND_net), .I1(n47_adj_4544), .I2(n116_adj_4545), 
            .I3(GND_net), .O(n9508[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_2 (.CI(GND_net), .I0(n47_adj_4544), .I1(n116_adj_4545), 
            .CO(n27065));
    SB_LUT4 add_5069_11_lut (.I0(GND_net), .I1(n9508[8]), .I2(n770_adj_4546), 
            .I3(n27064), .O(n9496[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_10_lut (.I0(GND_net), .I1(n9508[7]), .I2(n697_adj_4547), 
            .I3(n27063), .O(n9496[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_10 (.CI(n27063), .I0(n9508[7]), .I1(n697_adj_4547), 
            .CO(n27064));
    SB_LUT4 add_5069_9_lut (.I0(GND_net), .I1(n9508[6]), .I2(n624_adj_4548), 
            .I3(n27062), .O(n9496[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_9 (.CI(n27062), .I0(n9508[6]), .I1(n624_adj_4548), 
            .CO(n27063));
    SB_LUT4 add_5069_8_lut (.I0(GND_net), .I1(n9508[5]), .I2(n551_adj_4549), 
            .I3(n27061), .O(n9496[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_8 (.CI(n27061), .I0(n9508[5]), .I1(n551_adj_4549), 
            .CO(n27062));
    SB_LUT4 add_5069_7_lut (.I0(GND_net), .I1(n9508[4]), .I2(n478_adj_4550), 
            .I3(n27060), .O(n9496[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_7 (.CI(n27060), .I0(n9508[4]), .I1(n478_adj_4550), 
            .CO(n27061));
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4551));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5069_6_lut (.I0(GND_net), .I1(n9508[3]), .I2(n405_adj_4552), 
            .I3(n27059), .O(n9496[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_6 (.CI(n27059), .I0(n9508[3]), .I1(n405_adj_4552), 
            .CO(n27060));
    SB_LUT4 add_5069_5_lut (.I0(GND_net), .I1(n9508[2]), .I2(n332_adj_4553), 
            .I3(n27058), .O(n9496[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_5 (.CI(n27058), .I0(n9508[2]), .I1(n332_adj_4553), 
            .CO(n27059));
    SB_LUT4 add_5069_4_lut (.I0(GND_net), .I1(n9508[1]), .I2(n259_adj_4554), 
            .I3(n27057), .O(n9496[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_4 (.CI(n27057), .I0(n9508[1]), .I1(n259_adj_4554), 
            .CO(n27058));
    SB_LUT4 add_5069_3_lut (.I0(GND_net), .I1(n9508[0]), .I2(n186_adj_4555), 
            .I3(n27056), .O(n9496[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_3 (.CI(n27056), .I0(n9508[0]), .I1(n186_adj_4555), 
            .CO(n27057));
    SB_LUT4 add_5069_2_lut (.I0(GND_net), .I1(n44_adj_4556), .I2(n113_adj_4557), 
            .I3(GND_net), .O(n9496[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_2 (.CI(GND_net), .I0(n44_adj_4556), .I1(n113_adj_4557), 
            .CO(n27056));
    SB_LUT4 add_5068_12_lut (.I0(GND_net), .I1(n9496[9]), .I2(n840_adj_4558), 
            .I3(n27055), .O(n9483[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5068_11_lut (.I0(GND_net), .I1(n9496[8]), .I2(n767_adj_4559), 
            .I3(n27054), .O(n9483[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_11 (.CI(n27054), .I0(n9496[8]), .I1(n767_adj_4559), 
            .CO(n27055));
    SB_LUT4 add_5068_10_lut (.I0(GND_net), .I1(n9496[7]), .I2(n694_adj_4560), 
            .I3(n27053), .O(n9483[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_10 (.CI(n27053), .I0(n9496[7]), .I1(n694_adj_4560), 
            .CO(n27054));
    SB_LUT4 add_5068_9_lut (.I0(GND_net), .I1(n9496[6]), .I2(n621_adj_4561), 
            .I3(n27052), .O(n9483[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_9 (.CI(n27052), .I0(n9496[6]), .I1(n621_adj_4561), 
            .CO(n27053));
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4562));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5068_8_lut (.I0(GND_net), .I1(n9496[5]), .I2(n548_adj_4563), 
            .I3(n27051), .O(n9483[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4564));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5068_8 (.CI(n27051), .I0(n9496[5]), .I1(n548_adj_4563), 
            .CO(n27052));
    SB_LUT4 add_5068_7_lut (.I0(GND_net), .I1(n9496[4]), .I2(n475_adj_4565), 
            .I3(n27050), .O(n9483[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28160_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n34332));
    defparam i28160_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_5068_7 (.CI(n27050), .I0(n9496[4]), .I1(n475_adj_4565), 
            .CO(n27051));
    SB_LUT4 add_5068_6_lut (.I0(GND_net), .I1(n9496[3]), .I2(n402_adj_4566), 
            .I3(n27049), .O(n9483[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_6 (.CI(n27049), .I0(n9496[3]), .I1(n402_adj_4566), 
            .CO(n27050));
    SB_LUT4 i28157_3_lut (.I0(n11_adj_4564), .I1(n9_adj_4562), .I2(n34332), 
            .I3(GND_net), .O(n34329));
    defparam i28157_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 add_5068_5_lut (.I0(GND_net), .I1(n9496[2]), .I2(n329_adj_4567), 
            .I3(n27048), .O(n9483[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_171_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n36254));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_171_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5068_5 (.CI(n27048), .I0(n9496[2]), .I1(n329_adj_4567), 
            .CO(n27049));
    SB_LUT4 add_5068_4_lut (.I0(GND_net), .I1(n9496[1]), .I2(n256_adj_4568), 
            .I3(n27047), .O(n9483[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_4 (.CI(n27047), .I0(n9496[1]), .I1(n256_adj_4568), 
            .CO(n27048));
    SB_LUT4 add_5068_3_lut (.I0(GND_net), .I1(n9496[0]), .I2(n183_adj_4569), 
            .I3(n27046), .O(n9483[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_3 (.CI(n27046), .I0(n9496[0]), .I1(n183_adj_4569), 
            .CO(n27047));
    SB_LUT4 add_5068_2_lut (.I0(GND_net), .I1(n41_adj_4570), .I2(n110_adj_4571), 
            .I3(GND_net), .O(n9483[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28524_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n36254), 
            .I2(IntegralLimit[7]), .I3(n34329), .O(n34698));
    defparam i28524_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5068_2 (.CI(GND_net), .I0(n41_adj_4570), .I1(n110_adj_4571), 
            .CO(n27046));
    SB_LUT4 add_5067_13_lut (.I0(GND_net), .I1(n9483[10]), .I2(n910_adj_4572), 
            .I3(n27045), .O(n9469[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5067_12_lut (.I0(GND_net), .I1(n9483[9]), .I2(n837_adj_4573), 
            .I3(n27044), .O(n9469[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_12 (.CI(n27044), .I0(n9483[9]), .I1(n837_adj_4573), 
            .CO(n27045));
    SB_LUT4 i28404_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4551), 
            .I2(IntegralLimit[9]), .I3(n34698), .O(n34578));
    defparam i28404_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5067_11_lut (.I0(GND_net), .I1(n9483[8]), .I2(n764_adj_4574), 
            .I3(n27043), .O(n9469[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_11 (.CI(n27043), .I0(n9483[8]), .I1(n764_adj_4574), 
            .CO(n27044));
    SB_LUT4 add_5067_10_lut (.I0(GND_net), .I1(n9483[7]), .I2(n691_adj_4575), 
            .I3(n27042), .O(n9469[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_10 (.CI(n27042), .I0(n9483[7]), .I1(n691_adj_4575), 
            .CO(n27043));
    SB_LUT4 add_5067_9_lut (.I0(GND_net), .I1(n9483[6]), .I2(n618_adj_4576), 
            .I3(n27041), .O(n9469[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_153_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n36236));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_153_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5067_9 (.CI(n27041), .I0(n9483[6]), .I1(n618_adj_4576), 
            .CO(n27042));
    SB_LUT4 add_5067_8_lut (.I0(GND_net), .I1(n9483[5]), .I2(n545_adj_4577), 
            .I3(n27040), .O(n9469[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_8 (.CI(n27040), .I0(n9483[5]), .I1(n545_adj_4577), 
            .CO(n27041));
    SB_LUT4 add_5067_7_lut (.I0(GND_net), .I1(n9483[4]), .I2(n472_adj_4578), 
            .I3(n27039), .O(n9469[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28402_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4551), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4562), .O(n34576));
    defparam i28402_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5067_7 (.CI(n27039), .I0(n9483[4]), .I1(n472_adj_4578), 
            .CO(n27040));
    SB_LUT4 add_5067_6_lut (.I0(GND_net), .I1(n9483[3]), .I2(n399_adj_4579), 
            .I3(n27038), .O(n9469[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_6 (.CI(n27038), .I0(n9483[3]), .I1(n399_adj_4579), 
            .CO(n27039));
    SB_LUT4 add_5067_5_lut (.I0(GND_net), .I1(n9483[2]), .I2(n326_adj_4580), 
            .I3(n27037), .O(n9469[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_5 (.CI(n27037), .I0(n9483[2]), .I1(n326_adj_4580), 
            .CO(n27038));
    SB_LUT4 i28400_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n36236), 
            .I2(IntegralLimit[11]), .I3(n34576), .O(n34574));
    defparam i28400_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5067_4_lut (.I0(GND_net), .I1(n9483[1]), .I2(n253_adj_4581), 
            .I3(n27036), .O(n9469[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_4 (.CI(n27036), .I0(n9483[1]), .I1(n253_adj_4581), 
            .CO(n27037));
    SB_LUT4 add_5067_3_lut (.I0(GND_net), .I1(n9483[0]), .I2(n180_adj_4582), 
            .I3(n27035), .O(n9469[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_3 (.CI(n27035), .I0(n9483[0]), .I1(n180_adj_4582), 
            .CO(n27036));
    SB_LUT4 add_5067_2_lut (.I0(GND_net), .I1(n38_adj_4583), .I2(n107_adj_4584), 
            .I3(GND_net), .O(n9469[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5067_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5067_2 (.CI(GND_net), .I0(n38_adj_4583), .I1(n107_adj_4584), 
            .CO(n27035));
    SB_LUT4 add_5066_14_lut (.I0(GND_net), .I1(n9469[11]), .I2(n980_adj_4585), 
            .I3(n27034), .O(n9454[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5066_13_lut (.I0(GND_net), .I1(n9469[10]), .I2(n907_adj_4586), 
            .I3(n27033), .O(n9454[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_13 (.CI(n27033), .I0(n9469[10]), .I1(n907_adj_4586), 
            .CO(n27034));
    SB_LUT4 add_5066_12_lut (.I0(GND_net), .I1(n9469[9]), .I2(n834_adj_4587), 
            .I3(n27032), .O(n9454[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_12 (.CI(n27032), .I0(n9469[9]), .I1(n834_adj_4587), 
            .CO(n27033));
    SB_LUT4 add_5066_11_lut (.I0(GND_net), .I1(n9469[8]), .I2(n761_adj_4588), 
            .I3(n27031), .O(n9454[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_11 (.CI(n27031), .I0(n9469[8]), .I1(n761_adj_4588), 
            .CO(n27032));
    SB_LUT4 add_5066_10_lut (.I0(GND_net), .I1(n9469[7]), .I2(n688_adj_4589), 
            .I3(n27030), .O(n9454[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_10 (.CI(n27030), .I0(n9469[7]), .I1(n688_adj_4589), 
            .CO(n27031));
    SB_LUT4 add_5066_9_lut (.I0(GND_net), .I1(n9469[6]), .I2(n615_adj_4590), 
            .I3(n27029), .O(n9454[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_9 (.CI(n27029), .I0(n9469[6]), .I1(n615_adj_4590), 
            .CO(n27030));
    SB_LUT4 add_5066_8_lut (.I0(GND_net), .I1(n9469[5]), .I2(n542_adj_4591), 
            .I3(n27028), .O(n9454[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_8 (.CI(n27028), .I0(n9469[5]), .I1(n542_adj_4591), 
            .CO(n27029));
    SB_LUT4 add_5066_7_lut (.I0(GND_net), .I1(n9469[4]), .I2(n469_adj_4592), 
            .I3(n27027), .O(n9454[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_7 (.CI(n27027), .I0(n9469[4]), .I1(n469_adj_4592), 
            .CO(n27028));
    SB_LUT4 add_5066_6_lut (.I0(GND_net), .I1(n9469[3]), .I2(n396_adj_4593), 
            .I3(n27026), .O(n9454[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_6 (.CI(n27026), .I0(n9469[3]), .I1(n396_adj_4593), 
            .CO(n27027));
    SB_LUT4 add_5066_5_lut (.I0(GND_net), .I1(n9469[2]), .I2(n323_adj_4594), 
            .I3(n27025), .O(n9454[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_5 (.CI(n27025), .I0(n9469[2]), .I1(n323_adj_4594), 
            .CO(n27026));
    SB_LUT4 add_5066_4_lut (.I0(GND_net), .I1(n9469[1]), .I2(n250_adj_4595), 
            .I3(n27024), .O(n9454[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_4 (.CI(n27024), .I0(n9469[1]), .I1(n250_adj_4595), 
            .CO(n27025));
    SB_LUT4 add_5066_3_lut (.I0(GND_net), .I1(n9469[0]), .I2(n177_adj_4596), 
            .I3(n27023), .O(n9454[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5066_3 (.CI(n27023), .I0(n9469[0]), .I1(n177_adj_4596), 
            .CO(n27024));
    SB_LUT4 add_5066_2_lut (.I0(GND_net), .I1(n35_adj_4597), .I2(n104_adj_4598), 
            .I3(GND_net), .O(n9454[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5066_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5066_2 (.CI(GND_net), .I0(n35_adj_4597), .I1(n104_adj_4598), 
            .CO(n27023));
    SB_LUT4 add_5065_15_lut (.I0(GND_net), .I1(n9454[12]), .I2(n1050_adj_4600), 
            .I3(n27022), .O(n9438[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5065_14_lut (.I0(GND_net), .I1(n9454[11]), .I2(n977_adj_4601), 
            .I3(n27021), .O(n9438[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5065_12_lut (.I0(GND_net), .I1(n9454[9]), .I2(n831), .I3(n27019), 
            .O(n9438[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n25702), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n25703));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_147_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n36230));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_147_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28082_4_lut (.I0(n27), .I1(n15_adj_4366), .I2(n13_adj_4392), 
            .I3(n11_adj_4412), .O(n34254));
    defparam i28082_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28088_4_lut (.I0(n21_adj_4353), .I1(n19_adj_4354), .I2(n17_adj_4362), 
            .I3(n9_adj_4414), .O(n34260));
    defparam i28088_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n25762), .I0(GND_net), .I1(n1_adj_4633[15]), 
            .CO(n25763));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[14]), 
            .I3(n25761), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_4320), .I3(GND_net), 
            .O(n16_adj_4605));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i28057_2_lut (.I0(n43_adj_4320), .I1(n19_adj_4354), .I2(GND_net), 
            .I3(GND_net), .O(n34229));
    defparam i28057_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n25702));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n25761), .I0(GND_net), .I1(n1_adj_4633[14]), 
            .CO(n25762));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4362), .I3(GND_net), 
            .O(n8_adj_4607));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4605), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_4319), .I3(GND_net), 
            .O(n24_adj_4609));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i28101_2_lut (.I0(n7_adj_4419), .I1(n5_adj_4421), .I2(GND_net), 
            .I3(GND_net), .O(n34273));
    defparam i28101_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_12_8 (.CI(n25619), .I0(n106[6]), .I1(n155[6]), .CO(n25620));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[13]), 
            .I3(n25760), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28376_4_lut (.I0(n13_adj_4392), .I1(n11_adj_4412), .I2(n9_adj_4414), 
            .I3(n34273), .O(n34550));
    defparam i28376_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n25760), .I0(GND_net), .I1(n1_adj_4633[13]), 
            .CO(n25761));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[12]), 
            .I3(n25759), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n25759), .I0(GND_net), .I1(n1_adj_4633[12]), 
            .CO(n25760));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[11]), 
            .I3(n25758), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28372_4_lut (.I0(n19_adj_4354), .I1(n17_adj_4362), .I2(n15_adj_4366), 
            .I3(n34550), .O(n34546));
    defparam i28372_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n25758), .I0(GND_net), .I1(n1_adj_4633[11]), 
            .CO(n25759));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[10]), 
            .I3(n25757), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n25757), .I0(GND_net), .I1(n1_adj_4633[10]), 
            .CO(n25758));
    SB_LUT4 i28658_4_lut (.I0(n25_adj_4351), .I1(n23_adj_4352), .I2(n21_adj_4353), 
            .I3(n34546), .O(n34832));
    defparam i28658_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28502_4_lut (.I0(n31_adj_4348), .I1(n29_adj_4350), .I2(n27), 
            .I3(n34832), .O(n34676));
    defparam i28502_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[9]), 
            .I3(n25756), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n25756), .I0(GND_net), .I1(n1_adj_4633[9]), 
            .CO(n25757));
    SB_LUT4 i28689_4_lut (.I0(n37_adj_4345), .I1(n35_adj_4346), .I2(n33_adj_4347), 
            .I3(n34676), .O(n34863));
    defparam i28689_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[8]), 
            .I3(n25755), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n25755), .I0(GND_net), .I1(n1_adj_4633[8]), 
            .CO(n25756));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n25618), 
            .O(duty_23__N_3563[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[7]), 
            .I3(n25754), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n25754), .I0(GND_net), .I1(n1_adj_4633[7]), 
            .CO(n25755));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[6]), 
            .I3(n25753), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28406_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n36254), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4564), .O(n34580));
    defparam i28406_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_140_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n36223));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_140_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_7 (.CI(n25618), .I0(n106[5]), .I1(n155[5]), .CO(n25619));
    SB_LUT4 i28394_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n36223), 
            .I2(IntegralLimit[14]), .I3(n34580), .O(n34568));
    defparam i28394_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_135_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n36218));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_135_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4613));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28116_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n34288));
    defparam i28116_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_158_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n36241));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_158_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4614));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4613), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4615));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28590_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n36236), 
            .I2(IntegralLimit[11]), .I3(n34578), .O(n34764));
    defparam i28590_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n25753), .I0(GND_net), .I1(n1_adj_4633[6]), 
            .CO(n25754));
    SB_LUT4 i28140_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n36230), 
            .I2(IntegralLimit[13]), .I3(n34764), .O(n34312));
    defparam i28140_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_138_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n36221));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_138_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28518_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n36221), 
            .I2(IntegralLimit[15]), .I3(n34312), .O(n34692));
    defparam i28518_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_164_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n36247));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_164_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28663_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n36247), 
            .I2(IntegralLimit[17]), .I3(n34692), .O(n34837));
    defparam i28663_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_129_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n36212));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_129_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n25617), 
            .O(duty_23__N_3563[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28717_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n36212), 
            .I2(IntegralLimit[19]), .I3(n34837), .O(n34891));
    defparam i28717_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_126_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n36209));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_126_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4616));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28103_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n34275));
    defparam i28103_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[5]), 
            .I3(n25752), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n25752), .I0(GND_net), .I1(n1_adj_4633[5]), 
            .CO(n25753));
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4616), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4617));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4618));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28542_3_lut (.I0(n6_adj_4618), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n34716));   // verilog/motorControl.v(31[10:34])
    defparam i28542_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28543_3_lut (.I0(n34716), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n34717));   // verilog/motorControl.v(31[10:34])
    defparam i28543_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4633[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28105_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n36230), 
            .I2(IntegralLimit[21]), .I3(n34574), .O(n34277));
    defparam i28105_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_123_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n36206));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_123_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[4]), 
            .I3(n25751), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28484_4_lut (.I0(n24_adj_4617), .I1(n8_adj_4504), .I2(n36206), 
            .I3(n34275), .O(n34658));   // verilog/motorControl.v(31[10:34])
    defparam i28484_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28324_3_lut (.I0(n34717), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n34498));   // verilog/motorControl.v(31[10:34])
    defparam i28324_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3514 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4443), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4619));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i28532_3_lut (.I0(n4_adj_4619), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n34706));   // verilog/motorControl.v(31[38:63])
    defparam i28532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28533_3_lut (.I0(n34706), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4350), .I3(GND_net), .O(n34707));   // verilog/motorControl.v(31[38:63])
    defparam i28533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_4347), .I3(GND_net), 
            .O(n12_adj_4620));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i28068_2_lut (.I0(n33_adj_4347), .I1(n15_adj_4366), .I2(GND_net), 
            .I3(GND_net), .O(n34240));
    defparam i28068_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4392), .I3(GND_net), 
            .O(n10_adj_4621));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n25751), .I0(GND_net), .I1(n1_adj_4633[4]), 
            .CO(n25752));
    SB_CARRY add_12_6 (.CI(n25617), .I0(n106[4]), .I1(n155[4]), .CO(n25618));
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n25616), 
            .O(duty_23__N_3563[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4620), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4346), .I3(GND_net), 
            .O(n30_adj_4622));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i28078_4_lut (.I0(n33_adj_4347), .I1(n31_adj_4348), .I2(n29_adj_4350), 
            .I3(n34254), .O(n34250));
    defparam i28078_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5065_13 (.CI(n27020), .I0(n9454[10]), .I1(n904_adj_4408), 
            .CO(n27021));
    SB_LUT4 add_5065_13_lut (.I0(GND_net), .I1(n9454[10]), .I2(n904_adj_4408), 
            .I3(n27020), .O(n9438[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_14 (.CI(n27021), .I0(n9454[11]), .I1(n977_adj_4601), 
            .CO(n27022));
    SB_LUT4 i28675_4_lut (.I0(n30_adj_4622), .I1(n10_adj_4621), .I2(n35_adj_4346), 
            .I3(n34240), .O(n34849));   // verilog/motorControl.v(31[38:63])
    defparam i28675_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4601));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4598));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28336_3_lut (.I0(n34707), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_4348), .I3(GND_net), .O(n34510));   // verilog/motorControl.v(31[38:63])
    defparam i28336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28727_4_lut (.I0(n34510), .I1(n34849), .I2(n35_adj_4346), 
            .I3(n34250), .O(n34901));   // verilog/motorControl.v(31[38:63])
    defparam i28727_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4596));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4595));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4593));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4592));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4590));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28728_3_lut (.I0(n34901), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_4345), .I3(GND_net), .O(n34902));   // verilog/motorControl.v(31[38:63])
    defparam i28728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28700_3_lut (.I0(n34902), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4333), .I3(GND_net), .O(n34874));   // verilog/motorControl.v(31[38:63])
    defparam i28700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4589));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4419), .I3(GND_net), 
            .O(n6_adj_4623));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4587));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28534_3_lut (.I0(n6_adj_4623), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4353), .I3(GND_net), .O(n34708));   // verilog/motorControl.v(31[38:63])
    defparam i28534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28535_3_lut (.I0(n34708), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4352), .I3(GND_net), .O(n34709));   // verilog/motorControl.v(31[38:63])
    defparam i28535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28059_4_lut (.I0(n43_adj_4320), .I1(n25_adj_4351), .I2(n23_adj_4352), 
            .I3(n34260), .O(n34231));
    defparam i28059_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28486_4_lut (.I0(n24_adj_4609), .I1(n8_adj_4607), .I2(n45_adj_4319), 
            .I3(n34229), .O(n34660));   // verilog/motorControl.v(31[38:63])
    defparam i28486_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4584));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28334_3_lut (.I0(n34709), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4351), .I3(GND_net), .O(n34508));   // verilog/motorControl.v(31[38:63])
    defparam i28334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4583));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28061_4_lut (.I0(n43_adj_4320), .I1(n41_adj_4331), .I2(n39_adj_4333), 
            .I3(n34863), .O(n34233));
    defparam i28061_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i28638_4_lut (.I0(n34508), .I1(n34660), .I2(n45_adj_4319), 
            .I3(n34231), .O(n34812));   // verilog/motorControl.v(31[38:63])
    defparam i28638_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4582));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28342_3_lut (.I0(n34874), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4331), .I3(GND_net), .O(n34516));   // verilog/motorControl.v(31[38:63])
    defparam i28342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28687_4_lut (.I0(n34516), .I1(n34812), .I2(n45_adj_4319), 
            .I3(n34233), .O(n34861));   // verilog/motorControl.v(31[38:63])
    defparam i28687_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4581));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4624));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4580));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4579));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4633[3]), 
            .I3(n25750), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28540_3_lut (.I0(n4_adj_4624), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n34714));   // verilog/motorControl.v(31[10:34])
    defparam i28540_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28541_3_lut (.I0(n34714), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n34715));   // verilog/motorControl.v(31[10:34])
    defparam i28541_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_12_5 (.CI(n25616), .I0(n106[3]), .I1(n155[3]), .CO(n25617));
    SB_LUT4 i28118_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n36218), 
            .I2(IntegralLimit[16]), .I3(n34568), .O(n34290));
    defparam i28118_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i28673_4_lut (.I0(n30_adj_4615), .I1(n10_adj_4614), .I2(n36241), 
            .I3(n34288), .O(n34847));   // verilog/motorControl.v(31[10:34])
    defparam i28673_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i28326_3_lut (.I0(n34715), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n34500));   // verilog/motorControl.v(31[10:34])
    defparam i28326_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28725_4_lut (.I0(n34500), .I1(n34847), .I2(n36241), .I3(n34290), 
            .O(n34899));   // verilog/motorControl.v(31[10:34])
    defparam i28725_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28726_3_lut (.I0(n34899), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n34900));   // verilog/motorControl.v(31[10:34])
    defparam i28726_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4578));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28704_3_lut (.I0(n34900), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n34878));   // verilog/motorControl.v(31[10:34])
    defparam i28704_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28107_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n36209), 
            .I2(IntegralLimit[21]), .I3(n34891), .O(n34279));
    defparam i28107_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4577));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4576));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28636_4_lut (.I0(n34498), .I1(n34658), .I2(n36206), .I3(n34277), 
            .O(n34810));   // verilog/motorControl.v(31[10:34])
    defparam i28636_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4575));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28332_3_lut (.I0(n34878), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n34506));   // verilog/motorControl.v(31[10:34])
    defparam i28332_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i28688_3_lut (.I0(n34861), .I1(\PID_CONTROLLER.integral_23__N_3514 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3513 ));   // verilog/motorControl.v(31[38:63])
    defparam i28688_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4574));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4573));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28685_4_lut (.I0(n34506), .I1(n34810), .I2(n36206), .I3(n34279), 
            .O(n34859));   // verilog/motorControl.v(31[10:34])
    defparam i28685_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_831_4_lut  (.I0(n34859), .I1(\PID_CONTROLLER.integral_23__N_3513 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3511 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_831_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4572));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4571));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4570));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4569));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4568));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4567));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4566));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4565));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4563));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4561));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4559));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4558));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4556));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4555));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4553));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4552));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4550));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4549));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4547));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4546));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4543));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4541));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4540));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4538));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4537));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4534));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17837_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3511 ), 
            .I2(GND_net), .I3(GND_net), .O(n3005[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i17837_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4532));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4531));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4398));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4529));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4394));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4528));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4526));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4389));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4525));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4383));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4382));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4523));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4520));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4519));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4517));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4516));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4514));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4513));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1483 (.I0(n6_adj_4508), .I1(\Ki[4] ), .I2(n9553[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [18]), .O(n9546[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1483.LUT_INIT = 16'h965a;
    SB_LUT4 i20912_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3463 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [21]), .O(n9564[0]));   // verilog/motorControl.v(34[25:36])
    defparam i20912_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1484 (.I0(n4_adj_4510), .I1(\Ki[3] ), .I2(n9559[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [19]), .O(n9553[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1484.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1485 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3463 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [20]), .O(n12_adj_4625));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1485.LUT_INIT = 16'h9c50;
    SB_LUT4 i20848_4_lut (.I0(n9553[2]), .I1(\Ki[4] ), .I2(n6_adj_4508), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [18]), .O(n8_adj_4626));   // verilog/motorControl.v(34[25:36])
    defparam i20848_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1486 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3463 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [21]), .O(n11_adj_4627));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1486.LUT_INIT = 16'h6ca0;
    SB_LUT4 i20879_4_lut (.I0(n9559[1]), .I1(\Ki[3] ), .I2(n4_adj_4510), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [19]), .O(n6_adj_4628));   // verilog/motorControl.v(34[25:36])
    defparam i20879_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i20914_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3463 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [21]), .O(n25489));   // verilog/motorControl.v(34[25:36])
    defparam i20914_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1487 (.I0(n6_adj_4628), .I1(n11_adj_4627), .I2(n8_adj_4626), 
            .I3(n12_adj_4625), .O(n18_adj_4629));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1488 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3463 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3463 [22]), .O(n13_adj_4630));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1488.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1489 (.I0(n13_adj_4630), .I1(n18_adj_4629), .I2(n25489), 
            .I3(n4_adj_4511), .O(n32845));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4365));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4364));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4632[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4361));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4360));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4359));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4358));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4357));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4355));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4215));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20780_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n25332), 
            .I3(n9267[0]), .O(n4_adj_4499));   // verilog/motorControl.v(34[16:22])
    defparam i20780_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1490 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n9267[0]), 
            .I3(n25332), .O(n9262[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1490.LUT_INIT = 16'h8778;
    SB_LUT4 i20769_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n25332));   // verilog/motorControl.v(34[16:22])
    defparam i20769_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20767_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n9262[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20767_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20749_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n25298), 
            .I3(n9262[0]), .O(n4_adj_4492));   // verilog/motorControl.v(34[16:22])
    defparam i20749_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n9262[0]), 
            .I3(n25298), .O(n9256[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h8778;
    SB_LUT4 i20736_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n9256[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20736_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20738_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n25298));   // verilog/motorControl.v(34[16:22])
    defparam i20738_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20718_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4631), 
            .I3(n9256[1]), .O(n6_adj_4491));   // verilog/motorControl.v(34[16:22])
    defparam i20718_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1492 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n9256[1]), 
            .I3(n4_adj_4631), .O(n9249[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1492.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1493 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n9256[0]), 
            .I3(n25255), .O(n9249[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1493.LUT_INIT = 16'h8778;
    SB_LUT4 i20710_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n25255), 
            .I3(n9256[0]), .O(n4_adj_4631));   // verilog/motorControl.v(34[16:22])
    defparam i20710_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20699_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n25255));   // verilog/motorControl.v(34[16:22])
    defparam i20699_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20697_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n9249[0]));   // verilog/motorControl.v(34[16:22])
    defparam i20697_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4356));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3463 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, clk32MHz, 
            data_o, ENCODER1_A_c_1, reg_B, n33025, VCC_net, ENCODER1_B_c_0, 
            n18059, n18544) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    input ENCODER1_A_c_1;
    output [1:0]reg_B;
    output n33025;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n18059;
    input n18544;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2856;
    
    wire n2833, n25828, count_enable, B_delayed, A_delayed, n25829, 
        n25827, n25826, n25825, n25824, n25823, n25822, n25821, 
        n25820, n25819, n25818, n25817, n25816, n25815, n25814, 
        n25813, n25812, n25811, n25810, count_direction, n25809, 
        n25832, n25831, n25830;
    
    SB_LUT4 add_658_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2833), 
            .I3(n25828), .O(n2856[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_658_21 (.CI(n25828), .I0(encoder1_position[19]), .I1(n2833), 
            .CO(n25829));
    SB_LUT4 add_658_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2833), 
            .I3(n25827), .O(n2856[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_20 (.CI(n25827), .I0(encoder1_position[18]), .I1(n2833), 
            .CO(n25828));
    SB_LUT4 add_658_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2833), 
            .I3(n25826), .O(n2856[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_19 (.CI(n25826), .I0(encoder1_position[17]), .I1(n2833), 
            .CO(n25827));
    SB_LUT4 add_658_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2833), 
            .I3(n25825), .O(n2856[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[23]));   // quad.v(35[10] 41[6])
    SB_CARRY add_658_18 (.CI(n25825), .I0(encoder1_position[16]), .I1(n2833), 
            .CO(n25826));
    SB_LUT4 add_658_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2833), 
            .I3(n25824), .O(n2856[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_17 (.CI(n25824), .I0(encoder1_position[15]), .I1(n2833), 
            .CO(n25825));
    SB_LUT4 add_658_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2833), 
            .I3(n25823), .O(n2856[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_16 (.CI(n25823), .I0(encoder1_position[14]), .I1(n2833), 
            .CO(n25824));
    SB_LUT4 add_658_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2833), 
            .I3(n25822), .O(n2856[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_15 (.CI(n25822), .I0(encoder1_position[13]), .I1(n2833), 
            .CO(n25823));
    SB_LUT4 add_658_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2833), 
            .I3(n25821), .O(n2856[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_14 (.CI(n25821), .I0(encoder1_position[12]), .I1(n2833), 
            .CO(n25822));
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[22]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_658_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2833), 
            .I3(n25820), .O(n2856[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_13 (.CI(n25820), .I0(encoder1_position[11]), .I1(n2833), 
            .CO(n25821));
    SB_LUT4 add_658_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2833), 
            .I3(n25819), .O(n2856[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_12 (.CI(n25819), .I0(encoder1_position[10]), .I1(n2833), 
            .CO(n25820));
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2856[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_658_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2833), 
            .I3(n25818), .O(n2856[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_11 (.CI(n25818), .I0(encoder1_position[9]), .I1(n2833), 
            .CO(n25819));
    SB_LUT4 add_658_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2833), 
            .I3(n25817), .O(n2856[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_10 (.CI(n25817), .I0(encoder1_position[8]), .I1(n2833), 
            .CO(n25818));
    SB_LUT4 add_658_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2833), 
            .I3(n25816), .O(n2856[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_9 (.CI(n25816), .I0(encoder1_position[7]), .I1(n2833), 
            .CO(n25817));
    SB_LUT4 add_658_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2833), 
            .I3(n25815), .O(n2856[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_8 (.CI(n25815), .I0(encoder1_position[6]), .I1(n2833), 
            .CO(n25816));
    SB_LUT4 add_658_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2833), 
            .I3(n25814), .O(n2856[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_7 (.CI(n25814), .I0(encoder1_position[5]), .I1(n2833), 
            .CO(n25815));
    SB_LUT4 add_658_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2833), 
            .I3(n25813), .O(n2856[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_6 (.CI(n25813), .I0(encoder1_position[4]), .I1(n2833), 
            .CO(n25814));
    SB_LUT4 add_658_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2833), 
            .I3(n25812), .O(n2856[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_5 (.CI(n25812), .I0(encoder1_position[3]), .I1(n2833), 
            .CO(n25813));
    SB_LUT4 add_658_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2833), 
            .I3(n25811), .O(n2856[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_4 (.CI(n25811), .I0(encoder1_position[2]), .I1(n2833), 
            .CO(n25812));
    SB_LUT4 add_658_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2833), 
            .I3(n25810), .O(n2856[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_3 (.CI(n25810), .I0(encoder1_position[1]), .I1(n2833), 
            .CO(n25811));
    SB_LUT4 add_658_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n25809), .O(n2856[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_2 (.CI(n25809), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n25810));
    SB_CARRY add_658_1 (.CI(GND_net), .I0(n2833), .I1(n2833), .CO(n25809));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1105_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2833));   // quad.v(37[5] 40[8])
    defparam i1105_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_658_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2833), 
            .I3(n25832), .O(n2856[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_658_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2833), 
            .I3(n25831), .O(n2856[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_24 (.CI(n25831), .I0(encoder1_position[22]), .I1(n2833), 
            .CO(n25832));
    SB_LUT4 add_658_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2833), 
            .I3(n25830), .O(n2856[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_23 (.CI(n25830), .I0(encoder1_position[21]), .I1(n2833), 
            .CO(n25831));
    SB_LUT4 add_658_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2833), 
            .I3(n25829), .O(n2856[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_658_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_658_22 (.CI(n25829), .I0(encoder1_position[20]), .I1(n2833), 
            .CO(n25830));
    \grp_debouncer(2,100)  debounce (.ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .GND_net(GND_net), .n33025(n33025), .VCC_net(VCC_net), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n18059(n18059), .data_o({data_o}), 
            .n18544(n18544));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (ENCODER1_A_c_1, clk32MHz, reg_B, GND_net, 
            n33025, VCC_net, ENCODER1_B_c_0, n18059, data_o, n18544);
    input ENCODER1_A_c_1;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n33025;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n18059;
    output [1:0]data_o;
    input n18544;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [6:0]n33;
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n26334, n12, n26333, n2, cnt_next_6__N_3647, n26332, n26331, 
        n26330, n26329;
    
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1468_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n26334), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 cnt_reg_1468_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n26333), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n33025));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n33025), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_CARRY cnt_reg_1468_add_4_7 (.CI(n26333), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n26334));
    SB_LUT4 cnt_reg_1468_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n26332), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1468_add_4_6 (.CI(n26332), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n26333));
    SB_LUT4 cnt_reg_1468_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n26331), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1468_add_4_5 (.CI(n26331), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n26332));
    SB_LUT4 cnt_reg_1468_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n26330), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1468_add_4_4 (.CI(n26330), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n26331));
    SB_LUT4 cnt_reg_1468_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n26329), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1468_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1468_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1468_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n26329));
    SB_CARRY cnt_reg_1468_add_4_3 (.CI(n26329), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n26330));
    SB_DFFSR cnt_reg_1468__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18059));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18544));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1468__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1468__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1468__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1468__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1468__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1468__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3647));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (\state[2] , \state[0] , \state[3] , GND_net, n21828, 
            n21898, n4604, n21826, CLK_c, scl_enable, \state_7__N_3815[0] , 
            sda_enable, VCC_net, n5019, n34058, \state_7__N_3831[3] , 
            n10, n5, n882, n8, n11) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[2] ;
    output \state[0] ;
    output \state[3] ;
    input GND_net;
    output n21828;
    output n21898;
    output n4604;
    output n21826;
    input CLK_c;
    output scl_enable;
    output \state_7__N_3815[0] ;
    output sda_enable;
    input VCC_net;
    input n5019;
    output n34058;
    output \state_7__N_3831[3] ;
    input n10;
    input n5;
    output [0:0]n882;
    input n8;
    output n11;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    i2c_controller i2c (.\state[2] (\state[2] ), .\state[0] (\state[0] ), 
            .\state[3] (\state[3] ), .GND_net(GND_net), .n21828(n21828), 
            .n21898(n21898), .n4604(n4604), .n21826(n21826), .CLK_c(CLK_c), 
            .scl_enable(scl_enable), .\state_7__N_3815[0] (\state_7__N_3815[0] ), 
            .sda_enable(sda_enable), .VCC_net(VCC_net), .n5019(n5019), 
            .n34058(n34058), .\state_7__N_3831[3] (\state_7__N_3831[3] ), 
            .n10(n10), .n5(n5), .n882({n882}), .n8(n8), .n11(n11)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(59[16] 72[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state[2] , \state[0] , \state[3] , GND_net, 
            n21828, n21898, n4604, n21826, CLK_c, scl_enable, \state_7__N_3815[0] , 
            sda_enable, VCC_net, n5019, n34058, \state_7__N_3831[3] , 
            n10, n5, n882, n8, n11) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[2] ;
    output \state[0] ;
    output \state[3] ;
    input GND_net;
    output n21828;
    output n21898;
    output n4604;
    output n21826;
    input CLK_c;
    output scl_enable;
    output \state_7__N_3815[0] ;
    output sda_enable;
    input VCC_net;
    input n5019;
    output n34058;
    output \state_7__N_3831[3] ;
    input n10;
    input n5;
    output [0:0]n882;
    input n8;
    output n11;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(40[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n883;
    
    wire n17861;
    wire [7:0]counter;   // verilog/i2c_controller.v(35[12:19])
    
    wire n18019;
    wire [7:0]state;   // verilog/i2c_controller.v(32[12:17])
    
    wire n33991, n11_c, n34096, n7, n33, n37, n17958, n34, n39, 
        counter2_7__N_3802, n10024;
    wire [7:0]counter2;   // verilog/i2c_controller.v(36[12:20])
    
    wire n6, i2c_clk_N_3907, n15, n22761, n10_c, n17717, n4597, 
        n11_adj_4207, n34088, n30257, scl_enable_N_3908, enable_slow_N_3918, 
        n9882, n4896, n30123, sda_out;
    wire [4:0]n25;
    
    wire n26338, n26337, n25808, n25807, n26336, n25806, n25805, 
        n25804, n26335, n25803, n25802, n10_adj_4208, n14, n31270, 
        n22072, n32894, n22630;
    
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n17861), .D(n883[5]), 
            .R(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i28213_4_lut (.I0(counter[1]), .I1(state[1]), .I2(counter[0]), 
            .I3(counter[2]), .O(n33991));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam i28213_4_lut.LUT_INIT = 16'hc004;
    SB_LUT4 i28149_4_lut (.I0(n33991), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11_c), .O(n34096));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam i28149_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 i1_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(state[1]), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n17958));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_1474 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_1474.LUT_INIT = 16'heeee;
    SB_LUT4 i17258_2_lut_4_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n21828));
    defparam i17258_2_lut_4_lut_4_lut.LUT_INIT = 16'hfdfb;
    SB_LUT4 i5525_2_lut (.I0(i2c_clk), .I1(counter2_7__N_3802), .I2(GND_net), 
            .I3(GND_net), .O(n10024));   // verilog/i2c_controller.v(68[8:33])
    defparam i5525_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17327_2_lut (.I0(state[1]), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n21898));
    defparam i17327_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1475 (.I0(counter2[0]), .I1(counter2[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_1475.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[2]), .I2(counter2[1]), 
            .I3(n6), .O(counter2_7__N_3802));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1476 (.I0(i2c_clk), .I1(counter2_7__N_3802), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_3907));
    defparam i1_2_lut_adj_1476.LUT_INIT = 16'h6666;
    SB_LUT4 i28988_3_lut (.I0(n4604), .I1(n15), .I2(n21828), .I3(GND_net), 
            .O(n22761));
    defparam i28988_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 state_7__I_0_144_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // verilog/i2c_controller.v(137[5:14])
    defparam state_7__I_0_144_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i28775_4_lut (.I0(n17717), .I1(n4597), .I2(n11_adj_4207), 
            .I3(n21826), .O(n4604));
    defparam i28775_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut (.I0(state[1]), .I1(n7), .I2(n34088), .I3(\state[0] ), 
            .O(n30257));   // verilog/i2c_controller.v(90[4] 154[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n17861), .D(n883[4]), 
            .R(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n17861), .D(n883[3]), 
            .R(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n17861), .D(n883[2]), 
            .S(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_3907));   // verilog/i2c_controller.v(57[9] 69[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_3908));   // verilog/i2c_controller.v(74[12] 80[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_3815[0] ), .C(CLK_c), .E(n10024), 
            .D(enable_slow_N_3918));   // verilog/i2c_controller.v(57[9] 69[5])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n4896), 
            .D(n9882), .S(n17958));   // verilog/i2c_controller.v(162[12] 197[6])
    SB_DFFNE sda_out_133 (.Q(sda_out), .C(i2c_clk), .E(n30123), .D(n34096));   // verilog/i2c_controller.v(162[12] 197[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n17861), .D(n883[0]), 
            .S(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 counter2_1469_1470_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n26338), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1469_1470_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1469_1470_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n26337), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1469_1470_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_89_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n25808), .O(n883[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1469_1470_add_4_5 (.CI(n26337), .I0(GND_net), .I1(counter2[3]), 
            .CO(n26338));
    SB_LUT4 sub_89_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n25807), .O(n883[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_8 (.CI(n25807), .I0(counter[6]), .I1(VCC_net), 
            .CO(n25808));
    SB_LUT4 counter2_1469_1470_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n26336), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1469_1470_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1469_1470_add_4_4 (.CI(n26336), .I0(GND_net), .I1(counter2[2]), 
            .CO(n26337));
    SB_LUT4 sub_89_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n25806), .O(n883[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_7 (.CI(n25806), .I0(counter[5]), .I1(VCC_net), 
            .CO(n25807));
    SB_LUT4 sub_89_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n25805), .O(n883[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_6 (.CI(n25805), .I0(counter[4]), .I1(VCC_net), 
            .CO(n25806));
    SB_LUT4 sub_89_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n25804), .O(n883[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_5 (.CI(n25804), .I0(counter[3]), .I1(VCC_net), 
            .CO(n25805));
    SB_LUT4 counter2_1469_1470_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n26335), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1469_1470_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_89_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n25803), .O(n883[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1469_1470_add_4_3 (.CI(n26335), .I0(GND_net), .I1(counter2[1]), 
            .CO(n26336));
    SB_CARRY sub_89_add_2_4 (.CI(n25803), .I0(counter[2]), .I1(VCC_net), 
            .CO(n25804));
    SB_LUT4 sub_89_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n25802), .O(n883[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_3 (.CI(n25802), .I0(counter[1]), .I1(VCC_net), 
            .CO(n25803));
    SB_LUT4 sub_89_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n883[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_89_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_89_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n25802));
    SB_LUT4 counter2_1469_1470_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1469_1470_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1469_1470_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n26335));
    SB_DFFSR counter2_1469_1470__i1 (.Q(counter2[0]), .C(CLK_c), .D(n25[0]), 
            .R(counter2_7__N_3802));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n17861), .D(n883[1]), 
            .S(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i2_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4208));   // verilog/i2c_controller.v(107[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(counter[7]), .I1(counter[4]), .I2(counter[5]), 
            .I3(counter[6]), .O(n14));   // verilog/i2c_controller.v(107[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(counter[0]), .I1(n14), .I2(n10_adj_4208), .I3(counter[3]), 
            .O(n4597));   // verilog/i2c_controller.v(107[10:22])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n4597), .I1(n31270), .I2(n5019), .I3(n37), 
            .O(n17861));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 equal_86_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(75[27:43])
    defparam equal_86_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(state[1]), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i28167_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(n10_c), 
            .I3(n22072), .O(n34058));   // verilog/i2c_controller.v(137[5:14])
    defparam i28167_3_lut_4_lut.LUT_INIT = 16'hfb00;
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n4604), .D(n30257), 
            .S(n32894));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state_7__N_3831[3] ), 
            .I3(n10), .O(n22072));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n4604), .D(n22630), 
            .S(n22761));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n17717));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4207));   // verilog/i2c_controller.v(137[5:14])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i25061_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n31270), .O(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i25061_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i25111_2_lut_3_lut (.I0(sda_out), .I1(sda_enable), .I2(n15), 
            .I3(GND_net), .O(n31270));
    defparam i25111_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(state[1]), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1514;
    SB_DFFE state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(VCC_net), .D(n5));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i17353_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(n882[0]));   // verilog/i2c_controller.v(44[19:55])
    defparam i17353_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1707_2_lut (.I0(sda_out), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(\state_7__N_3831[3] ));   // verilog/i2c_controller.v(45[9:16])
    defparam i1707_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFSR counter2_1469_1470__i2 (.Q(counter2[1]), .C(CLK_c), .D(n25[1]), 
            .R(counter2_7__N_3802));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1469_1470__i3 (.Q(counter2[2]), .C(CLK_c), .D(n25[2]), 
            .R(counter2_7__N_3802));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1469_1470__i4 (.Q(counter2[3]), .C(CLK_c), .D(n25[3]), 
            .R(counter2_7__N_3802));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1469_1470__i5 (.Q(counter2[4]), .C(CLK_c), .D(n25[4]), 
            .R(counter2_7__N_3802));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n17861), .D(n883[7]), 
            .R(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n17861), .D(n883[6]), 
            .R(n18019));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i28804_4_lut_4_lut (.I0(state[1]), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n30123));
    defparam i28804_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i28093_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(sda_out), 
            .I3(sda_enable), .O(n34088));   // verilog/i2c_controller.v(90[4] 154[11])
    defparam i28093_3_lut_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i28991_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(state[1]), 
            .I3(n4604), .O(n32894));
    defparam i28991_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i17813_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n21826));
    defparam i17813_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i18271_3_lut_4_lut (.I0(n15), .I1(state[1]), .I2(\state[0] ), 
            .I3(\state[2] ), .O(scl_enable_N_3908));
    defparam i18271_3_lut_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i13349_1_lut_2_lut (.I0(i2c_clk), .I1(counter2_7__N_3802), .I2(GND_net), 
            .I3(GND_net), .O(enable_slow_N_3918));
    defparam i13349_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state[3] ), 
            .I3(GND_net), .O(n11_c));
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i2_3_lut_4_lut_adj_1477 (.I0(\state[0] ), .I1(state[1]), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(75[27:43])
    defparam i2_3_lut_4_lut_adj_1477.LUT_INIT = 16'hfdff;
    SB_LUT4 i28791_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(n10_c), 
            .I3(n22072), .O(n22630));   // verilog/i2c_controller.v(75[27:43])
    defparam i28791_3_lut_4_lut.LUT_INIT = 16'h02ff;
    SB_LUT4 i28806_4_lut_4_lut (.I0(\state[2] ), .I1(n11_c), .I2(state[1]), 
            .I3(n39), .O(n4896));
    defparam i28806_4_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i28815_2_lut_3_lut (.I0(\state[2] ), .I1(n11_c), .I2(\state[0] ), 
            .I3(GND_net), .O(n9882));
    defparam i28815_2_lut_3_lut.LUT_INIT = 16'h0404;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n34753, VCC_net, INHA_c, clk32MHz, n16458, GND_net, 
            pwm_counter, n16456) /* synthesis syn_module_defined=1 */ ;
    input n34753;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n16458;
    input GND_net;
    output [31:0]pwm_counter;
    input n16456;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n133;
    
    wire n26282, n26281, n26280, n26279, n26278, n26277, n26276, 
        n26275, n26274, n26273, n26272, n26271, n26270, n26269, 
        n26268, n26267, n26266, n26265, n26264, n26263, n26262, 
        n26261, n26260, n26259, n26258, n26257, n26256, n26255, 
        n26254, n26253, n26252, n32061, n18, n24, n22, n26, 
        n21, pwm_counter_31__N_602;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n34753), 
            .R(n16458));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_1462_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n26282), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1462_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n26281), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_32 (.CI(n26281), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n26282));
    SB_LUT4 pwm_counter_1462_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n26280), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_31 (.CI(n26280), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n26281));
    SB_LUT4 pwm_counter_1462_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n26279), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_30 (.CI(n26279), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n26280));
    SB_LUT4 pwm_counter_1462_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n26278), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_29 (.CI(n26278), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n26279));
    SB_LUT4 pwm_counter_1462_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n26277), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_28 (.CI(n26277), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n26278));
    SB_LUT4 pwm_counter_1462_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n26276), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_27 (.CI(n26276), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n26277));
    SB_LUT4 pwm_counter_1462_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n26275), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_26 (.CI(n26275), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n26276));
    SB_LUT4 pwm_counter_1462_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n26274), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_25 (.CI(n26274), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n26275));
    SB_LUT4 pwm_counter_1462_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n26273), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_24 (.CI(n26273), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n26274));
    SB_LUT4 pwm_counter_1462_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n26272), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_23 (.CI(n26272), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n26273));
    SB_LUT4 pwm_counter_1462_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n26271), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_22 (.CI(n26271), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n26272));
    SB_LUT4 pwm_counter_1462_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n26270), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_21 (.CI(n26270), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n26271));
    SB_LUT4 pwm_counter_1462_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n26269), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_20 (.CI(n26269), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n26270));
    SB_LUT4 pwm_counter_1462_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n26268), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_19 (.CI(n26268), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n26269));
    SB_LUT4 pwm_counter_1462_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n26267), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_18 (.CI(n26267), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n26268));
    SB_LUT4 pwm_counter_1462_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n26266), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_17 (.CI(n26266), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n26267));
    SB_LUT4 pwm_counter_1462_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n26265), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_16 (.CI(n26265), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n26266));
    SB_LUT4 pwm_counter_1462_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n26264), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_15 (.CI(n26264), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n26265));
    SB_LUT4 pwm_counter_1462_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n26263), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_14 (.CI(n26263), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n26264));
    SB_LUT4 pwm_counter_1462_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n26262), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_13 (.CI(n26262), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n26263));
    SB_LUT4 pwm_counter_1462_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n26261), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_12 (.CI(n26261), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n26262));
    SB_LUT4 pwm_counter_1462_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n26260), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_11 (.CI(n26260), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n26261));
    SB_LUT4 pwm_counter_1462_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n26259), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_10 (.CI(n26259), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n26260));
    SB_LUT4 pwm_counter_1462_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n26258), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_9 (.CI(n26258), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n26259));
    SB_LUT4 pwm_counter_1462_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n26257), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_8 (.CI(n26257), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n26258));
    SB_LUT4 pwm_counter_1462_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n26256), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_7 (.CI(n26256), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n26257));
    SB_LUT4 pwm_counter_1462_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n26255), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_6 (.CI(n26255), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n26256));
    SB_LUT4 pwm_counter_1462_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n26254), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_5 (.CI(n26254), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n26255));
    SB_LUT4 pwm_counter_1462_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n26253), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_4 (.CI(n26253), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n26254));
    SB_LUT4 pwm_counter_1462_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n26252), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_3 (.CI(n26252), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n26253));
    SB_LUT4 pwm_counter_1462_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1462_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1462_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n26252));
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n32061));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n32061), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(pwm_counter[18]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[21]), .I1(n16456), .I2(pwm_counter[16]), 
            .I3(pwm_counter[12]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(pwm_counter[15]), .I1(n24), .I2(n18), .I3(pwm_counter[19]), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[11]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17464_4_lut (.I0(n21), .I1(pwm_counter[31]), .I2(n26), .I3(n22), 
            .O(pwm_counter_31__N_602));   // verilog/pwm.v(18[8:40])
    defparam i17464_4_lut.LUT_INIT = 16'h3332;
    SB_DFFSR pwm_counter_1462__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1462__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_602));   // verilog/pwm.v(17[20:33])
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, GND_net, \data_out_frame[14] , \data_out_frame[13] , 
            \data_out_frame[12] , \data_out_frame[18] , \data_out_frame[19] , 
            \data_out_frame[15] , \data_out_frame[17] , n30471, \data_out_frame[16] , 
            \data_out_frame[9] , \data_out_frame[11] , \data_out_frame[5] , 
            \data_out_frame[7] , \data_out_frame[8] , \data_out_frame[6] , 
            \data_out_frame[10] , \data_out_frame[5][7] , \FRAME_MATCHER.state[0] , 
            \data_out_frame[5][6] , n30475, \data_out_frame[23] , \data_out_frame[25] , 
            \FRAME_MATCHER.state[3] , n22632, \data_in_frame[1] , \data_in_frame[2] , 
            \data_in_frame[1][6] , \data_in_frame[1][7] , n16613, n4922, 
            n122, n16606, n3303, n63, n5, n36350, \data_in_frame[3] , 
            n63_adj_3, n2696, n4452, n16621, n13810, n771, n9711, 
            n123, \FRAME_MATCHER.state_31__N_2579[1] , \data_in[0] , \data_in[1] , 
            \data_in[2] , \data_in[3] , rx_data, \data_in_frame[11] , 
            \data_in_frame[9] , \data_in_frame[4] , \data_in_frame[13] , 
            \data_in_frame[21] , control_mode, n32040, \data_in_frame[12] , 
            \data_in_frame[10] , \data_in_frame[8] , rx_data_ready, setpoint, 
            \data_in_frame[6] , \data_in_frame[5] , \data_out_frame[20] , 
            n18102, n18101, n18100, n16614, n18099, n18098, \control_mode[6] , 
            \control_mode[7] , \control_mode[4] , \control_mode[5] , n15, 
            \state[2] , \state[3] , n10, n15_adj_4, tx_active, \data_out_frame[24] , 
            n18097, n18096, n18095, DE_c, n18091, n18090, n18089, 
            n18088, n18087, PWMLimit, n18086, n18085, n18084, n18083, 
            n18082, n18081, n18080, n18079, n18078, n18077, n18076, 
            n18075, n18074, n18073, n18072, n18071, n18070, n18069, 
            n18068, n18067, n18066, n18065, n35879, n35882, LED_c, 
            n32812, \state[0] , n5019, n18536, IntegralLimit, n18535, 
            n18534, n18533, n18532, n18531, n18530, n18529, n18528, 
            n18527, n18526, n18525, n18524, n18523, n18522, n18521, 
            n18520, n18519, n18518, n18517, n18516, n18515, n18514, 
            n18513, n18512, n18511, n18510, n18509, n18508, n18507, 
            n18506, n18505, n18504, n18503, n18502, n18501, n18500, 
            n18499, n18498, n18497, n18496, n18495, n18494, n18493, 
            n18492, n18491, n18490, n18489, n18485, n18484, n18483, 
            n18482, n18481, n18480, n18479, \Kp[1] , n18478, \Kp[2] , 
            n18477, \Kp[3] , n18476, \Kp[4] , n18475, \Kp[5] , n18474, 
            \Kp[6] , n18473, \Kp[7] , n18472, \Kp[8] , n18471, \Kp[9] , 
            n18470, \Kp[10] , n18469, \Kp[11] , n18468, \Kp[12] , 
            n18467, \Kp[13] , n18466, \Kp[14] , n18465, \Kp[15] , 
            n18464, \Ki[1] , n18463, \Ki[2] , n18462, \Ki[3] , n18461, 
            \Ki[4] , n18460, \Ki[5] , n18459, \Ki[6] , n18458, \Ki[7] , 
            n18457, \Ki[8] , n18456, \Ki[9] , n18455, \Ki[10] , 
            n18454, \Ki[11] , n18453, \Ki[12] , n18452, \Ki[13] , 
            n18451, \Ki[14] , n18450, \Ki[15] , n18447, n18446, 
            n18445, n18444, n18443, n18442, n18441, n18440, n18439, 
            n18438, n18437, n18436, n18435, n18434, n18433, n18432, 
            n18431, n18430, n18429, n18428, n18427, n18426, n18425, 
            n18424, n18423, n18422, n18421, n18420, n18419, n18418, 
            n18417, n18416, n18415, n18414, n18413, n18412, n18411, 
            n18410, n18409, n18408, n18407, n18406, n18405, n18404, 
            n18403, n18402, n18401, n18400, n18399, n18398, n18397, 
            n18396, n18395, n18394, n18393, n18392, n18391, n18390, 
            n18389, n18388, n18387, n18386, n18385, n18384, n18383, 
            n18382, n18381, n18380, n18379, n18378, n18377, n18376, 
            n18375, n18374, n18373, n18372, n18371, n18370, n18369, 
            n18368, n18367, n18366, n18365, n18364, n18363, n18362, 
            n18361, n18360, n18359, n18358, n18357, n18356, n18355, 
            n18354, n18353, n18352, n18351, n18350, n18349, n18348, 
            n29947, n18347, n18346, n18345, n18344, n18343, n18342, 
            n18341, n18055, n18340, n18339, n18338, n18337, n18336, 
            n18335, n18334, n18333, n18332, n18331, n18330, n18329, 
            n18328, n18327, n18326, n18325, n18324, n18323, n18317, 
            n18316, n18315, n18314, n18313, n18312, n18311, n18310, 
            n18309, n18308, n18307, n18306, n18305, n18304, n18303, 
            n18302, n18301, n18300, n18052, neopxl_color, n18051, 
            \Ki[0] , n18050, \Kp[0] , n18049, n18299, n18298, n18297, 
            n18296, n18295, n18294, n18293, n18040, n18292, n18291, 
            n18290, n18289, n18288, n18287, n18286, n18285, n18284, 
            n18283, n18282, n18281, n18280, n18279, n18278, n18277, 
            n18276, n18275, n18274, n18273, n18272, n18271, n18270, 
            n18230, n18229, n18228, n18227, n18226, n18225, n18224, 
            n18223, n18166, n18165, n18164, n18163, n18162, n18161, 
            n18160, n18159, n19, \motor_state_23__N_74[0] , \encoder0_position_scaled[0] , 
            motor_state, \motor_state_23__N_74[1] , \encoder0_position_scaled[1] , 
            \motor_state_23__N_74[2] , \encoder0_position_scaled[2] , \motor_state_23__N_74[3] , 
            \encoder0_position_scaled[3] , \motor_state_23__N_74[4] , \encoder0_position_scaled[4] , 
            \motor_state_23__N_74[5] , \encoder0_position_scaled[5] , \motor_state_23__N_74[6] , 
            \encoder0_position_scaled[6] , \motor_state_23__N_74[7] , \encoder0_position_scaled[7] , 
            \motor_state_23__N_74[8] , \encoder0_position_scaled[8] , \motor_state_23__N_74[9] , 
            \encoder0_position_scaled[9] , \motor_state_23__N_74[10] , \encoder0_position_scaled[10] , 
            \motor_state_23__N_74[11] , \encoder0_position_scaled[11] , 
            \motor_state_23__N_74[12] , \encoder0_position_scaled[12] , 
            \motor_state_23__N_74[13] , \encoder0_position_scaled[13] , 
            \motor_state_23__N_74[14] , \encoder0_position_scaled[14] , 
            \motor_state_23__N_74[15] , \encoder0_position_scaled[15] , 
            \motor_state_23__N_74[16] , \encoder0_position_scaled[16] , 
            \motor_state_23__N_74[17] , \encoder0_position_scaled[17] , 
            \motor_state_23__N_74[18] , \encoder0_position_scaled[18] , 
            \motor_state_23__N_74[19] , \encoder0_position_scaled[19] , 
            \motor_state_23__N_74[20] , \encoder0_position_scaled[20] , 
            \motor_state_23__N_74[21] , \encoder0_position_scaled[22] , 
            \motor_state_23__N_74[23] , \motor_state_23__N_74[22] , n13933, 
            n30466, VCC_net, n17831, n17982, r_SM_Main, \r_SM_Main_2__N_3404[1] , 
            tx_o, \r_Bit_Index[0] , n4, n18322, n18058, n35944, 
            n9799, tx_enable, n17825, n17980, \r_Bit_Index[0]_adj_5 , 
            n16549, n4_adj_6, r_Rx_Data, RX_N_2, n18488, n21943, 
            n4_adj_7, n4_adj_8, n16544, n18540, n18048, n18047, 
            n18046, n18045, n18044, n18043, n18042) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    input GND_net;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[17] ;
    output n30471;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[10] ;
    output \data_out_frame[5][7] ;
    output \FRAME_MATCHER.state[0] ;
    output \data_out_frame[5][6] ;
    output n30475;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[25] ;
    output \FRAME_MATCHER.state[3] ;
    output n22632;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output \data_in_frame[1][6] ;
    output \data_in_frame[1][7] ;
    output n16613;
    input n4922;
    output n122;
    output n16606;
    output n3303;
    output n63;
    output n5;
    output n36350;
    output [7:0]\data_in_frame[3] ;
    input n63_adj_3;
    output n2696;
    output n4452;
    output n16621;
    output n13810;
    output n771;
    output n9711;
    output n123;
    output \FRAME_MATCHER.state_31__N_2579[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[21] ;
    output [7:0]control_mode;
    output n32040;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[8] ;
    output rx_data_ready;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_out_frame[20] ;
    input n18102;
    input n18101;
    input n18100;
    output n16614;
    input n18099;
    input n18098;
    output \control_mode[6] ;
    output \control_mode[7] ;
    output \control_mode[4] ;
    output \control_mode[5] ;
    output n15;
    input \state[2] ;
    input \state[3] ;
    output n10;
    output n15_adj_4;
    output tx_active;
    output [7:0]\data_out_frame[24] ;
    input n18097;
    input n18096;
    input n18095;
    output DE_c;
    input n18091;
    input n18090;
    input n18089;
    input n18088;
    input n18087;
    output [23:0]PWMLimit;
    input n18086;
    input n18085;
    input n18084;
    input n18083;
    input n18082;
    input n18081;
    input n18080;
    input n18079;
    input n18078;
    input n18077;
    input n18076;
    input n18075;
    input n18074;
    input n18073;
    input n18072;
    input n18071;
    input n18070;
    input n18069;
    input n18068;
    input n18067;
    input n18066;
    input n18065;
    input n35879;
    input n35882;
    output LED_c;
    output n32812;
    input \state[0] ;
    output n5019;
    input n18536;
    output [23:0]IntegralLimit;
    input n18535;
    input n18534;
    input n18533;
    input n18532;
    input n18531;
    input n18530;
    input n18529;
    input n18528;
    input n18527;
    input n18526;
    input n18525;
    input n18524;
    input n18523;
    input n18522;
    input n18521;
    input n18520;
    input n18519;
    input n18518;
    input n18517;
    input n18516;
    input n18515;
    input n18514;
    input n18513;
    input n18512;
    input n18511;
    input n18510;
    input n18509;
    input n18508;
    input n18507;
    input n18506;
    input n18505;
    input n18504;
    input n18503;
    input n18502;
    input n18501;
    input n18500;
    input n18499;
    input n18498;
    input n18497;
    input n18496;
    input n18495;
    input n18494;
    input n18493;
    input n18492;
    input n18491;
    input n18490;
    input n18489;
    input n18485;
    input n18484;
    input n18483;
    input n18482;
    input n18481;
    input n18480;
    input n18479;
    output \Kp[1] ;
    input n18478;
    output \Kp[2] ;
    input n18477;
    output \Kp[3] ;
    input n18476;
    output \Kp[4] ;
    input n18475;
    output \Kp[5] ;
    input n18474;
    output \Kp[6] ;
    input n18473;
    output \Kp[7] ;
    input n18472;
    output \Kp[8] ;
    input n18471;
    output \Kp[9] ;
    input n18470;
    output \Kp[10] ;
    input n18469;
    output \Kp[11] ;
    input n18468;
    output \Kp[12] ;
    input n18467;
    output \Kp[13] ;
    input n18466;
    output \Kp[14] ;
    input n18465;
    output \Kp[15] ;
    input n18464;
    output \Ki[1] ;
    input n18463;
    output \Ki[2] ;
    input n18462;
    output \Ki[3] ;
    input n18461;
    output \Ki[4] ;
    input n18460;
    output \Ki[5] ;
    input n18459;
    output \Ki[6] ;
    input n18458;
    output \Ki[7] ;
    input n18457;
    output \Ki[8] ;
    input n18456;
    output \Ki[9] ;
    input n18455;
    output \Ki[10] ;
    input n18454;
    output \Ki[11] ;
    input n18453;
    output \Ki[12] ;
    input n18452;
    output \Ki[13] ;
    input n18451;
    output \Ki[14] ;
    input n18450;
    output \Ki[15] ;
    input n18447;
    input n18446;
    input n18445;
    input n18444;
    input n18443;
    input n18442;
    input n18441;
    input n18440;
    input n18439;
    input n18438;
    input n18437;
    input n18436;
    input n18435;
    input n18434;
    input n18433;
    input n18432;
    input n18431;
    input n18430;
    input n18429;
    input n18428;
    input n18427;
    input n18426;
    input n18425;
    input n18424;
    input n18423;
    input n18422;
    input n18421;
    input n18420;
    input n18419;
    input n18418;
    input n18417;
    input n18416;
    input n18415;
    input n18414;
    input n18413;
    input n18412;
    input n18411;
    input n18410;
    input n18409;
    input n18408;
    input n18407;
    input n18406;
    input n18405;
    input n18404;
    input n18403;
    input n18402;
    input n18401;
    input n18400;
    input n18399;
    input n18398;
    input n18397;
    input n18396;
    input n18395;
    input n18394;
    input n18393;
    input n18392;
    input n18391;
    input n18390;
    input n18389;
    input n18388;
    input n18387;
    input n18386;
    input n18385;
    input n18384;
    input n18383;
    input n18382;
    input n18381;
    input n18380;
    input n18379;
    input n18378;
    input n18377;
    input n18376;
    input n18375;
    input n18374;
    input n18373;
    input n18372;
    input n18371;
    input n18370;
    input n18369;
    input n18368;
    input n18367;
    input n18366;
    input n18365;
    input n18364;
    input n18363;
    input n18362;
    input n18361;
    input n18360;
    input n18359;
    input n18358;
    input n18357;
    input n18356;
    input n18355;
    input n18354;
    input n18353;
    input n18352;
    input n18351;
    input n18350;
    input n18349;
    input n18348;
    input n29947;
    input n18347;
    input n18346;
    input n18345;
    input n18344;
    input n18343;
    input n18342;
    input n18341;
    input n18055;
    input n18340;
    input n18339;
    input n18338;
    input n18337;
    input n18336;
    input n18335;
    input n18334;
    input n18333;
    input n18332;
    input n18331;
    input n18330;
    input n18329;
    input n18328;
    input n18327;
    input n18326;
    input n18325;
    input n18324;
    input n18323;
    input n18317;
    input n18316;
    input n18315;
    input n18314;
    input n18313;
    input n18312;
    input n18311;
    input n18310;
    input n18309;
    input n18308;
    input n18307;
    input n18306;
    input n18305;
    input n18304;
    input n18303;
    input n18302;
    input n18301;
    input n18300;
    input n18052;
    output [23:0]neopxl_color;
    input n18051;
    output \Ki[0] ;
    input n18050;
    output \Kp[0] ;
    input n18049;
    input n18299;
    input n18298;
    input n18297;
    input n18296;
    input n18295;
    input n18294;
    input n18293;
    input n18040;
    input n18292;
    input n18291;
    input n18290;
    input n18289;
    input n18288;
    input n18287;
    input n18286;
    input n18285;
    input n18284;
    input n18283;
    input n18282;
    input n18281;
    input n18280;
    input n18279;
    input n18278;
    input n18277;
    input n18276;
    input n18275;
    input n18274;
    input n18273;
    input n18272;
    input n18271;
    input n18270;
    input n18230;
    input n18229;
    input n18228;
    input n18227;
    input n18226;
    input n18225;
    input n18224;
    input n18223;
    input n18166;
    input n18165;
    input n18164;
    input n18163;
    input n18162;
    input n18161;
    input n18160;
    input n18159;
    output n19;
    input \motor_state_23__N_74[0] ;
    input \encoder0_position_scaled[0] ;
    output [23:0]motor_state;
    input \motor_state_23__N_74[1] ;
    input \encoder0_position_scaled[1] ;
    input \motor_state_23__N_74[2] ;
    input \encoder0_position_scaled[2] ;
    input \motor_state_23__N_74[3] ;
    input \encoder0_position_scaled[3] ;
    input \motor_state_23__N_74[4] ;
    input \encoder0_position_scaled[4] ;
    input \motor_state_23__N_74[5] ;
    input \encoder0_position_scaled[5] ;
    input \motor_state_23__N_74[6] ;
    input \encoder0_position_scaled[6] ;
    input \motor_state_23__N_74[7] ;
    input \encoder0_position_scaled[7] ;
    input \motor_state_23__N_74[8] ;
    input \encoder0_position_scaled[8] ;
    input \motor_state_23__N_74[9] ;
    input \encoder0_position_scaled[9] ;
    input \motor_state_23__N_74[10] ;
    input \encoder0_position_scaled[10] ;
    input \motor_state_23__N_74[11] ;
    input \encoder0_position_scaled[11] ;
    input \motor_state_23__N_74[12] ;
    input \encoder0_position_scaled[12] ;
    input \motor_state_23__N_74[13] ;
    input \encoder0_position_scaled[13] ;
    input \motor_state_23__N_74[14] ;
    input \encoder0_position_scaled[14] ;
    input \motor_state_23__N_74[15] ;
    input \encoder0_position_scaled[15] ;
    input \motor_state_23__N_74[16] ;
    input \encoder0_position_scaled[16] ;
    input \motor_state_23__N_74[17] ;
    input \encoder0_position_scaled[17] ;
    input \motor_state_23__N_74[18] ;
    input \encoder0_position_scaled[18] ;
    input \motor_state_23__N_74[19] ;
    input \encoder0_position_scaled[19] ;
    input \motor_state_23__N_74[20] ;
    input \encoder0_position_scaled[20] ;
    input \motor_state_23__N_74[21] ;
    input \encoder0_position_scaled[22] ;
    input \motor_state_23__N_74[23] ;
    input \motor_state_23__N_74[22] ;
    output n13933;
    output n30466;
    input VCC_net;
    output n17831;
    output n17982;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3404[1] ;
    output tx_o;
    output \r_Bit_Index[0] ;
    output n4;
    input n18322;
    input n18058;
    input n35944;
    output n9799;
    output tx_enable;
    output n17825;
    output n17980;
    output \r_Bit_Index[0]_adj_5 ;
    output n16549;
    output n4_adj_6;
    output r_Rx_Data;
    input RX_N_2;
    input n18488;
    output n21943;
    output n4_adj_7;
    output n4_adj_8;
    output n16544;
    input n18540;
    input n18048;
    input n18047;
    input n18046;
    input n18045;
    input n18044;
    input n18043;
    input n18042;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n30913, n20, n16, n30556, n31662, n18120;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n30852, n24, n28088, n28, n28125, n8, n16954, n17350, 
        n26, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n18119, n16878, n30502, n17336, n16702, n30524, n7, 
        n32089, n2112, n30949, n30703, n30493, n16666, n30714, 
        n31093, n28782, n28681, n6, n28740, n18118;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n30817, n27756, n28767, n30773, n30468, n31090, n30617, 
        n30843, n17490, n6_adj_3925, n28723, n30814, n27790, n30887, 
        n27774, n28784, n28654, n30987, n30742, n1835, n31096, 
        n30, n34, n30823, n30905, n32, n30737, n28648, n33, 
        n30783, n28656, n31, n4_c, n16895, n16963, n27, n16246, 
        n17356, n5_c, n10_c, n17481, n25, n6_adj_3926, n28791, 
        n32882, n30649, n6_adj_3927, n30799, n14900, n6_adj_3928, 
        n27848, n16263, n16736, n6_adj_3929, n17600, n30499, n30884, 
        n17046, n30837, n28736, n28725, n28685, n30505, n12, n31004, 
        n31049, n17053, n14, n30834, n15_c, n16279, n32935, n4_adj_3930, 
        n30635, n1180, n30515, n30489, n10_adj_3931, n27801, n16660, 
        n28707, n31_adj_3932, n31040, n31114, n16891, n16631, n30632, 
        n28310, n31111, n35, n30899, n30623, n34_adj_3933;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n14151, n4752, n30890, n33_adj_3934, n30508, n22, n37, 
        n29, n1241, n39, n17057, n27850, n30749;
    wire [7:0]n8825;
    
    wire n17751;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n17965, n30662;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n33103, n12_adj_3935, n13, n30929, n30598, n10_adj_3936, 
        n18117;
    wire [7:0]\data_out_frame[5]_c ;   // verilog/coms.v(97[12:26])
    
    wire n30689, n10_adj_3937, n30711, n30879, n18116, n30626, n4_adj_3938, 
        n17040, n30553, n30550, n22967, n22634, n13_adj_3939, n6_adj_3940, 
        n32017, n48, n46, n30717, n47, n45, n44, n43, n54, 
        n49, n11, n22829, n17773, n30546, n6_adj_3941, n30846, 
        n6_adj_3942, n16697, n12_adj_3943, n13_adj_3944, n12_adj_3945, 
        n16888, n7_adj_3946, n9, n30473, n6_adj_3947, n28748, n28637, 
        n30521;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n31073, n32357, n30361, n31340, n17807;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(96[12:25])
    
    wire n38, n25_adj_3948, n16797, n33151, n33153, n39_adj_3949, 
        n43_adj_3950, n33159;
    wire [31:0]\FRAME_MATCHER.state_31__N_2515 ;
    
    wire n4_adj_3951, n14112, n7_adj_3952, n16608, n29945, n9_adj_3953, 
        n29837, n6_adj_3954, n29839, n30019, n29841, n13865, n2_adj_3955, 
        n22624, n16429, n30017, n29843, n30015, n30013, n30011, 
        n30009, n30007, n30005, n16619, n29931, n16583, n31439, 
        n5_adj_3956, n6_adj_3957, n30394, n30003, n30001, n29999, 
        n29997, n29995, n18115, n29993, n29991, n29989, n63_c, 
        n63_adj_3958, n29987, n29985, n29983, n29981, n29979, n29977, 
        n29975, n29973, n4753, n29935;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n4776, n4775, n4774, n4773, n18114, n4772, n4771, n29971, 
        n29969, n4770, n4769, n4768, n16607, n6_adj_3962, n4767, 
        n22650, n4766, n4765, n4764, n4763, n4762, n4761, n8_adj_3963, 
        n16594, n4760, n18113, n18112, n22775, n5_adj_3964, tx_transmit_N_3304, 
        n18111, n4759, n4758, n4757, n5_adj_3965, n32365, n32475, 
        n32363, n4756, n14_adj_3966, n4755, n20_adj_3967, n32221, 
        n18, n22_adj_3968, n16441, n14_adj_3969, n16597, n15_adj_3970, 
        n16459, n16_adj_3971, n17, n16541, n10_adj_3972, n10_adj_3973, 
        n14_adj_3974, n16538, n18_adj_3975, n20_adj_3976, n15_adj_3977, 
        n16_adj_3978, n17_adj_3979, n20_adj_3980, n19_c, n33155, n8_adj_3981, 
        n18175, n32881, n13914, n21822, n16611, n11_adj_3982, n29967, 
        n18_adj_3983, n18176, n18177, n2026;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n30946, n16242, n13_adj_3984, n11_adj_3985, n16686, n28787, 
        Kp_23__N_1591, n31075, n30709;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n10_adj_3986, n30809, n28603, n30972, n30695, n31087, n31776, 
        n31081, n31123, n10_adj_3987, n31064, n31043, n27714, n18_adj_3988, 
        n31013, n16714, n16_adj_3989, n30614, n20_adj_3990, n31117, 
        n31058, n30658, n7_adj_3991, n31126, n30955, n16_adj_3992, 
        n27739, n30938, Kp_23__N_1092, n22_adj_3993;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n30620, n20_adj_3994, n31070, n24_adj_3995, n17378, n16978, 
        n30732, n10_adj_3996, n30638, n14_adj_3997, n30671, n28732, 
        n12_adj_3998, n16323, n31836, n32679, n31129, n18092, n8_adj_3999, 
        Kp_23__N_652, n60, Kp_23__N_1293, n31099, n31007, n58, n18093, 
        n4754, n30793, n30752, n59, n18178, n30761, n57, n31132, 
        n31019, n56, n55, n63_adj_4000, n31028, n30960, n62, n68, 
        n30995, n17656, n16657, n61, n69, n32512, n30700, n28_adj_4001, 
        n28650, n30684, n26_adj_4002, n31120, n27_adj_4003, n30866, 
        n28673, n25_adj_4004, n32292, n30611, n30592, n27501, n12_adj_4005, 
        n16927, n30935, n32560, n27776, n30896, n27688, n28614, 
        n12_adj_4006, n30720, n30978, n28756, n32366, n17312, n17529, 
        Kp_23__N_1097, n31_adj_4007;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(130[14:26])
    
    wire n18094, n16785, n30533, n13_adj_4008, n11_adj_4009, n18179, 
        n14_adj_4010, n30787, n15_adj_4011, n17252, n18110;
    wire [0:0]n3276;
    wire [2:0]r_SM_Main_2__N_3407;
    
    wire n31148, n30849, n30902, n15030, n17297, n14_adj_4012, n10_adj_4013, 
        n30764, Kp_23__N_1076, n12_adj_4014, n31010, n31815, n31472, 
        n4854, n31272, n30767, Kp_23__N_1082, n8_adj_4015, n30857, 
        n30796, n30559, n17114, n30963, Kp_23__N_986, n16937, \FRAME_MATCHER.rx_data_ready_prev , 
        n30769, n15_adj_4016, n14_adj_4017, n17642, n24_adj_4018, 
        n22_adj_4019, n26_adj_4020, n30958, n16882, n8_adj_4021, n15023, 
        n14_adj_4022, n10_adj_4023, n30666, n25555, n25556, n30655, 
        n17636, n12_adj_4024, n30745, n28620, n17342, n10_adj_4025, 
        n10_adj_4026, n30629, n32203, n36139, n8_adj_4027, n32739, 
        n32209, n27881, n32713, n7_adj_4028, n10_adj_4029, n32875, 
        n6_adj_4030, n32519, n33080, n22_adj_4031, n33082, n21, 
        n18180, n33084, n30595, n19_adj_4032, n30_adj_4033, n32133, 
        n25_adj_4034, n18181, n18182, n10_adj_4035, n30451, n18167, 
        n18168, n18169, n18170, n18109, n18108, n18171, n18107, 
        n18172, n18173, n18174, n17391, n2_adj_4036, n25584, n25613;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n30920, n30790, n30569, n30923, n30537, n30496, n10_adj_4037, 
        n16_adj_4038, n17_adj_4039, n34084, n34083, n16_adj_4040, 
        n17_adj_4041, n34081, n34080, n16_adj_4042, n6_adj_4043, n5_adj_4044, 
        n17_adj_4045, n33932, n7_adj_4046, n34078, n35618, n35606, 
        n14_adj_4047, n34077, n35690, n34085, n16_adj_4048, n17_adj_4049, 
        n34075, n34074, n16_adj_4050, n2_adj_4051, n25554, n2_adj_4052, 
        n25583, n17_adj_4053, n34072, n34071, n17134, n30755, n10_adj_4054, 
        n17452, n33191, n33192, n16_adj_4055, n17_adj_4056, n30952, 
        n6_adj_4057, n34069, n33183, n33182, n34068, n16910, n10_adj_4058, 
        n17265, n6_adj_4059, n2_adj_4060, n25582, n34376, n5_adj_4061, 
        n16_adj_4062, n17315, n17_adj_4063, n7_adj_4064, n16840, n6_adj_4065, 
        n35576, n35570, n14_adj_4066, n35642, n34063, n34370, n5_adj_4067, 
        n8_adj_4068, n18151, n7_adj_4069, n35552, n35624, n14_adj_4070, 
        n18152, n35648, n34066, n2_adj_4071, n25581, n25612, n25611, 
        n16863, n6_adj_4072, n34364, n5_adj_4073, n7_adj_4074, n34065, 
        n2_adj_4075, n25580, n34064, n35612, n35546, n14_adj_4076, 
        n35660, n34070, n10_adj_4077, n6_adj_4078, n30652, n17277, 
        n14_adj_4079, n16_adj_4080, n5_adj_4081, n7_adj_4082, n17290, 
        n18153, n17_adj_4083, n30981, n34087, n34086, Kp_23__N_855, 
        n35516, n35504, n14_adj_4084, n35666, n34073, n30587, Kp_23__N_779, 
        n17135, n10_adj_4085, n6_adj_4086, n30840, n2_adj_4087, n25579, 
        n27737, Kp_23__N_784, n6_adj_4088, Kp_23__N_884, n30566, n25610, 
        n18154, n30831, n30604, n18155, n16730, n30512, n6_adj_4089, 
        n16832, n30572, n5_adj_4090, n7_adj_4091, n29939, n30584, 
        n25609, n29927, n29923, n29919, n29915, n29911, n29907, 
        n29903, n21837, n30725, n29899, n29895, n29891, n29887, 
        n29883, n35510, n35654, n14_adj_4092, n29879, n29875, n29871, 
        n29867, n29863, n29859, n29855, n29851, n29847, n15796, 
        n29835, n35672, n34076, n31067, n6_adj_4093, n2_adj_4094, 
        n25578, n31055, n5_adj_4095, n7_adj_4096, n25608, n30932, 
        n28_adj_4097, n18156, n14_adj_4098, n2_adj_4099, n25577, n30926, 
        n15_adj_4100, n32550, n32_adj_4101, n35678, n34079, n30601, 
        n30_adj_4102, n18157, n31_adj_4103, Kp_23__N_811, n29_adj_4104, 
        n34344, n18158, n5_adj_4105, n32090;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n7_adj_4106, n25607, n21993, n18143, n16999, n35564, n35558, 
        n14_adj_4107, n12_adj_4108, n35684, n34082, n18_adj_4109, 
        n18144, n2_adj_4110, n25576, n18145, n18146, n18147, n32617, 
        n18148, n31607, n30542, n32125, n31666, n30861, n32161, 
        n31697;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n32219, n32412, n31422, n31772, n32037, n31747, n32377, 
        n3_adj_4111, n18149, n18150, n10_adj_4112, n30455, n18135, 
        n18136, n3_adj_4113, n3_adj_4114, n3_adj_4115, n3_adj_4116, 
        n3_adj_4117, n3_adj_4118, n3_adj_4119, n3_adj_4120, n2_adj_4121, 
        n3_adj_4122, n2_adj_4123, n3_adj_4124, n25575, n2_adj_4125, 
        n3_adj_4126, n2_adj_4127, n3_adj_4128, n2_adj_4129, n3_adj_4130, 
        n2_adj_4131, n3_adj_4132, n2_adj_4133, n3_adj_4134, n2_adj_4135, 
        n3_adj_4136, n2_adj_4137, n3_adj_4138, n2_adj_4139, n3_adj_4140, 
        n2_adj_4141, n3_adj_4142, n2_adj_4143, n3_adj_4144, n2_adj_4145, 
        n3_adj_4146, n2_adj_4147, n3_adj_4148, n2_adj_4149, n3_adj_4150, 
        n2_adj_4151, n3_adj_4152, n2_adj_4153, n3_adj_4154, n2_adj_4155, 
        n3_adj_4156, n2_adj_4157, n3_adj_4158, n2_adj_4159, n3_adj_4160, 
        n2_adj_4161, n3_adj_4162, n25574, n3_adj_4163, n25573, n18137, 
        n25572, n18138, n25571, n18139, n18140, n18141, n25570, 
        n161, n25569, n18142, n30447, n18127, n18106, n18128, 
        n18129, n18130, n18131, n18132, n18133, n18105, n18104, 
        n18103, n25568, n18134, n10_adj_4164, n14_adj_4165, n25567, 
        n25566, n21985, n21830, n32888, n25565, n10_adj_4166, n21709, 
        n21710, n28_adj_4168, n26_adj_4171, n25564, n25563, n27_adj_4172, 
        n25_adj_4173, n35456, n35729;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n35462, n35723, n35630, n35468, n35717, n25562, n35474, 
        n35711, n35480, n35705, n35486, n35699, n35492, n35693, 
        n35687, n35681, n35675, n35669, n35663, n35657, n35651, 
        n35645, n25561, n35639, n35627, n35621, n35615, n35609, 
        n35603, n35498, n35579, n35573, n35567, n35561, n35555, 
        n35549, n35543, n25560, n35513, n30562, n9_adj_4174, n14898, 
        n30802, n25559, n27823, n31016, n6_adj_4175, n2483, n6_adj_4176, 
        n25558, n17262, n14_adj_4177, n10_adj_4178, n31034, n21861, 
        n10_adj_4179, n30463, n31025, n30739, n10_adj_4180, n30486, 
        n31052, n25557, n30770, n16671, n28699, n4_adj_4181, n28702, 
        n16822, n30828, n30860, n30575, n31061, n6_adj_4182, n28622, 
        n30969, n32847, n28667, n2196, n10_adj_4183, n17937, n28697, 
        n6_adj_4184, n16604, n28610, n32564, n31084, n30643, n8_adj_4185, 
        n31102, n27760, n35507, n18449, n18448, n18054, n18263, 
        n18264, n18265, n18266, n18267, n18268, n30874, n18269, 
        n18053, n35501, n30459, n18121, n18122, n18123, n18124, 
        n18262, n18261, n18260, n18259, n18258, n18257, n18256, 
        n18255, n18254, n18253, n18252, n18251, n18250, n18249, 
        n18248, n18247, n18246, n18245, n18244, n18243, n18242, 
        n18241, n18240, n18239, n18238, n18237, n18236, n18235, 
        n18234, n18233, n18232, n18231, n18222, n18221, n18125, 
        n18220, n18219, n18218, n18217, n18216, n18215, n18214, 
        n18213, n18212, n18211, n18210, n18209, n18208, n18207, 
        n18126, n18206, n18205, n18204, n18203, n18202, n18201, 
        n18200, n18199, n18198, n18197, n18196, n18195, n18194, 
        n18193, n18192, n18191, n18190, n18189, n18188, n18187, 
        n18186, n18185, n18184, n18183, n30863, n35495, n35489, 
        n35483, n30870, n18_adj_4187, n31078, n20_adj_4188, n28404, 
        n15_adj_4189, n31901, n28379, n30778, n14_adj_4190, n31022, 
        n30806, n17226, n31108, n35477, n31712, n10_adj_4191, n30966, 
        n1, n30_adj_4192, n34_adj_4193, n32_adj_4194, n30729, n33_adj_4195, 
        n35471, n17457, n31_adj_4196, n17440, n28631, n27784, n30541, 
        n30998, n31001, n30992, n15_adj_4197, n10_adj_4198, n30758, 
        n30820, n2066, n12_adj_4199, n28730, n12_adj_4200, n14_adj_4201, 
        n32095, n30527, n35465, n35459, n35453, n33129, n13703;
    
    SB_LUT4 i10_4_lut (.I0(n30913), .I1(n20), .I2(n16), .I3(n30556), 
            .O(n31662));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18120));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_3_lut (.I0(n30852), .I1(n24), .I2(n28088), .I3(GND_net), 
            .O(n28));
    defparam i12_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i10_4_lut_adj_841 (.I0(n28125), .I1(n8), .I2(n16954), .I3(n17350), 
            .O(n26));
    defparam i10_4_lut_adj_841.LUT_INIT = 16'hffef;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18119));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[14] [1]), .I1(n16878), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n30502));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut (.I0(\data_out_frame[12] [0]), .I1(n30502), .I2(n17336), 
            .I3(GND_net), .O(n16702));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30524));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(n30524), .I2(n32089), .I3(n2112), 
            .O(n30949));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_842 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n30703));
    defparam i2_3_lut_adj_842.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[19] [1]), .I1(n30703), .I2(n30493), 
            .I3(\data_out_frame[19] [6]), .O(n2112));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_843 (.I0(\data_out_frame[13] [4]), .I1(n16666), 
            .I2(n30714), .I3(GND_net), .O(n31093));
    defparam i1_3_lut_adj_843.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_844 (.I0(\data_out_frame[15] [2]), .I1(n28782), 
            .I2(n28681), .I3(n6), .O(n28740));
    defparam i4_4_lut_adj_844.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18118));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[15] [5]), .I1(n30714), .I2(n30817), 
            .I3(n27756), .O(n28767));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_845 (.I0(n28767), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30773));
    defparam i1_2_lut_adj_845.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n30468), .I3(\FRAME_MATCHER.i [0]), .O(n30471));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n31090));
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_847 (.I0(n30617), .I1(n30843), .I2(GND_net), 
            .I3(GND_net), .O(n17490));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_848 (.I0(n16666), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3925));
    defparam i1_2_lut_adj_848.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_849 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[13] [2]), 
            .I2(n28681), .I3(n6_adj_3925), .O(n28723));
    defparam i4_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_850 (.I0(\data_out_frame[15] [3]), .I1(n30814), 
            .I2(n17490), .I3(n27756), .O(n27790));
    defparam i3_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_851 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30887));
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_852 (.I0(n27790), .I1(\data_out_frame[17] [5]), 
            .I2(n28723), .I3(GND_net), .O(n27774));
    defparam i2_3_lut_adj_852.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_853 (.I0(n28784), .I1(n28654), .I2(GND_net), 
            .I3(GND_net), .O(n30987));
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_854 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30742));
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(71[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut (.I0(n31096), .I1(n1835), .I2(n30742), .I3(n30987), 
            .O(n30));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n27774), .I1(n30), .I2(\data_out_frame[16] [0]), 
            .I3(n30887), .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n31090), .I1(n30823), .I2(n30905), .I3(n30773), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(n30737), .I1(n16878), .I2(n28740), .I3(n28648), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(n30783), .I1(n28656), .I2(n32089), .I3(\data_out_frame[17] [7]), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_855 (.I0(n4_c), .I1(n31662), .I2(n16895), .I3(n16963), 
            .O(n27));
    defparam i11_4_lut_adj_855.LUT_INIT = 16'hfeff;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n16246));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17356), .I1(n5_c), .I2(n10_c), .I3(n17481), 
            .O(n25));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_856 (.I0(\data_in_frame[19] [6]), .I1(n6_adj_3926), 
            .I2(n28791), .I3(\data_in_frame[19] [5]), .O(n32882));
    defparam i3_4_lut_adj_856.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_857 (.I0(\data_out_frame[19] [0]), .I1(n30649), 
            .I2(n2112), .I3(n6_adj_3927), .O(n30799));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_858 (.I0(n14900), .I1(n30799), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3928));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_859 (.I0(\data_out_frame[18] [6]), .I1(n27848), 
            .I2(\data_out_frame[18] [4]), .I3(n6_adj_3928), .O(n16263));
    defparam i4_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_860 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[11] [6]), 
            .I2(n16736), .I3(n6_adj_3929), .O(n17600));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_860.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_861 (.I0(n30499), .I1(n30884), .I2(\data_out_frame[5] [5]), 
            .I3(GND_net), .O(n17046));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_861.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_862 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[13] [0]), 
            .I2(n30837), .I3(n28736), .O(n28725));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_863 (.I0(\data_out_frame[17] [2]), .I1(n28648), 
            .I2(n28725), .I3(GND_net), .O(n28784));
    defparam i1_3_lut_adj_863.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut (.I0(n28685), .I1(n31096), .I2(n17046), .I3(n30505), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[12] [2]), .I1(n12), .I2(\data_out_frame[17] [0]), 
            .I3(n31004), .O(n30823));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30493));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_865 (.I0(\data_out_frame[12] [0]), .I1(n30905), 
            .I2(GND_net), .I3(GND_net), .O(n31049));
    defparam i1_2_lut_adj_865.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut (.I0(n17053), .I1(\data_out_frame[19] [0]), .I2(n30823), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_866 (.I0(n31049), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[14] [2]), .I3(n30834), .O(n15_c));
    defparam i6_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_c), .I1(n17600), .I2(n14), .I3(\data_out_frame[16] [4]), 
            .O(n16279));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_867 (.I0(\data_out_frame[14] [3]), .I1(n32935), 
            .I2(GND_net), .I3(GND_net), .O(n30505));
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_868 (.I0(\data_out_frame[7] [5]), .I1(n4_adj_3930), 
            .I2(n30635), .I3(n1180), .O(n16878));
    defparam i3_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_869 (.I0(n30515), .I1(\data_out_frame[16] [5]), 
            .I2(n17053), .I3(GND_net), .O(n27848));
    defparam i2_3_lut_adj_869.LUT_INIT = 16'h9696;
    SB_LUT4 i392_2_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1180));   // verilog/coms.v(74[16:27])
    defparam i392_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_870 (.I0(\data_out_frame[14] [4]), .I1(n30884), 
            .I2(n30489), .I3(\data_out_frame[12] [2]), .O(n10_adj_3931));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_871 (.I0(\data_out_frame[14] [5]), .I1(n32935), 
            .I2(n27801), .I3(n16660), .O(n28707));
    defparam i3_4_lut_adj_871.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_872 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n31_adj_3932));
    defparam i15_4_lut_adj_872.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_873 (.I0(n31040), .I1(n31114), .I2(n16891), .I3(GND_net), 
            .O(n30489));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_873.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_874 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16631));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_874.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_875 (.I0(\data_out_frame[6] [3]), .I1(n30632), 
            .I2(\data_out_frame[10] [5]), .I3(n16631), .O(n30843));
    defparam i3_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_876 (.I0(n28310), .I1(n30843), .I2(\data_out_frame[14] [7]), 
            .I3(GND_net), .O(n28736));
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_877 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n31114));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_877.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_878 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3930));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_878.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_879 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[8] [6]), .I3(n31111), .O(n35));
    defparam i14_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_880 (.I0(n30899), .I1(n30499), .I2(n30623), 
            .I3(\data_out_frame[6] [2]), .O(n34_adj_3933));
    defparam i13_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_881 (.I0(n31_adj_3932), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n14151), .I3(GND_net), .O(n4752));
    defparam i2_3_lut_adj_881.LUT_INIT = 16'h0404;
    SB_LUT4 i12_4_lut_adj_882 (.I0(n31114), .I1(\data_out_frame[6] [0]), 
            .I2(n30890), .I3(\data_out_frame[10] [1]), .O(n33_adj_3934));
    defparam i12_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n16891), .I1(n30508), .I2(\data_out_frame[6] [4]), 
            .I3(n22), .O(n37));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_883 (.I0(n35), .I1(n29), .I2(\data_out_frame[5] [4]), 
            .I3(n1241), .O(n39));
    defparam i18_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n39), .I1(n37), .I2(n33_adj_3934), .I3(n34_adj_3933), 
            .O(n32935));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_884 (.I0(\data_out_frame[13] [5]), .I1(n17057), 
            .I2(n30714), .I3(GND_net), .O(n27850));
    defparam i1_3_lut_adj_884.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30749));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n17751), .D(n8825[7]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_886 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30662));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_886.LUT_INIT = 16'h6666;
    SB_LUT4 i26934_2_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33103));
    defparam i26934_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_887 (.I0(\data_out_frame[9] [0]), .I1(n30662), 
            .I2(\data_out_frame[11] [1]), .I3(\data_out_frame[6] [3]), .O(n12_adj_3935));   // verilog/coms.v(85[17:63])
    defparam i5_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_888 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [6]), .O(n13));
    defparam i5_4_lut_adj_888.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(n33103), .I2(\data_in_frame[0] [1]), 
            .I3(\data_in_frame[0] [5]), .O(n14151));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_889 (.I0(\data_out_frame[6] [6]), .I1(n12_adj_3935), 
            .I2(n30749), .I3(\data_out_frame[10] [7]), .O(n27756));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_890 (.I0(n30929), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[11] [0]), .I3(n30598), .O(n28681));
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n17751), .D(n8825[6]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16660));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_892 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[11] [2]), .I3(n30623), .O(n10_adj_3936));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18117));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[5]_c [1]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30508));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30689));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_out_frame[5][7] ), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n31040));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n17751), .D(n8825[5]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_896 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[11] [5]), .I3(n30890), .O(n10_adj_3937));
    defparam i4_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_897 (.I0(\data_out_frame[5]_c [0]), .I1(n10_adj_3937), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n17336));
    defparam i5_3_lut_adj_897.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_898 (.I0(\data_out_frame[5]_c [1]), .I1(\data_out_frame[5]_c [0]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n16736));
    defparam i2_3_lut_adj_898.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_899 (.I0(\data_out_frame[11] [4]), .I1(n30711), 
            .I2(n16736), .I3(\data_out_frame[9] [2]), .O(n17057));
    defparam i3_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30879));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n17751), .D(n8825[4]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n17751), .D(n8825[3]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18116));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_901 (.I0(\data_out_frame[5]_c [1]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[11] [7]), .O(n30635));
    defparam i3_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(n30626), .I1(\data_out_frame[11] [3]), .I2(\data_out_frame[6] [5]), 
            .I3(n4_adj_3938), .O(n30714));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_902 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17040));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_903 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[9] [2]), .O(n30626));
    defparam i3_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30553));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_905 (.I0(n30929), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[6] [4]), .O(n30617));   // verilog/coms.v(76[16:43])
    defparam i2_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30550));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_907 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30817));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n28310), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28782));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_909 (.I0(n27801), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n30837));
    defparam i2_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_910 (.I0(\FRAME_MATCHER.state[0] ), .I1(n14151), 
            .I2(n22967), .I3(n22634), .O(n13_adj_3939));
    defparam i5_4_lut_adj_910.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_911 (.I0(n28782), .I1(\data_out_frame[13] [5]), 
            .I2(n30817), .I3(n6_adj_3940), .O(n32017));
    defparam i4_4_lut_adj_911.LUT_INIT = 16'h9669;
    SB_LUT4 i20_4_lut_adj_912 (.I0(n30550), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[10] [5]), .I3(\data_out_frame[9] [0]), .O(n48));
    defparam i20_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_913 (.I0(n30553), .I1(n17057), .I2(\data_out_frame[7] [4]), 
            .I3(\data_out_frame[12] [0]), .O(n46));
    defparam i18_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n31111), .I1(n30635), .I2(n30717), .I3(n30598), 
            .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n30626), .I1(n17040), .I2(n30714), .I3(n30711), 
            .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_914 (.I0(n17336), .I1(n31040), .I2(n30689), 
            .I3(\data_out_frame[11] [6]), .O(n44));
    defparam i16_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_915 (.I0(n27850), .I1(n32017), .I2(n32935), 
            .I3(n30617), .O(n43));
    defparam i15_4_lut_adj_915.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n16666), .I1(n16660), .I2(n28681), .I3(n27756), 
            .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i28778_4_lut (.I0(n13_adj_3939), .I1(n11), .I2(n22829), .I3(\FRAME_MATCHER.state [2]), 
            .O(n17773));
    defparam i28778_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(n28656));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_916 (.I0(\data_out_frame[5][7] ), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30632));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_916.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_917 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30546));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[5][6] ), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16891));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_919 (.I0(n1241), .I1(n30546), .I2(\data_out_frame[10] [4]), 
            .I3(n6_adj_3941), .O(n30846));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[5][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3942));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_921 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(n30899), .I3(n6_adj_3942), .O(n27801));
    defparam i4_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_922 (.I0(\data_out_frame[12] [5]), .I1(n27801), 
            .I2(n30846), .I3(GND_net), .O(n30717));
    defparam i1_3_lut_adj_922.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16697));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_924 (.I0(\data_out_frame[14] [5]), .I1(n12_adj_3943), 
            .I2(n28656), .I3(\data_out_frame[14] [6]), .O(n28685));
    defparam i6_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_925 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [4]), .I3(\data_out_frame[15] [0]), 
            .O(n13_adj_3944));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_926 (.I0(n13_adj_3944), .I1(n27801), .I2(n12_adj_3945), 
            .I3(n30617), .O(n28648));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_926.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_927 (.I0(n16888), .I1(n28648), .I2(\data_out_frame[17] [1]), 
            .I3(n28685), .O(n7_adj_3946));
    defparam i1_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_928 (.I0(n9), .I1(n7_adj_3946), .I2(\data_out_frame[12] [3]), 
            .I3(n32935), .O(n28654));
    defparam i5_4_lut_adj_928.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_929 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n30473), .I3(\FRAME_MATCHER.i [0]), .O(n30475));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_929.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_adj_930 (.I0(n28707), .I1(n30515), .I2(\data_out_frame[16] [6]), 
            .I3(GND_net), .O(n32089));
    defparam i2_3_lut_adj_930.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_931 (.I0(\data_out_frame[18] [7]), .I1(n30834), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3947));
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_932 (.I0(n32089), .I1(\data_out_frame[19] [2]), 
            .I2(n28654), .I3(n6_adj_3947), .O(n28748));
    defparam i4_4_lut_adj_932.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_933 (.I0(n28748), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28637));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30521));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_935 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [2]), 
            .I2(n31073), .I3(GND_net), .O(n32357));
    defparam i2_3_lut_adj_935.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_936 (.I0(\FRAME_MATCHER.state[3] ), .I1(n22632), 
            .I2(GND_net), .I3(GND_net), .O(n30361));
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_937 (.I0(n22829), .I1(n22967), .I2(n22634), .I3(GND_net), 
            .O(n31340));
    defparam i2_3_lut_adj_937.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_938 (.I0(\FRAME_MATCHER.state [1]), .I1(n31340), 
            .I2(n30361), .I3(GND_net), .O(n17807));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[7] [6]), .O(n30499));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_939 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[1]_c [2]), .O(n38));
    defparam i14_4_lut_adj_939.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[1]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3948));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h8888;
    SB_LUT4 i26979_4_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(n16797), .I3(\data_in_frame[2] [0]), .O(n33151));
    defparam i26979_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26981_4_lut (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[0] [1]), .O(n33153));
    defparam i26981_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_941 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1]_c [1]), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[2] [5]), .O(n39_adj_3949));
    defparam i15_4_lut_adj_941.LUT_INIT = 16'h0002;
    SB_LUT4 i19_4_lut_adj_942 (.I0(n25_adj_3948), .I1(n38), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[1][7] ), .O(n43_adj_3950));
    defparam i19_4_lut_adj_942.LUT_INIT = 16'h0800;
    SB_LUT4 i26987_4_lut (.I0(n33151), .I1(\data_in_frame[2] [6]), .I2(n33103), 
            .I3(\data_in_frame[0] [0]), .O(n33159));
    defparam i26987_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n33159), .I1(n43_adj_3950), .I2(n39_adj_3949), 
            .I3(n33153), .O(\FRAME_MATCHER.state_31__N_2515 [3]));
    defparam i23_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i1_4_lut_adj_943 (.I0(\FRAME_MATCHER.state[3] ), .I1(n16613), 
            .I2(n4_adj_3951), .I3(n14112), .O(n7_adj_3952));
    defparam i1_4_lut_adj_943.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_944 (.I0(\FRAME_MATCHER.state [2]), .I1(n7_adj_3952), 
            .I2(n16608), .I3(\FRAME_MATCHER.state_31__N_2515 [3]), .O(n29945));
    defparam i1_4_lut_adj_944.LUT_INIT = 16'hcdcc;
    SB_LUT4 i1_2_lut_adj_945 (.I0(\FRAME_MATCHER.state [4]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29837));
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_946 (.I0(\FRAME_MATCHER.state [4]), .I1(n6_adj_3954), 
            .I2(GND_net), .I3(GND_net), .O(n29839));
    defparam i1_2_lut_adj_946.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\FRAME_MATCHER.state [5]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30019));
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\FRAME_MATCHER.state [5]), .I1(n6_adj_3954), 
            .I2(GND_net), .I3(GND_net), .O(n29841));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n13865), .I1(n2_adj_3955), .I2(n22624), 
            .I3(n16429), .O(n6_adj_3954));
    defparam i1_4_lut_adj_949.LUT_INIT = 16'hccec;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\FRAME_MATCHER.state [6]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30017));
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\FRAME_MATCHER.state [6]), .I1(n6_adj_3954), 
            .I2(GND_net), .I3(GND_net), .O(n29843));
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_952 (.I0(\FRAME_MATCHER.state [7]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30015));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\FRAME_MATCHER.state [8]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30013));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\FRAME_MATCHER.state [9]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30011));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\FRAME_MATCHER.state [10]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30009));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\FRAME_MATCHER.state [11]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30007));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\FRAME_MATCHER.state [12]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30005));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [29]), .O(n29931));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hf400;
    SB_LUT4 i28920_3_lut (.I0(n22632), .I1(n31340), .I2(n16583), .I3(GND_net), 
            .O(n31439));
    defparam i28920_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i28986_4_lut (.I0(n16583), .I1(n4922), .I2(n5_adj_3956), .I3(n6_adj_3957), 
            .O(n30394));
    defparam i28986_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\FRAME_MATCHER.state [13]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30003));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_959 (.I0(\FRAME_MATCHER.state [14]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n30001));
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\FRAME_MATCHER.state [15]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29999));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_961 (.I0(\FRAME_MATCHER.state [16]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29997));
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_962 (.I0(\FRAME_MATCHER.state [17]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29995));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18115));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_963 (.I0(\FRAME_MATCHER.state [18]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29993));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\FRAME_MATCHER.state [19]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29991));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_965 (.I0(\FRAME_MATCHER.state [20]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29989));
    defparam i1_2_lut_adj_965.LUT_INIT = 16'h8888;
    SB_LUT4 i17502_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), .I2(n63_adj_3958), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i17502_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_404_Select_2_i5_4_lut (.I0(n122), .I1(n16606), .I2(n3303), 
            .I3(n63), .O(n5));
    defparam select_404_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_966 (.I0(\FRAME_MATCHER.state [21]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29987));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_967 (.I0(\FRAME_MATCHER.state [22]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29985));
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\FRAME_MATCHER.state [23]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29983));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\FRAME_MATCHER.state [24]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29981));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\FRAME_MATCHER.state [25]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29979));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_971 (.I0(\FRAME_MATCHER.state [26]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29977));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h8888;
    SB_LUT4 i17496_rep_267_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n36350));   // verilog/coms.v(142[4] 144[7])
    defparam i17496_rep_267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\FRAME_MATCHER.state [27]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29975));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\FRAME_MATCHER.state [28]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29973));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1266_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4752), .I3(GND_net), .O(n4753));
    defparam mux_1266_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_974 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [30]), .O(n29935));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_974.LUT_INIT = 16'hf400;
    SB_LUT4 mux_1266_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1][7] ), 
            .I2(n4752), .I3(GND_net), .O(n4776));
    defparam mux_1266_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[13] [2]), .I3(GND_net), .O(n30814));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_975 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[18] [3]), .I3(GND_net), .O(n30649));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_975.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1266_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1][6] ), 
            .I2(n4752), .I3(GND_net), .O(n4775));
    defparam mux_1266_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4752), .I3(GND_net), .O(n4774));
    defparam mux_1266_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4752), .I3(GND_net), .O(n4773));
    defparam mux_1266_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18114));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1266_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n4752), .I3(GND_net), .O(n4772));
    defparam mux_1266_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1]_c [2]), 
            .I2(n4752), .I3(GND_net), .O(n4771));
    defparam mux_1266_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_976 (.I0(\FRAME_MATCHER.state [29]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29971));
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_977 (.I0(\FRAME_MATCHER.state [30]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29969));
    defparam i1_2_lut_adj_977.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1266_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n4752), .I3(GND_net), .O(n4770));
    defparam mux_1266_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1]_c [0]), 
            .I2(n4752), .I3(GND_net), .O(n4769));
    defparam mux_1266_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4752), .I3(GND_net), .O(n4768));
    defparam mux_1266_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_978 (.I0(n16607), .I1(n63_adj_3), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3962));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h8888;
    SB_LUT4 mux_1266_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4752), .I3(GND_net), .O(n4767));
    defparam mux_1266_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_979 (.I0(n16608), .I1(n22650), .I2(n16619), .I3(n6_adj_3962), 
            .O(n2696));
    defparam i4_4_lut_adj_979.LUT_INIT = 16'h8000;
    SB_LUT4 mux_1266_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4752), .I3(GND_net), .O(n4766));
    defparam mux_1266_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4752), .I3(GND_net), .O(n4765));
    defparam mux_1266_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4752), .I3(GND_net), .O(n4764));
    defparam mux_1266_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4752), .I3(GND_net), .O(n4763));
    defparam mux_1266_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4752), .I3(GND_net), .O(n4762));
    defparam mux_1266_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4752), .I3(GND_net), .O(n4761));
    defparam mux_1266_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17473_4_lut (.I0(n8_adj_3963), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n16594), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i17473_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 mux_1266_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4752), .I3(GND_net), .O(n4760));
    defparam mux_1266_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18112));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28757_2_lut (.I0(n22775), .I1(n5_adj_3964), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3304));
    defparam i28757_2_lut.LUT_INIT = 16'h1111;
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18111));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_980 (.I0(n16621), .I1(n4452), .I2(n13810), .I3(GND_net), 
            .O(n2_adj_3955));
    defparam i1_3_lut_adj_980.LUT_INIT = 16'h1010;
    SB_LUT4 mux_1266_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4752), .I3(GND_net), .O(n4759));
    defparam mux_1266_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4752), .I3(GND_net), .O(n4758));
    defparam mux_1266_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1266_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4752), .I3(GND_net), .O(n4757));
    defparam mux_1266_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17471_4_lut (.I0(n5_adj_3965), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i17471_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i3_4_lut_adj_981 (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(\FRAME_MATCHER.i [7]), .I3(\FRAME_MATCHER.i [9]), .O(n32365));
    defparam i3_4_lut_adj_981.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_982 (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [6]), .I3(\FRAME_MATCHER.i [8]), .O(n32475));
    defparam i3_4_lut_adj_982.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_983 (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [23]), .I3(\FRAME_MATCHER.i [19]), .O(n32363));
    defparam i3_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1266_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4752), .I3(GND_net), .O(n4756));
    defparam mux_1266_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_984 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n32365), .O(n14_adj_3966));
    defparam i2_4_lut_adj_984.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1266_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4752), .I3(GND_net), .O(n4755));
    defparam mux_1266_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_985 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [29]), 
            .I2(n32475), .I3(\FRAME_MATCHER.i [24]), .O(n20_adj_3967));
    defparam i8_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_986 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [16]), .I3(\FRAME_MATCHER.i [14]), .O(n32221));
    defparam i3_4_lut_adj_986.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(GND_net), .I3(GND_net), .O(n18));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_987 (.I0(n32221), .I1(n20_adj_3967), .I2(n14_adj_3966), 
            .I3(n32363), .O(n22_adj_3968));
    defparam i10_4_lut_adj_987.LUT_INIT = 16'hfffe;
    SB_LUT4 i5218_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n9711));   // verilog/coms.v(157[6] 159[9])
    defparam i5218_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11_4_lut_adj_988 (.I0(\FRAME_MATCHER.i [30]), .I1(n22_adj_3968), 
            .I2(n18), .I3(\FRAME_MATCHER.i [18]), .O(n16594));
    defparam i11_4_lut_adj_988.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_989 (.I0(\FRAME_MATCHER.i [4]), .I1(n16594), .I2(GND_net), 
            .I3(GND_net), .O(n16441));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_989.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_990 (.I0(n63), .I1(n3303), .I2(n123), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2579[1] ));
    defparam i2_3_lut_adj_990.LUT_INIT = 16'hfdfd;
    SB_LUT4 i5_3_lut_adj_991 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_3969));
    defparam i5_3_lut_adj_991.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_992 (.I0(\data_in[0] [6]), .I1(n16597), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_3970));
    defparam i6_4_lut_adj_992.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_993 (.I0(n15_adj_3970), .I1(\data_in[2] [2]), .I2(n14_adj_3969), 
            .I3(\data_in[3] [0]), .O(n16459));
    defparam i8_4_lut_adj_993.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_994 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3971));
    defparam i6_4_lut_adj_994.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_995 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_995.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_996 (.I0(n17), .I1(\data_in[1] [6]), .I2(n16_adj_3971), 
            .I3(\data_in[3] [7]), .O(n16541));
    defparam i9_4_lut_adj_996.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_997 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3972));
    defparam i4_4_lut_adj_997.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_998 (.I0(\data_in[3] [4]), .I1(n10_adj_3972), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n16597));
    defparam i5_3_lut_adj_998.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3973));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_999 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3974));
    defparam i6_4_lut_adj_999.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1000 (.I0(\data_in[3] [6]), .I1(n14_adj_3974), 
            .I2(n10_adj_3973), .I3(\data_in[2] [1]), .O(n16538));
    defparam i7_4_lut_adj_1000.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1001 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n16538), .I3(\data_in[1] [0]), .O(n18_adj_3975));
    defparam i7_4_lut_adj_1001.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1002 (.I0(\data_in[1] [4]), .I1(n18_adj_3975), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n20_adj_3976));
    defparam i9_4_lut_adj_1002.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_1003 (.I0(n15_adj_3977), .I1(n20_adj_3976), .I2(n16541), 
            .I3(\data_in[0] [6]), .O(n63_c));
    defparam i10_4_lut_adj_1003.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1004 (.I0(\data_in[3] [6]), .I1(n16459), .I2(\data_in[2] [1]), 
            .I3(\data_in[0] [7]), .O(n16_adj_3978));
    defparam i6_4_lut_adj_1004.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1005 (.I0(n16541), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [5]), .O(n17_adj_3979));
    defparam i7_4_lut_adj_1005.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1006 (.I0(n17_adj_3979), .I1(\data_in[3] [3]), 
            .I2(n16_adj_3978), .I3(\data_in[3] [1]), .O(n63_adj_3958));
    defparam i9_4_lut_adj_1006.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_1007 (.I0(n16459), .I1(n16538), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [5]), .O(n20_adj_3980));
    defparam i8_4_lut_adj_1007.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_1008 (.I0(\data_in[2] [5]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[2] [6]), .O(n19_c));
    defparam i7_4_lut_adj_1008.LUT_INIT = 16'hfffd;
    SB_LUT4 i26983_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[0] [1]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n33155));
    defparam i26983_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n33155), .I1(n19_c), .I2(n20_adj_3980), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i13595_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n18175));
    defparam i13595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17472_4_lut (.I0(n32881), .I1(\FRAME_MATCHER.i [31]), .I2(n16441), 
            .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i17472_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(n3303), .I1(n13810), .I2(GND_net), 
            .I3(GND_net), .O(n13914));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(n13810), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n14112));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n21822), .I1(n14112), .I2(n13914), 
            .I3(n16611), .O(n11_adj_3982));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'ha0ec;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\FRAME_MATCHER.state [31]), .I1(n9_adj_3953), 
            .I2(GND_net), .I3(GND_net), .O(n29967));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut_4_lut (.I0(n8), .I1(\data_in_frame[9] [5]), .I2(\data_in_frame[9] [7]), 
            .I3(\data_in_frame[9] [6]), .O(n18_adj_3983));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13596_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n18176));
    defparam i13596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut_4_lut_adj_1013 (.I0(n30489), .I1(n30879), .I2(\data_out_frame[5] [4]), 
            .I3(n28736), .O(n12_adj_3945));   // verilog/coms.v(71[16:27])
    defparam i4_2_lut_4_lut_adj_1013.LUT_INIT = 16'h9669;
    SB_LUT4 i13597_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n18177));
    defparam i13597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18077_1_lut (.I0(n22650), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2026));
    defparam i18077_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut_adj_1014 (.I0(\data_in_frame[14] [1]), .I1(n30946), 
            .I2(n16242), .I3(\data_in_frame[11] [3]), .O(n13_adj_3984));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1015 (.I0(n13_adj_3984), .I1(n11_adj_3985), .I2(n16686), 
            .I3(n28787), .O(Kp_23__N_1591));   // verilog/coms.v(70[16:27])
    defparam i7_4_lut_adj_1015.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1016 (.I0(\data_in_frame[18] [4]), .I1(n31075), 
            .I2(n30709), .I3(\data_in_frame[16] [3]), .O(n10_adj_3986));
    defparam i4_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1017 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[11] [6]), 
            .I2(n30809), .I3(n28603), .O(n30972));
    defparam i3_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1018 (.I0(n30695), .I1(n31087), .I2(n30972), 
            .I3(n30946), .O(n31776));
    defparam i3_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1019 (.I0(n31081), .I1(\data_in_frame[18] [0]), 
            .I2(n10_c), .I3(n31123), .O(n10_adj_3987));
    defparam i4_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1020 (.I0(n31064), .I1(n31043), .I2(n27714), 
            .I3(\data_in_frame[4] [7]), .O(n18_adj_3988));
    defparam i7_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(n31013), .I1(n16714), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_3989));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1021 (.I0(n16686), .I1(n18_adj_3988), .I2(\data_in_frame[14] [2]), 
            .I3(n30614), .O(n20_adj_3990));
    defparam i9_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1022 (.I0(n31117), .I1(n20_adj_3990), .I2(n16_adj_3989), 
            .I3(n31058), .O(n30709));
    defparam i10_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1023 (.I0(\data_in_frame[19] [0]), .I1(n30658), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3991));
    defparam i2_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1024 (.I0(n7_adj_3991), .I1(\data_in_frame[16] [4]), 
            .I2(n30709), .I3(n31126), .O(n30955));
    defparam i4_4_lut_adj_1024.LUT_INIT = 16'h9669;
    SB_LUT4 i3_2_lut (.I0(n16954), .I1(n17481), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_3992));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1025 (.I0(\data_in_frame[17] [4]), .I1(n27739), 
            .I2(n30938), .I3(Kp_23__N_1092), .O(n22_adj_3993));
    defparam i9_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(\data_in_frame[15] [3]), .I1(n30620), .I2(\data_in_frame[15] [2]), 
            .I3(GND_net), .O(n20_adj_3994));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1026 (.I0(\data_in_frame[11] [1]), .I1(n22_adj_3993), 
            .I2(n16_adj_3992), .I3(n31070), .O(n24_adj_3995));
    defparam i11_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1027 (.I0(n17378), .I1(n24_adj_3995), .I2(n20_adj_3994), 
            .I3(\data_in_frame[13] [0]), .O(n16978));
    defparam i12_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30695));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(n8), .I1(\data_in_frame[13] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n30938));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1030 (.I0(n30732), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3996));
    defparam i2_2_lut_adj_1030.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1031 (.I0(n30938), .I1(n30638), .I2(n30695), 
            .I3(\data_in_frame[15] [5]), .O(n14_adj_3997));
    defparam i6_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1032 (.I0(\data_in_frame[9] [1]), .I1(n14_adj_3997), 
            .I2(n10_adj_3996), .I3(n30671), .O(n31081));
    defparam i7_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1033 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[17] [0]), .I3(n28732), .O(n30658));
    defparam i3_4_lut_adj_1033.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1034 (.I0(\data_in_frame[21] [0]), .I1(n12_adj_3998), 
            .I2(n16323), .I3(n31836), .O(n32679));
    defparam i6_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n31129));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i17148_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n32040), .I3(GND_net), .O(n18092));
    defparam i17148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1036 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[19] [5]), .O(n8_adj_3999));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1037 (.I0(\data_in_frame[19] [4]), .I1(n8_adj_3999), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [1]), .O(Kp_23__N_652));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[14] [2]), 
            .I2(\data_in_frame[12] [4]), .I3(\data_in_frame[14] [3]), .O(n60));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(Kp_23__N_1293), .I1(n31099), .I2(n31129), .I3(n31007), 
            .O(n58));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17145_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1]_c [2]), 
            .I2(n32040), .I3(GND_net), .O(n18093));
    defparam i17145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1266_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4752), .I3(GND_net), .O(n4754));
    defparam mux_1266_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_4_lut_adj_1038 (.I0(n30793), .I1(\data_in_frame[13] [2]), 
            .I2(n30752), .I3(\data_in_frame[16] [2]), .O(n59));
    defparam i23_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i13598_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n18178));
    defparam i13598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21_4_lut_adj_1039 (.I0(n30761), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[16] [5]), .I3(\data_in_frame[14] [7]), .O(n57));
    defparam i21_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1040 (.I0(n31070), .I1(n31132), .I2(\data_in_frame[12] [0]), 
            .I3(n31019), .O(n56));
    defparam i20_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1041 (.I0(n30809), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[14] [5]), .I3(n31123), .O(n55));
    defparam i19_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_1042 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[11] [0]), 
            .I2(n16963), .I3(\data_in_frame[9] [6]), .O(n63_adj_4000));
    defparam i27_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut_adj_1043 (.I0(\data_in_frame[11] [2]), .I1(n31028), 
            .I2(n31117), .I3(n30960), .O(n62));
    defparam i26_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i32_3_lut (.I0(n63_adj_4000), .I1(n55), .I2(n56), .I3(GND_net), 
            .O(n68));
    defparam i32_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(\data_in_frame[15] [4]), .I1(n30995), .I2(n17656), 
            .I3(n16657), .O(n61));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n57), .I1(n59), .I2(n58), .I3(n60), .O(n69));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n69), .I1(n61), .I2(n68), .I3(n62), .O(n32512));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30700));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1045 (.I0(n16978), .I1(n28791), .I2(\data_in_frame[18] [1]), 
            .I3(\data_in_frame[18] [5]), .O(n28_adj_4001));
    defparam i12_4_lut_adj_1045.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1046 (.I0(n31081), .I1(n28650), .I2(n30684), 
            .I3(n32512), .O(n26_adj_4002));
    defparam i10_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1047 (.I0(n31120), .I1(n30700), .I2(n30960), 
            .I3(n30658), .O(n27_adj_4003));
    defparam i11_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1048 (.I0(\data_in_frame[17] [7]), .I1(n30866), 
            .I2(\data_in_frame[18] [4]), .I3(n28673), .O(n25_adj_4004));
    defparam i9_4_lut_adj_1048.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1049 (.I0(n25_adj_4004), .I1(n27_adj_4003), .I2(n26_adj_4002), 
            .I3(n28_adj_4001), .O(n32292));
    defparam i15_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(n16895), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30611));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1051 (.I0(n30592), .I1(n30611), .I2(n27501), 
            .I3(\data_in_frame[8] [4]), .O(n12_adj_4005));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1052 (.I0(n16927), .I1(n12_adj_4005), .I2(n30935), 
            .I3(\data_in_frame[8] [0]), .O(n32560));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1053 (.I0(\data_in_frame[12] [0]), .I1(n27776), 
            .I2(\data_in_frame[11] [7]), .I3(n32560), .O(n31043));
    defparam i3_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1054 (.I0(\data_in_frame[9] [2]), .I1(n30896), 
            .I2(n27688), .I3(n28614), .O(n12_adj_4006));
    defparam i5_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1055 (.I0(\data_in_frame[11] [5]), .I1(n12_adj_4006), 
            .I2(n31043), .I3(\data_in_frame[13] [7]), .O(n16242));
    defparam i6_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1056 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[14] [1]), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n30752));
    defparam i2_3_lut_adj_1056.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1057 (.I0(n32292), .I1(n30720), .I2(Kp_23__N_652), 
            .I3(GND_net), .O(n30978));
    defparam i2_3_lut_adj_1057.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1058 (.I0(n30752), .I1(n16242), .I2(\data_in_frame[18] [5]), 
            .I3(n28756), .O(n32366));
    defparam i3_4_lut_adj_1058.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1059 (.I0(\data_in_frame[11] [1]), .I1(n17312), 
            .I2(n17529), .I3(\data_in_frame[15] [4]), .O(n30732));
    defparam i3_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1060 (.I0(Kp_23__N_1097), .I1(\data_in_frame[15] [3]), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[13] [1]), .O(n31007));
    defparam i3_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1061 (.I0(n16607), .I1(n14151), .I2(n31_adj_4007), 
            .I3(GND_net), .O(n32040));
    defparam i2_3_lut_adj_1061.LUT_INIT = 16'hfefe;
    SB_LUT4 i17153_3_lut (.I0(control_mode_c[1]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n32040), .I3(GND_net), .O(n18094));
    defparam i17153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[11] [2]), .I1(n30592), 
            .I2(GND_net), .I3(GND_net), .O(n16785));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1063 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[16] [0]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n31099));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(n28088), .I1(n17350), .I2(GND_net), 
            .I3(GND_net), .O(n28614));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1065 (.I0(\data_in_frame[18] [0]), .I1(n31099), 
            .I2(n31087), .I3(n30533), .O(n13_adj_4008));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1066 (.I0(n13_adj_4008), .I1(n11_adj_4009), .I2(\data_in_frame[11] [4]), 
            .I3(n28787), .O(n30720));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1066.LUT_INIT = 16'h9669;
    SB_LUT4 i13599_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n18179));
    defparam i13599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1067 (.I0(\data_in_frame[13] [3]), .I1(n17378), 
            .I2(n30732), .I3(GND_net), .O(n14_adj_4010));
    defparam i5_3_lut_adj_1067.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1068 (.I0(n31007), .I1(\data_in_frame[17] [5]), 
            .I2(n16686), .I3(n30787), .O(n15_adj_4011));
    defparam i6_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1069 (.I0(n15_adj_4011), .I1(n16785), .I2(n14_adj_4010), 
            .I3(n17252), .O(n28791));
    defparam i8_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18110));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3407[0]), .C(clk32MHz), 
            .D(n3276[0]), .R(n31148));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1070 (.I0(n30849), .I1(n30902), .I2(\data_in_frame[13] [0]), 
            .I3(GND_net), .O(n30793));
    defparam i2_3_lut_adj_1070.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17529));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n31132));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[10] [3]), .I1(n17356), 
            .I2(GND_net), .I3(GND_net), .O(n16657));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1074 (.I0(n15030), .I1(\data_in_frame[10] [7]), 
            .I2(n17297), .I3(\data_in_frame[13] [1]), .O(n14_adj_4012));
    defparam i6_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1075 (.I0(n30620), .I1(n14_adj_4012), .I2(n10_adj_4013), 
            .I3(\data_in_frame[17] [3]), .O(n30764));
    defparam i7_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1076 (.I0(Kp_23__N_1076), .I1(n30793), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[10] [6]), .O(n12_adj_4014));
    defparam i5_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1077 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_4014), 
            .I2(n31010), .I3(n17378), .O(n31815));
    defparam i6_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(n31815), .I1(n30764), .I2(GND_net), 
            .I3(GND_net), .O(n28673));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h9999;
    SB_LUT4 i28893_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n31148), .I2(n22632), 
            .I3(GND_net), .O(n31472));
    defparam i28893_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i29248_4_lut (.I0(n31148), .I1(\FRAME_MATCHER.state[3] ), .I2(n4854), 
            .I3(n4922), .O(n31272));
    defparam i29248_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(n28125), .I1(n30767), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1082));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i28763_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4854));   // verilog/coms.v(145[4] 299[11])
    defparam i28763_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[9] [7]), 
            .I2(n31028), .I3(GND_net), .O(n8_adj_4015));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(Kp_23__N_1082), .I1(n30857), .I2(n8_adj_4015), 
            .I3(n28088), .O(n31013));
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(\data_in_frame[14] [3]), .I1(n30796), 
            .I2(n31013), .I3(\data_in_frame[12] [2]), .O(n28756));
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n31126));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1083 (.I0(\data_in_frame[18] [7]), .I1(n30559), 
            .I2(\data_in_frame[14] [5]), .I3(n17114), .O(n31120));
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1084 (.I0(n31120), .I1(n31126), .I2(n28756), 
            .I3(GND_net), .O(n30963));
    defparam i2_3_lut_adj_1084.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17656));
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16686));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(Kp_23__N_986), .I1(n5_c), .I2(GND_net), 
            .I3(GND_net), .O(n17312));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1088 (.I0(\data_in_frame[8] [6]), .I1(n8), .I2(GND_net), 
            .I3(GND_net), .O(n16937));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1089 (.I0(n10_c), .I1(n16895), .I2(GND_net), 
            .I3(GND_net), .O(n31019));
    defparam i1_2_lut_adj_1089.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(n28088), .I1(n16954), .I2(GND_net), 
            .I3(GND_net), .O(n28603));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(n16954), .I1(n30767), .I2(GND_net), 
            .I3(GND_net), .O(n30769));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1092 (.I0(n31019), .I1(n16963), .I2(n16937), 
            .I3(n30852), .O(n15_adj_4016));
    defparam i6_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1093 (.I0(n15_adj_4016), .I1(n17350), .I2(n14_adj_4017), 
            .I3(n17312), .O(n27739));
    defparam i8_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n17350), .I1(n16895), .I2(GND_net), 
            .I3(GND_net), .O(n17642));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(n10_c), .I1(\data_in_frame[9] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n30866));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1096 (.I0(n17642), .I1(n27739), .I2(n30769), 
            .I3(n28603), .O(n30787));
    defparam i3_4_lut_adj_1096.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_in_frame[10] [7]), .I1(n30787), 
            .I2(GND_net), .I3(GND_net), .O(n28650));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1098 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[13] [3]), 
            .I2(\data_in_frame[11] [1]), .I3(\data_in_frame[15] [7]), .O(n24_adj_4018));
    defparam i10_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1099 (.I0(n30533), .I1(n28650), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[9] [1]), .O(n22_adj_4019));
    defparam i8_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1100 (.I0(\data_in_frame[13] [4]), .I1(n24_adj_4018), 
            .I2(n18_adj_3983), .I3(n17350), .O(n26_adj_4020));
    defparam i12_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1101 (.I0(\data_in_frame[17] [7]), .I1(n26_adj_4020), 
            .I2(n22_adj_4019), .I3(\data_in_frame[16] [0]), .O(n30958));
    defparam i13_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16927));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30902));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1104 (.I0(n28125), .I1(n16882), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n8_adj_4021));
    defparam i3_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1105 (.I0(\data_in_frame[10] [1]), .I1(n15023), 
            .I2(n8_adj_4021), .I3(\data_in_frame[9] [7]), .O(n30796));
    defparam i1_4_lut_adj_1105.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17297));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1107 (.I0(\data_in_frame[12] [3]), .I1(n30796), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n30559));
    defparam i2_3_lut_adj_1107.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1108 (.I0(n4_c), .I1(n5_c), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1076));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1109 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n30761));
    defparam i2_3_lut_adj_1109.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n17751), .D(n8825[2]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1110 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[10] [5]), 
            .I2(n30559), .I3(n17297), .O(n14_adj_4022));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1111 (.I0(\data_in_frame[17] [1]), .I1(n14_adj_4022), 
            .I2(n10_adj_4023), .I3(n30902), .O(n30684));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1097));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1112 (.I0(n30666), .I1(n30935), .I2(\data_in_frame[1]_c [3]), 
            .I3(GND_net), .O(n15023));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1112.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1113 (.I0(n17481), .I1(n15023), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n15030));
    defparam i2_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[10] [3]), .I1(n15030), 
            .I2(GND_net), .I3(GND_net), .O(n17114));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_CARRY add_43_4 (.CI(n25555), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n25556));
    SB_LUT4 i5_4_lut_adj_1115 (.I0(n30655), .I1(n30666), .I2(n30852), 
            .I3(n17636), .O(n12_adj_4024));
    defparam i5_4_lut_adj_1115.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(\data_in_frame[3] [4]), .I1(n12_adj_4024), 
            .I2(n30745), .I3(\data_in_frame[1]_c [2]), .O(n28620));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1117 (.I0(n28620), .I1(\data_in_frame[10] [2]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n31010));
    defparam i2_4_lut_adj_1117.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30849));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(n27501), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27714));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_16__7__I_0_3896_2_lut (.I0(\data_in_frame[16] [7]), 
            .I1(\data_in_frame[16] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1293));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_16__7__I_0_3896_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(n30849), .I1(n17342), .I2(\data_in_frame[10] [4]), 
            .I3(n31010), .O(n10_adj_4025));
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1121 (.I0(n28732), .I1(\data_in_frame[17] [0]), 
            .I2(Kp_23__N_1293), .I3(n30995), .O(n10_adj_4026));
    defparam i4_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1122 (.I0(n28620), .I1(n30684), .I2(n10_adj_4026), 
            .I3(n30761), .O(n16323));
    defparam i1_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1123 (.I0(\data_in_frame[19] [2]), .I1(n30629), 
            .I2(n16323), .I3(\data_in_frame[21] [4]), .O(n32203));
    defparam i3_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_56_2_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36139));   // verilog/coms.v(85[17:28])
    defparam i1_rep_56_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1124 (.I0(\data_in_frame[18] [1]), .I1(n30958), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n8_adj_4027));
    defparam i3_3_lut_adj_1124.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1125 (.I0(\data_in_frame[21] [3]), .I1(n30963), 
            .I2(n30684), .I3(n36139), .O(n32739));
    defparam i3_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1126 (.I0(\data_in_frame[21] [7]), .I1(n30764), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3926));
    defparam i2_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1127 (.I0(\data_in_frame[21] [5]), .I1(n30629), 
            .I2(n28673), .I3(\data_in_frame[19] [4]), .O(n32209));
    defparam i3_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1128 (.I0(\data_in_frame[20] [1]), .I1(n30958), 
            .I2(n27881), .I3(GND_net), .O(n32713));
    defparam i2_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1129 (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4028));
    defparam i2_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1130 (.I0(n16978), .I1(\data_in_frame[20] [0]), 
            .I2(\data_in_frame[19] [6]), .I3(n31073), .O(n10_adj_4029));
    defparam i4_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1131 (.I0(n32366), .I1(n30978), .I2(\data_in_frame[19] [0]), 
            .I3(\data_in_frame[20] [7]), .O(n32875));
    defparam i3_4_lut_adj_1131.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1132 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[20] [4]), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n6_adj_4030));
    defparam i2_3_lut_adj_1132.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(n7_adj_4028), .I1(n16978), .I2(\data_in_frame[21] [6]), 
            .I3(n31815), .O(n32519));
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h9669;
    SB_LUT4 i26912_4_lut (.I0(\data_in_frame[21] [2]), .I1(n32203), .I2(n30955), 
            .I3(\data_in_frame[19] [1]), .O(n33080));
    defparam i26912_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i6_4_lut_adj_1134 (.I0(\data_in_frame[20] [3]), .I1(n32739), 
            .I2(n8_adj_4027), .I3(n31776), .O(n22_adj_4031));
    defparam i6_4_lut_adj_1134.LUT_INIT = 16'h7bb7;
    SB_LUT4 i26914_4_lut (.I0(n32519), .I1(Kp_23__N_1591), .I2(n6_adj_4030), 
            .I3(n31776), .O(n33082));
    defparam i26914_4_lut.LUT_INIT = 16'h2882;
    SB_LUT4 i5_4_lut_adj_1135 (.I0(n28791), .I1(n32875), .I2(n10_adj_4029), 
            .I3(n27881), .O(n21));
    defparam i5_4_lut_adj_1135.LUT_INIT = 16'hedde;
    SB_LUT4 i13600_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n18180));
    defparam i13600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_2_lut_4_lut (.I0(n30489), .I1(n30879), .I2(\data_out_frame[5] [4]), 
            .I3(n31004), .O(n9));   // verilog/coms.v(71[16:27])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26916_4_lut (.I0(n32209), .I1(n30963), .I2(n30978), .I3(\data_in_frame[21] [1]), 
            .O(n33084));
    defparam i26916_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1136 (.I0(n32713), .I1(n32366), .I2(n30595), 
            .I3(\data_in_frame[20] [6]), .O(n19_adj_4032));
    defparam i3_4_lut_adj_1136.LUT_INIT = 16'h7dd7;
    SB_LUT4 i14_4_lut_adj_1137 (.I0(n21), .I1(n33082), .I2(n22_adj_4031), 
            .I3(n33080), .O(n30_adj_4033));
    defparam i14_4_lut_adj_1137.LUT_INIT = 16'hfbff;
    SB_LUT4 i9_4_lut_adj_1138 (.I0(n32679), .I1(n32357), .I2(n32882), 
            .I3(n32133), .O(n25_adj_4034));
    defparam i9_4_lut_adj_1138.LUT_INIT = 16'hfffb;
    SB_LUT4 i15_4_lut_adj_1139 (.I0(n25_adj_4034), .I1(n30_adj_4033), .I2(n19_adj_4032), 
            .I3(n33084), .O(n31_adj_4007));
    defparam i15_4_lut_adj_1139.LUT_INIT = 16'hfeff;
    SB_LUT4 i13601_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n18181));
    defparam i13601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n17773), .D(n4753));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13602_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30468), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n18182));
    defparam i13602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13587_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n18167));
    defparam i13587_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13588_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n18168));
    defparam i13588_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13589_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n18169));
    defparam i13589_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13590_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n18170));
    defparam i13590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18108));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13591_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n18171));
    defparam i13591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n17751), .D(n8825[1]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18107));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13592_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n18172));
    defparam i13592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13593_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n18173));
    defparam i13593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13594_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30451), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n18174));
    defparam i13594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17391));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_33_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n25584), .O(n2_adj_4036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n25613), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n31064));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1142 (.I0(n17391), .I1(n30920), .I2(n30790), 
            .I3(\data_in_frame[5] [7]), .O(n16882));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1143 (.I0(n16882), .I1(n30569), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n17481));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(n30923), .I1(n31064), .I2(n30537), 
            .I3(GND_net), .O(n10_c));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1145 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[8] [5]), .I3(n30496), .O(n10_adj_4037));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4038));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4039));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28171_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34084));
    defparam i28171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28175_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34083));
    defparam i28175_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4040));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4041));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28177_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34081));
    defparam i28177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28179_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34080));
    defparam i28179_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4042));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5]_c [0]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4043));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'ha300;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4044));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4045));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut (.I0(n5_adj_4044), 
            .I1(n6_adj_4043), .I2(n33932), .I3(GND_net), .O(n7_adj_4046));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28182_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34078));
    defparam i28182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1860170_i1_3_lut (.I0(n35618), .I1(n35606), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4047));
    defparam i1860170_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28184_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34077));
    defparam i28184_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28174_2_lut (.I0(n35690), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34085));
    defparam i28174_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4048));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4049));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28186_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34075));
    defparam i28186_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28188_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34074));
    defparam i28188_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4050));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_3_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n25554), .O(n2_adj_4051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n25583), .O(n2_adj_4052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4053));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28191_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34072));
    defparam i28191_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28194_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34071));
    defparam i28194_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_32 (.CI(n25583), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n25584));
    SB_LUT4 i4_4_lut_adj_1146 (.I0(\data_in_frame[5] [3]), .I1(n17134), 
            .I2(\data_in_frame[5] [2]), .I3(n30755), .O(n10_adj_4054));
    defparam i4_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1147 (.I0(n17452), .I1(n10_adj_4054), .I2(\data_in_frame[7] [4]), 
            .I3(GND_net), .O(n30614));
    defparam i5_3_lut_adj_1147.LUT_INIT = 16'h9696;
    SB_LUT4 i27019_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n33191));
    defparam i27019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27020_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n33192));
    defparam i27020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4055));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4056));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1148 (.I0(\data_in_frame[7] [2]), .I1(n17452), 
            .I2(n30952), .I3(n6_adj_4057), .O(n17350));
    defparam i4_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i28196_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34069));
    defparam i28196_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i27011_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n33183));
    defparam i27011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27010_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n33182));
    defparam i27010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28215_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34068));
    defparam i28215_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1149 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[8] [7]), 
            .I2(n16910), .I3(n30556), .O(n10_adj_4058));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1150 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n17265), .I3(n6_adj_4059), .O(n28125));
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_31_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n25582), .O(n2_adj_4060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28203_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n34376));   // verilog/coms.v(106[34:55])
    defparam i28203_2_lut.LUT_INIT = 16'hdddd;
    SB_CARRY add_43_31 (.CI(n25582), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n25583));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4061));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4062));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n17315));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4063));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_3 (.CI(n25554), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n25555));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_4_lut (.I0(n5_adj_4061), 
            .I1(n34376), .I2(n33932), .I3(byte_transmit_counter[0]), .O(n7_adj_4064));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i4_4_lut_adj_1152 (.I0(\data_in_frame[3] [7]), .I1(n16840), 
            .I2(n17315), .I3(n6_adj_4065), .O(n30569));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i1853738_i1_3_lut (.I0(n35576), .I1(n35570), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4066));
    defparam i1853738_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28216_2_lut (.I0(n35642), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34063));
    defparam i28216_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28197_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n34370));   // verilog/coms.v(106[34:55])
    defparam i28197_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4067));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13571_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n18151));
    defparam i13571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_4_lut (.I0(n5_adj_4067), 
            .I1(n34370), .I2(n33932), .I3(byte_transmit_counter[0]), .O(n7_adj_4069));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i1854341_i1_3_lut (.I0(n35552), .I1(n35624), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4070));
    defparam i1854341_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13572_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18152));
    defparam i13572_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28205_2_lut (.I0(n35648), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34066));
    defparam i28205_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_30_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n25581), .O(n2_adj_4071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n25612), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_8 (.CI(n25612), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n25613));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n25611), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_30 (.CI(n25581), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n25582));
    SB_LUT4 i4_4_lut_adj_1153 (.I0(n16863), .I1(n17315), .I2(\data_in_frame[1][7] ), 
            .I3(n6_adj_4072), .O(n17342));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n34364));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4073));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_4_lut (.I0(n5_adj_4073), 
            .I1(byte_transmit_counter[0]), .I2(n33932), .I3(n34364), .O(n7_adj_4074));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i28202_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34065));
    defparam i28202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_43_29_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n25580), .O(n2_adj_4075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28206_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34064));
    defparam i28206_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1854944_i1_3_lut (.I0(n35612), .I1(n35546), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4076));
    defparam i1854944_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28199_2_lut (.I0(n35660), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34070));
    defparam i28199_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_adj_1154 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4077));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4078));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n30652), .I1(n17277), .I2(n16714), 
            .I3(\data_in_frame[7] [0]), .O(n14_adj_4079));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_7 (.CI(n25611), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n25612));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4080));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4081));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut (.I0(n5_adj_4081), 
            .I1(n6_adj_4078), .I2(n33932), .I3(GND_net), .O(n7_adj_4082));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(n17290), .I1(n14_adj_4079), .I2(n10_adj_4077), 
            .I3(\data_in_frame[6] [6]), .O(n16895));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i13573_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18153));
    defparam i13573_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1157 (.I0(n17342), .I1(n30569), .I2(\data_in_frame[8] [3]), 
            .I3(GND_net), .O(n4_c));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4083));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30981));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i28096_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34087));
    defparam i28096_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28092_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n34086));
    defparam i28092_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1159 (.I0(\data_in_frame[18] [3]), .I1(n30595), 
            .I2(Kp_23__N_1591), .I3(\data_in_frame[20] [5]), .O(n32133));   // verilog/coms.v(268[9:85])
    defparam i3_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_855));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1855547_i1_3_lut (.I0(n35516), .I1(n35504), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4084));
    defparam i1855547_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_29 (.CI(n25580), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n25581));
    SB_LUT4 i28193_2_lut (.I0(n35666), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34073));
    defparam i28193_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_in_frame[4] [7]), .I1(n30587), 
            .I2(GND_net), .I3(GND_net), .O(n30923));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1161 (.I0(n17134), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_779), .I3(GND_net), .O(n17135));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(\data_in_frame[5] [1]), .I1(n17135), 
            .I2(\data_in_frame[5] [2]), .I3(n30923), .O(n10_adj_4085));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1163 (.I0(\data_in_frame[3] [1]), .I1(n10_adj_4085), 
            .I2(\data_in_frame[7] [3]), .I3(GND_net), .O(n28088));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4086));
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1165 (.I0(n30790), .I1(Kp_23__N_855), .I2(n30840), 
            .I3(n6_adj_4086), .O(n30852));
    defparam i4_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_28_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n25579), .O(n2_adj_4087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_in_frame[8] [1]), .I1(n27737), 
            .I2(GND_net), .I3(GND_net), .O(n30745));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1167 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1] [5]), 
            .I2(Kp_23__N_784), .I3(n6_adj_4088), .O(Kp_23__N_884));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[6] [2]), .I3(GND_net), .O(n30566));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16910));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1170 (.I0(\data_in_frame[6] [4]), .I1(n30913), 
            .I2(\data_in_frame[6] [2]), .I3(\data_in_frame[6] [0]), .O(n31058));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n25610), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13574_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18154));
    defparam i13574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30952));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1172 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3] [7]), .I3(GND_net), .O(n30831));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n30604));
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i13575_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n18155));
    defparam i13575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1174 (.I0(\data_in_frame[5] [4]), .I1(n30755), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n16730));
    defparam i2_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n17290));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30512));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4089));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\data_in_frame[2] [1]), .I1(n17290), 
            .I2(GND_net), .I3(GND_net), .O(n16832));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30572));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_CARRY add_43_28 (.CI(n25579), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n25580));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4090));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut (.I0(n5_adj_4090), 
            .I1(n6_adj_4089), .I2(n33932), .I3(GND_net), .O(n7_adj_4091));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut.LUT_INIT = 16'hacac;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n29939), .S(n29967));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16863));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n29935), .S(n29969));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_6 (.CI(n25610), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n25611));
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n29931), .S(n29971));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1]_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30584));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n25609), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n29927), .S(n29973));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n30920));   // verilog/coms.v(96[12:25])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n29923), .S(n29975));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_784));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n29919), .S(n29977));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n29915), .S(n29979));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n29911), .S(n29981));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n29907), .S(n29983));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n29903), .S(n29985));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n21837), .S(n29987));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1182 (.I0(Kp_23__N_784), .I1(n30920), .I2(n30584), 
            .I3(\data_in_frame[1]_c [1]), .O(Kp_23__N_779));   // verilog/coms.v(96[12:25])
    defparam i3_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30725));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n29899), .S(n29989));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n29895), .S(n29991));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_5 (.CI(n25609), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n25610));
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n29891), .S(n29993));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n29887), .S(n29995));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n29883), .S(n29997));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1856150_i1_3_lut (.I0(n35510), .I1(n35654), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4092));
    defparam i1856150_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n29879), .S(n29999));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n29875), .S(n30001));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n29871), .S(n30003));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n29867), .S(n30005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n29863), .S(n30007));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n29859), .S(n30009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n29855), .S(n30011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n29851), .S(n30013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n29847), .S(n30015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n29843), .S(n30017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n29841), .S(n30019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n29839), .S(n29837));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1184 (.I0(\data_in_frame[1]_c [0]), .I1(Kp_23__N_779), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n15796));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n29835), .S(n29945));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28187_2_lut (.I0(n35672), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34076));
    defparam i28187_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1185 (.I0(n15796), .I1(n30587), .I2(\data_in_frame[2] [7]), 
            .I3(GND_net), .O(n31067));
    defparam i2_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_4093));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha003;
    SB_LUT4 add_43_27_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n25578), .O(n2_adj_4094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n31055));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4095));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut (.I0(n5_adj_4095), 
            .I1(n6_adj_4093), .I2(n33932), .I3(GND_net), .O(n7_adj_4096));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n25608), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_27 (.CI(n25578), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n25579));
    SB_CARRY add_3971_4 (.CI(n25608), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n25609));
    SB_LUT4 i1_2_lut_adj_1187 (.I0(n30537), .I1(n31058), .I2(GND_net), 
            .I3(GND_net), .O(n30896));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1188 (.I0(\data_in_frame[4] [6]), .I1(n30932), 
            .I2(n16840), .I3(\data_in_frame[4] [0]), .O(n28_adj_4097));
    defparam i10_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i13576_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n18156));
    defparam i13576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1189 (.I0(\data_in_frame[0] [1]), .I1(n17277), 
            .I2(n31067), .I3(GND_net), .O(n14_adj_4098));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_1189.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_26_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n25577), .O(n2_adj_4099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n25577), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n25578));
    SB_LUT4 i6_4_lut_adj_1190 (.I0(\data_in_frame[0] [6]), .I1(n16863), 
            .I2(n30926), .I3(n30572), .O(n15_adj_4100));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1191 (.I0(n15_adj_4100), .I1(\data_in_frame[0] [7]), 
            .I2(n14_adj_4098), .I3(n30512), .O(n32550));   // verilog/coms.v(70[16:27])
    defparam i8_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i14_3_lut (.I0(\data_in_frame[4] [7]), .I1(n28_adj_4097), .I2(n16730), 
            .I3(GND_net), .O(n32_adj_4101));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i28183_2_lut (.I0(n35678), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34079));
    defparam i28183_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1192 (.I0(n32550), .I1(n30831), .I2(n30952), 
            .I3(n30601), .O(n30_adj_4102));
    defparam i12_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i13577_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n18157));
    defparam i13577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1193 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[5] [2]), .O(n31_adj_4103));
    defparam i13_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i27748_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n33932));   // verilog/coms.v(106[34:55])
    defparam i27748_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_4_lut_adj_1194 (.I0(Kp_23__N_811), .I1(\data_in_frame[3] [4]), 
            .I2(n30604), .I3(\data_in_frame[4] [4]), .O(n29_adj_4104));
    defparam i11_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i28172_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5]_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34344));   // verilog/coms.v(106[34:55])
    defparam i28172_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i13578_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30468), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18158));
    defparam i13578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17_4_lut_adj_1195 (.I0(n29_adj_4104), .I1(n31_adj_4103), .I2(n30_adj_4102), 
            .I3(n32_adj_4101), .O(n27737));
    defparam i17_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4105));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n17807), .D(n32090));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[1]_c [1]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30601));   // verilog/coms.v(96[12:25])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_4_lut (.I0(n5_adj_4105), 
            .I1(n34344), .I2(n33932), .I3(byte_transmit_counter[0]), .O(n7_adj_4106));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n25607), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13563_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n18143));
    defparam i13563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1197 (.I0(\data_in_frame[7] [7]), .I1(n16999), 
            .I2(n17265), .I3(\data_in_frame[5] [5]), .O(n30935));   // verilog/coms.v(75[16:27])
    defparam i1_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1858361_i1_3_lut (.I0(n35564), .I1(n35558), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4107));
    defparam i1858361_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1198 (.I0(\data_in_frame[2] [0]), .I1(n30725), 
            .I2(\data_in_frame[6] [5]), .I3(n16832), .O(n12_adj_4108));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i28178_2_lut (.I0(n35684), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n34082));
    defparam i28178_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1199 (.I0(\data_in_frame[4] [4]), .I1(n12_adj_4108), 
            .I2(n30981), .I3(\data_in_frame[1][6] ), .O(Kp_23__N_986));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1200 (.I0(Kp_23__N_986), .I1(n30840), .I2(\data_in_frame[8] [6]), 
            .I3(n30935), .O(n24));
    defparam i8_4_lut_adj_1200.LUT_INIT = 16'hde7b;
    SB_LUT4 i7_4_lut_adj_1201 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[6] [3]), 
            .I2(n30566), .I3(n27776), .O(n18_adj_4109));
    defparam i7_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1202 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16));
    defparam i5_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1203 (.I0(\data_in_frame[1]_c [3]), .I1(n18_adj_4109), 
            .I2(n30496), .I3(n31055), .O(n20));
    defparam i9_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i13564_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n18144));
    defparam i13564_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_3971_3 (.CI(n25607), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n25608));
    SB_LUT4 add_43_25_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n25576), .O(n2_adj_4110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3304), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3304), 
            .CO(n25607));
    SB_LUT4 i13565_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n18145));
    defparam i13565_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13566_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n18146));
    defparam i13566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13567_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n18147));
    defparam i13567_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n17807), .D(n32617));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13568_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n18148));
    defparam i13568_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n17807), .D(n31607));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n17807), .D(n30542));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n17807), .D(n32125));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n17807), .D(n31666));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n17807), .D(n30861));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n17807), .D(n32161));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n17807), .D(n31697));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n17807), .D(n32219));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n17807), .D(n32412));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n17807), .D(n31422));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n17807), .D(n31772));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n17807), .D(n32037));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n17807), .D(n31747));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n17807), .D(n32377));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4036), .S(n3_adj_4111));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13569_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n18149));
    defparam i13569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13570_3_lut_4_lut (.I0(n21993), .I1(n30468), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n18150));
    defparam i13570_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13555_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18135));
    defparam i13555_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13556_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18136));
    defparam i13556_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_25 (.CI(n25576), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n25577));
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4052), .S(n3_adj_4113));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4060), .S(n3_adj_4114));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4071), .S(n3_adj_4115));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4075), .S(n3_adj_4116));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4087), .S(n3_adj_4117));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4094), .S(n3_adj_4118));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4099), .S(n3_adj_4119));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4110), .S(n3_adj_4120));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4121), .S(n3_adj_4122));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4123), .S(n3_adj_4124));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_24_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n25575), .O(n2_adj_4121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n25575), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n25576));
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4125), .S(n3_adj_4126));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4127), .S(n3_adj_4128));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4129), .S(n3_adj_4130));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4131), .S(n3_adj_4132));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4133), .S(n3_adj_4134));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4135), .S(n3_adj_4136));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4137), .S(n3_adj_4138));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4139), .S(n3_adj_4140));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4141), .S(n3_adj_4142));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4143), .S(n3_adj_4144));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4145), .S(n3_adj_4146));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4147), .S(n3_adj_4148));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4149), .S(n3_adj_4150));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4151), .S(n3_adj_4152));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4153), .S(n3_adj_4154));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4155), .S(n3_adj_4156));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4157), .S(n3_adj_4158));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4159), .S(n3_adj_4160));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4161), .S(n3_adj_4162));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1204 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[14] [4]), .I3(\data_out_frame[14] [3]), 
            .O(n16888));
    defparam i2_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_23_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n25574), .O(n2_adj_4123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4051), .S(n3_adj_4163));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_23 (.CI(n25574), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n25575));
    SB_LUT4 add_43_22_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n25573), .O(n2_adj_4125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13557_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18137));
    defparam i13557_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_22 (.CI(n25573), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n25574));
    SB_LUT4 add_43_21_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n25572), .O(n2_adj_4127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13558_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18138));
    defparam i13558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_21 (.CI(n25572), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n25573));
    SB_LUT4 add_43_20_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n25571), .O(n2_adj_4129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13559_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18139));
    defparam i13559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13560_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18140));
    defparam i13560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13561_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18141));
    defparam i13561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_20 (.CI(n25571), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n25572));
    SB_LUT4 add_43_19_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n25570), .O(n2_adj_4131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_19 (.CI(n25570), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n25571));
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n25554));
    SB_LUT4 add_43_18_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n25569), .O(n2_adj_4133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13562_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30455), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18142));
    defparam i13562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_18 (.CI(n25569), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n25570));
    SB_LUT4 i13547_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n18127));
    defparam i13547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18106));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13548_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n18128));
    defparam i13548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13549_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n18129));
    defparam i13549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13550_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n18130));
    defparam i13550_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13551_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n18131));
    defparam i13551_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13552_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n18132));
    defparam i13552_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13553_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n18133));
    defparam i13553_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18100));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_17_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n25568), .O(n2_adj_4135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13554_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30447), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n18134));
    defparam i13554_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1205 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4164));
    defparam i2_2_lut_adj_1205.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1206 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[1]_c [1]), .I3(\data_in_frame[3] [2]), .O(n30755));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [13]), .I3(\FRAME_MATCHER.state [14]), 
            .O(n14_adj_4165));
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_17 (.CI(n25568), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n25569));
    SB_LUT4 i7_4_lut_adj_1208 (.I0(\FRAME_MATCHER.state [15]), .I1(n14_adj_4165), 
            .I2(n10_adj_4164), .I3(\FRAME_MATCHER.state [11]), .O(n22829));
    defparam i7_4_lut_adj_1208.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1209 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[3] [0]), .I3(GND_net), .O(n30932));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_16_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n25567), .O(n2_adj_4137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n25567), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n25568));
    SB_LUT4 add_43_15_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n25566), .O(n2_adj_4139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_15 (.CI(n25566), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n25567));
    SB_LUT4 i2_3_lut_adj_1210 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n5_adj_3964));
    defparam i2_3_lut_adj_1210.LUT_INIT = 16'hfefe;
    SB_LUT4 i17414_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n21985));
    defparam i17414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1211 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n21985), .I3(byte_transmit_counter[2]), .O(n22775));
    defparam i2_4_lut_adj_1211.LUT_INIT = 16'h8880;
    SB_LUT4 i24996_3_lut (.I0(n22632), .I1(n16614), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n31148));
    defparam i24996_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n16714));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1213 (.I0(n22775), .I1(n22624), .I2(n21830), 
            .I3(n5_adj_3964), .O(n32888));
    defparam i3_4_lut_adj_1213.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_847_i1_3_lut (.I0(n32888), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n4922), .I3(GND_net), .O(n3276[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_847_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18098));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1214 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [6]), .O(n30587));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_14_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n25565), .O(n2_adj_4141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1215 (.I0(control_mode[2]), .I1(\control_mode[6] ), 
            .I2(\control_mode[7] ), .I3(\control_mode[4] ), .O(n10_adj_4166));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1215.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1216 (.I0(\control_mode[5] ), .I1(n10_adj_4166), 
            .I2(control_mode[3]), .I3(GND_net), .O(n21709));   // verilog/coms.v(127[12] 300[6])
    defparam i5_3_lut_adj_1216.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(control_mode_c[1]), .I1(n21710), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'hdddd;
    SB_LUT4 i12_4_lut_adj_1218 (.I0(\FRAME_MATCHER.state [31]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [24]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n28_adj_4168));
    defparam i12_4_lut_adj_1218.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_14 (.CI(n25565), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n25566));
    SB_LUT4 i2_3_lut_4_lut_adj_1219 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_884), 
            .I2(\data_in_frame[8] [4]), .I3(n17342), .O(n5_c));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i25083_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i25083_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1220 (.I0(control_mode_c[1]), .I1(n21709), .I2(control_mode_c[0]), 
            .I3(GND_net), .O(n15_adj_4));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_1220.LUT_INIT = 16'hefef;
    SB_LUT4 i17260_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3407[0]), .I2(GND_net), 
            .I3(GND_net), .O(n21830));
    defparam i17260_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n16619), .I1(n63_adj_3), .I2(GND_net), 
            .I3(GND_net), .O(n17965));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_884), 
            .I2(n10_adj_4037), .I3(n17277), .O(n17356));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1222 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [18]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n26_adj_4171));
    defparam i10_4_lut_adj_1222.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1223 (.I0(n16895), .I1(n30866), .I2(\data_in_frame[13] [6]), 
            .I3(\data_in_frame[11] [5]), .O(n30533));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_13_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n25564), .O(n2_adj_4143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_13 (.CI(n25564), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n25565));
    SB_LUT4 add_43_12_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n25563), .O(n2_adj_4145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11_4_lut_adj_1224 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [20]), 
            .I2(\FRAME_MATCHER.state [21]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n27_adj_4172));
    defparam i11_4_lut_adj_1224.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1225 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [22]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n25_adj_4173));
    defparam i9_4_lut_adj_1225.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n35456), .I2(n34082), .I3(byte_transmit_counter[4]), .O(n35729));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n35729_bdd_4_lut (.I0(n35729), .I1(n14_adj_4107), .I2(n7_adj_4106), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n35729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29507 (.I0(byte_transmit_counter[3]), 
            .I1(n35462), .I2(n34079), .I3(byte_transmit_counter[4]), .O(n35723));
    defparam byte_transmit_counter_3__bdd_4_lut_29507.LUT_INIT = 16'he4aa;
    SB_LUT4 n35723_bdd_4_lut (.I0(n35723), .I1(n35630), .I2(n7_adj_4096), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n35723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29502 (.I0(byte_transmit_counter[3]), 
            .I1(n35468), .I2(n34076), .I3(byte_transmit_counter[4]), .O(n35717));
    defparam byte_transmit_counter_3__bdd_4_lut_29502.LUT_INIT = 16'he4aa;
    SB_LUT4 n35717_bdd_4_lut (.I0(n35717), .I1(n14_adj_4092), .I2(n7_adj_4091), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n35717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15_4_lut_adj_1226 (.I0(n25_adj_4173), .I1(n27_adj_4172), .I2(n26_adj_4171), 
            .I3(n28_adj_4168), .O(n22967));
    defparam i15_4_lut_adj_1226.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_12 (.CI(n25563), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n25564));
    SB_LUT4 add_43_11_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n25562), .O(n2_adj_4147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n22634));
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'hfffe;
    SB_LUT4 i17252_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n21822));
    defparam i17252_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(n22634), .I1(n22967), .I2(n22829), 
            .I3(GND_net), .O(n16614));   // verilog/coms.v(254[5:25])
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1229 (.I0(\FRAME_MATCHER.state[3] ), .I1(n16614), 
            .I2(GND_net), .I3(GND_net), .O(n16429));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_adj_1229.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29497 (.I0(byte_transmit_counter[3]), 
            .I1(n35474), .I2(n34073), .I3(byte_transmit_counter[4]), .O(n35711));
    defparam byte_transmit_counter_3__bdd_4_lut_29497.LUT_INIT = 16'he4aa;
    SB_LUT4 n35711_bdd_4_lut (.I0(n35711), .I1(n14_adj_4084), .I2(n7_adj_4082), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n35711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16611));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'hbbbb;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29492 (.I0(byte_transmit_counter[3]), 
            .I1(n35480), .I2(n34070), .I3(byte_transmit_counter[4]), .O(n35705));
    defparam byte_transmit_counter_3__bdd_4_lut_29492.LUT_INIT = 16'he4aa;
    SB_LUT4 n35705_bdd_4_lut (.I0(n35705), .I1(n14_adj_4076), .I2(n7_adj_4074), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n35705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29487 (.I0(byte_transmit_counter[3]), 
            .I1(n35486), .I2(n34066), .I3(byte_transmit_counter[4]), .O(n35699));
    defparam byte_transmit_counter_3__bdd_4_lut_29487.LUT_INIT = 16'he4aa;
    SB_LUT4 n35699_bdd_4_lut (.I0(n35699), .I1(n14_adj_4070), .I2(n7_adj_4069), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n35699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29482 (.I0(byte_transmit_counter[3]), 
            .I1(n35492), .I2(n34063), .I3(byte_transmit_counter[4]), .O(n35693));
    defparam byte_transmit_counter_3__bdd_4_lut_29482.LUT_INIT = 16'he4aa;
    SB_LUT4 n35693_bdd_4_lut (.I0(n35693), .I1(n14_adj_4066), .I2(n7_adj_4064), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n35693_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n35687));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n35687_bdd_4_lut (.I0(n35687), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n35690));
    defparam n35687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29472 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n35681));
    defparam byte_transmit_counter_0__bdd_4_lut_29472.LUT_INIT = 16'he4aa;
    SB_LUT4 n35681_bdd_4_lut (.I0(n35681), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n35684));
    defparam n35681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_11 (.CI(n25562), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n25563));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29467 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n35675));
    defparam byte_transmit_counter_0__bdd_4_lut_29467.LUT_INIT = 16'he4aa;
    SB_LUT4 n35675_bdd_4_lut (.I0(n35675), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n35678));
    defparam n35675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29462 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n35669));
    defparam byte_transmit_counter_0__bdd_4_lut_29462.LUT_INIT = 16'he4aa;
    SB_LUT4 n35669_bdd_4_lut (.I0(n35669), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n35672));
    defparam n35669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29457 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n35663));
    defparam byte_transmit_counter_0__bdd_4_lut_29457.LUT_INIT = 16'he4aa;
    SB_LUT4 n35663_bdd_4_lut (.I0(n35663), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n35666));
    defparam n35663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29452 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n35657));
    defparam byte_transmit_counter_0__bdd_4_lut_29452.LUT_INIT = 16'he4aa;
    SB_LUT4 n35657_bdd_4_lut (.I0(n35657), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n35660));
    defparam n35657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29447 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n35651));
    defparam byte_transmit_counter_0__bdd_4_lut_29447.LUT_INIT = 16'he4aa;
    SB_LUT4 n35651_bdd_4_lut (.I0(n35651), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n35654));
    defparam n35651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29442 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n35645));
    defparam byte_transmit_counter_0__bdd_4_lut_29442.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1231 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[16] [6]), .I3(n28707), .O(n31096));
    defparam i2_3_lut_4_lut_adj_1231.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_10_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n25561), .O(n2_adj_4149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n35645_bdd_4_lut (.I0(n35645), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n35648));
    defparam n35645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29437 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n35639));
    defparam byte_transmit_counter_0__bdd_4_lut_29437.LUT_INIT = 16'he4aa;
    SB_LUT4 n35639_bdd_4_lut (.I0(n35639), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n35642));
    defparam n35639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n33182), .I2(n33183), .I3(byte_transmit_counter[2]), .O(n35627));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n35627_bdd_4_lut (.I0(n35627), .I1(n33192), .I2(n33191), .I3(byte_transmit_counter[2]), 
            .O(n35630));
    defparam n35627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29432 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n35621));
    defparam byte_transmit_counter_0__bdd_4_lut_29432.LUT_INIT = 16'he4aa;
    SB_LUT4 n35621_bdd_4_lut (.I0(n35621), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n35624));
    defparam n35621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29417 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n35615));
    defparam byte_transmit_counter_0__bdd_4_lut_29417.LUT_INIT = 16'he4aa;
    SB_LUT4 n35615_bdd_4_lut (.I0(n35615), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n35618));
    defparam n35615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[15] [7]), .I3(GND_net), .O(n30638));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_CARRY add_43_10 (.CI(n25561), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n25562));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29412 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n35609));
    defparam byte_transmit_counter_0__bdd_4_lut_29412.LUT_INIT = 16'he4aa;
    SB_LUT4 n35609_bdd_4_lut (.I0(n35609), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n35612));
    defparam n35609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29407 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n35603));
    defparam byte_transmit_counter_0__bdd_4_lut_29407.LUT_INIT = 16'he4aa;
    SB_LUT4 n35603_bdd_4_lut (.I0(n35603), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n35606));
    defparam n35603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_29477 (.I0(byte_transmit_counter[3]), 
            .I1(n35498), .I2(n34085), .I3(byte_transmit_counter[4]), .O(n35579));
    defparam byte_transmit_counter_3__bdd_4_lut_29477.LUT_INIT = 16'he4aa;
    SB_LUT4 n35579_bdd_4_lut (.I0(n35579), .I1(n14_adj_4047), .I2(n7_adj_4046), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n35579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29402 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n35573));
    defparam byte_transmit_counter_0__bdd_4_lut_29402.LUT_INIT = 16'he4aa;
    SB_LUT4 n35573_bdd_4_lut (.I0(n35573), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n35576));
    defparam n35573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29378 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n35567));
    defparam byte_transmit_counter_0__bdd_4_lut_29378.LUT_INIT = 16'he4aa;
    SB_LUT4 n35567_bdd_4_lut (.I0(n35567), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n35570));
    defparam n35567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29373 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n35561));
    defparam byte_transmit_counter_0__bdd_4_lut_29373.LUT_INIT = 16'he4aa;
    SB_LUT4 n35561_bdd_4_lut (.I0(n35561), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n35564));
    defparam n35561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29368 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n35555));
    defparam byte_transmit_counter_0__bdd_4_lut_29368.LUT_INIT = 16'he4aa;
    SB_LUT4 n35555_bdd_4_lut (.I0(n35555), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n35558));
    defparam n35555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29363 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n35549));
    defparam byte_transmit_counter_0__bdd_4_lut_29363.LUT_INIT = 16'he4aa;
    SB_LUT4 n35549_bdd_4_lut (.I0(n35549), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n35552));
    defparam n35549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29358 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n35543));
    defparam byte_transmit_counter_0__bdd_4_lut_29358.LUT_INIT = 16'he4aa;
    SB_LUT4 n35543_bdd_4_lut (.I0(n35543), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n35546));
    defparam n35543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_9_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n25560), .O(n2_adj_4151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n25560), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n25561));
    SB_LUT4 i1_2_lut_4_lut_adj_1233 (.I0(\data_in_frame[9] [0]), .I1(n27739), 
            .I2(n17356), .I3(Kp_23__N_1092), .O(n30767));
    defparam i1_2_lut_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1234 (.I0(\data_in_frame[9] [0]), .I1(n27739), 
            .I2(n17356), .I3(\data_in_frame[11] [7]), .O(n31028));
    defparam i1_2_lut_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1235 (.I0(n17356), .I1(n4_c), .I2(n28603), 
            .I3(n15030), .O(n14_adj_4017));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1236 (.I0(n17356), .I1(n4_c), .I2(\data_in_frame[12] [7]), 
            .I3(GND_net), .O(n17378));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29353 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n35513));
    defparam byte_transmit_counter_0__bdd_4_lut_29353.LUT_INIT = 16'he4aa;
    SB_LUT4 n35513_bdd_4_lut (.I0(n35513), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n35516));
    defparam n35513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_376_Select_1_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4163));
    defparam select_376_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_2_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4162));
    defparam select_376_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_1237 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[16] [2]), .I3(n17057), .O(n30562));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1238 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [6]), .I3(GND_net), .O(n9_adj_4174));
    defparam i1_2_lut_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_LUT4 select_376_Select_3_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4160));
    defparam select_376_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_1239 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[18] [4]), 
            .I2(n14898), .I3(\data_out_frame[23] [2]), .O(n30802));
    defparam i2_3_lut_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 select_376_Select_4_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4158));
    defparam select_376_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 add_43_8_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n25559), .O(n2_adj_4153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(\data_out_frame[23] [2]), .I1(n27823), 
            .I2(n31016), .I3(GND_net), .O(n6_adj_4175));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h9696;
    SB_CARRY add_43_8 (.CI(n25559), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n25560));
    SB_LUT4 select_376_Select_5_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4156));
    defparam select_376_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_6_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4154));
    defparam select_376_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_7_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4152));
    defparam select_376_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1241 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[25] [1]), 
            .I2(n2483), .I3(GND_net), .O(n6_adj_4176));
    defparam i1_2_lut_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_LUT4 select_376_Select_8_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4150));
    defparam select_376_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(n28791), .I1(n30720), .I2(\data_in_frame[19] [7]), 
            .I3(GND_net), .O(n27881));
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1243 (.I0(n28791), .I1(n30720), .I2(Kp_23__N_652), 
            .I3(n32292), .O(n31836));
    defparam i2_3_lut_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_7_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n25558), .O(n2_adj_4155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1244 (.I0(\data_out_frame[23] [0]), .I1(n16263), 
            .I2(n27823), .I3(GND_net), .O(n17262));
    defparam i1_2_lut_3_lut_adj_1244.LUT_INIT = 16'h9696;
    SB_LUT4 select_376_Select_9_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4148));
    defparam select_376_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_10_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4146));
    defparam select_376_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_11_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4144));
    defparam select_376_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i5_3_lut_4_lut_adj_1245 (.I0(n30737), .I1(\data_out_frame[15] [6]), 
            .I2(n28767), .I3(\data_out_frame[17] [6]), .O(n14_adj_4177));
    defparam i5_3_lut_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 select_376_Select_12_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4142));
    defparam select_376_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_13_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4140));
    defparam select_376_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_14_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4138));
    defparam select_376_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_15_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4136));
    defparam select_376_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_16_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4134));
    defparam select_376_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_17_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4132));
    defparam select_376_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_4_lut_adj_1246 (.I0(n16279), .I1(n28725), .I2(n10_adj_4178), 
            .I3(n28654), .O(n31034));
    defparam i1_2_lut_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(n21861), .I1(n10_adj_4179), .I2(GND_net), 
            .I3(GND_net), .O(n30463));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1248 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [4]), 
            .I2(n28088), .I3(n17350), .O(n17252));
    defparam i1_2_lut_3_lut_4_lut_adj_1248.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1249 (.I0(n28767), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n31025));
    defparam i1_2_lut_3_lut_adj_1249.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1250 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[17] [3]), .I3(GND_net), .O(n30739));
    defparam i1_2_lut_3_lut_adj_1250.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut (.I0(n28784), .I1(n28654), .I2(\data_out_frame[19] [3]), 
            .I3(GND_net), .O(n10_adj_4180));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_376_Select_18_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4130));
    defparam select_376_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1251 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[9] [6]), .I3(n30857), .O(Kp_23__N_1092));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 select_376_Select_19_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4128));
    defparam select_376_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1252 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(n16614), .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n16608));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1252.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1253 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(n16614), .I2(\FRAME_MATCHER.state [1]), .I3(n16611), .O(n16621));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1253.LUT_INIT = 16'hffef;
    SB_LUT4 select_376_Select_20_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4126));
    defparam select_376_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_21_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4124));
    defparam select_376_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_CARRY add_43_7 (.CI(n25558), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n25559));
    SB_LUT4 select_376_Select_22_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4122));
    defparam select_376_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18097));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n17751), .D(n8825[0]), .R(n17965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_376_Select_23_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4120));
    defparam select_376_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_24_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4119));
    defparam select_376_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_25_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4118));
    defparam select_376_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_26_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4117));
    defparam select_376_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_27_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4116));
    defparam select_376_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 add_43_4_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n25555), .O(n2_adj_4161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18095));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n31272), 
            .D(n4854), .R(n31472));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_376_Select_28_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4115));
    defparam select_376_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_29_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4114));
    defparam select_376_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_30_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4113));
    defparam select_376_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_DFF control_mode_i0_i1 (.Q(control_mode_c[1]), .C(clk32MHz), .D(n18094));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_376_Select_0_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_376_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_376_Select_31_i3_2_lut_4_lut (.I0(n22650), .I1(n16429), 
            .I2(n22632), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4111));
    defparam select_376_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_4_lut_adj_1254 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [2]), .I3(\data_out_frame[20] [1]), 
            .O(n30486));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1255 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n31052), .I3(n30799), .O(n27823));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1256 (.I0(\data_out_frame[14] [0]), .I1(n17600), 
            .I2(n16702), .I3(n30562), .O(n31052));
    defparam i2_3_lut_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_6_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n25557), .O(n2_adj_4157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n17773), .D(n4754));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(\data_out_frame[14] [0]), .I1(n17600), 
            .I2(\data_out_frame[13] [7]), .I3(GND_net), .O(n30770));
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1258 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[4] [6]), .O(n30652));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1259 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [3]), .I3(GND_net), .O(n16671));
    defparam i1_2_lut_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1260 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [5]), 
            .I2(n28699), .I3(n4_adj_4181), .O(n28702));
    defparam i1_2_lut_3_lut_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1261 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[1]_c [2]), .I3(n30655), .O(n16963));
    defparam i1_2_lut_3_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1262 (.I0(n16822), .I1(n28702), .I2(n30828), 
            .I3(n30860), .O(n32161));
    defparam i2_3_lut_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1263 (.I0(\data_in_frame[4] [5]), .I1(n16797), 
            .I2(\data_in_frame[2] [1]), .I3(n17290), .O(n30556));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n18093));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1264 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1]_c [3]), .I3(\data_in_frame[1]_c [2]), 
            .O(n30790));
    defparam i1_2_lut_3_lut_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1265 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n17290), .O(Kp_23__N_811));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1266 (.I0(n22650), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_4035), 
            .O(n30468));
    defparam i1_2_lut_3_lut_4_lut_adj_1266.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_4_lut_adj_1267 (.I0(n16822), .I1(n28702), .I2(n30575), 
            .I3(n31061), .O(n31666));
    defparam i2_3_lut_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1268 (.I0(\data_out_frame[18] [4]), .I1(n14898), 
            .I2(n28699), .I3(n16671), .O(n6_adj_4182));
    defparam i1_2_lut_3_lut_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1269 (.I0(\data_out_frame[20] [2]), .I1(n28622), 
            .I2(\data_out_frame[19] [7]), .I3(n30969), .O(n32847));
    defparam i2_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1270 (.I0(\data_out_frame[20] [2]), .I1(n28622), 
            .I2(\data_out_frame[20] [3]), .I3(n28667), .O(n2196));
    defparam i2_3_lut_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1271 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[11] [4]), .I3(n10_adj_3987), .O(n31073));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1272 (.I0(\data_out_frame[25] [1]), .I1(n10_adj_4183), 
            .I2(\data_out_frame[25] [4]), .I3(n31061), .O(n30828));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1273 (.I0(\data_out_frame[25] [1]), .I1(n10_adj_4183), 
            .I2(\data_out_frame[25] [4]), .I3(n30860), .O(n30861));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(n16895), .I1(n10_c), .I2(\data_in_frame[9] [2]), 
            .I3(\data_in_frame[11] [3]), .O(n11_adj_4009));   // verilog/coms.v(72[16:41])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1274 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_4112));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_adj_1274.LUT_INIT = 16'hfbfb;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n18092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(\control_mode[4] ), .C(clk32MHz), .D(n18091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(\control_mode[5] ), .C(clk32MHz), .D(n18090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk32MHz), .D(n18089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(\control_mode[7] ), .C(clk32MHz), .D(n18088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n35879));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1275 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[11] [4]), .I3(n16686), .O(n30960));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n17773), .D(n4755));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n17773), .D(n4756));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n17773), .D(n4757));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n17773), .D(n4758));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n17773), .D(n4759));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n17773), .D(n4760));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n17773), .D(n4761));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n17773), .D(n4762));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n17773), 
            .D(n4763));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n17773), 
            .D(n4764));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n17773), 
            .D(n4765));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n17773), 
            .D(n4766));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n17773), 
            .D(n4767));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n17773), 
            .D(n4768));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n17773), 
            .D(n4769));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n17773), 
            .D(n4770));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n17773), 
            .D(n4771));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n17773), 
            .D(n4772));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n17773), 
            .D(n4773));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n17773), 
            .D(n4774));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n17773), 
            .D(n4775));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n17773), 
            .D(n4776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n35882));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n30394), .D(n17937), 
            .R(n31439));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1276 (.I0(n28697), .I1(\data_out_frame[23] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(GND_net), .O(n6_adj_4184));
    defparam i1_2_lut_3_lut_adj_1276.LUT_INIT = 16'h9696;
    SB_LUT4 i17290_2_lut_3_lut (.I0(n22650), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n21861));
    defparam i17290_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1277 (.I0(n16606), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n16429), .O(n22650));
    defparam i2_3_lut_4_lut_adj_1277.LUT_INIT = 16'haa8a;
    SB_LUT4 i1_2_lut_3_lut_adj_1278 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n16604), .I3(GND_net), .O(n16606));   // verilog/coms.v(222[5:21])
    defparam i1_2_lut_3_lut_adj_1278.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1279 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n16614), .I3(GND_net), .O(n16604));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_adj_1279.LUT_INIT = 16'hfefe;
    SB_LUT4 i28784_3_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3407[0]), 
            .I2(n63_adj_3), .I3(n16619), .O(n17751));
    defparam i28784_3_lut_4_lut.LUT_INIT = 16'h0f1f;
    SB_LUT4 i1_2_lut_3_lut_adj_1280 (.I0(\FRAME_MATCHER.state[3] ), .I1(n16614), 
            .I2(n22624), .I3(GND_net), .O(n16619));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1280.LUT_INIT = 16'hefef;
    SB_LUT4 i5_3_lut_4_lut_adj_1281 (.I0(n16686), .I1(\data_in_frame[11] [4]), 
            .I2(n10_adj_3986), .I3(n30972), .O(n30595));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1282 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [2]), 
            .I2(n28610), .I3(n32564), .O(n31422));
    defparam i2_3_lut_4_lut_adj_1282.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_3_lut (.I0(n30684), .I1(n28791), .I2(n30955), .I3(GND_net), 
            .O(n12_adj_3998));
    defparam i5_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [2]), 
            .I2(n31084), .I3(n30643), .O(n8_adj_4185));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1283 (.I0(n31815), .I1(n30684), .I2(\data_in_frame[19] [3]), 
            .I3(GND_net), .O(n30629));
    defparam i1_2_lut_3_lut_adj_1283.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1284 (.I0(n31_adj_3932), .I1(n16608), .I2(n14151), 
            .I3(\FRAME_MATCHER.state [2]), .O(n32812));
    defparam i3_4_lut_adj_1284.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_4_lut (.I0(n30739), .I1(n31102), .I2(n31025), .I3(\data_out_frame[19] [7]), 
            .O(n27760));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29330 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n35507));
    defparam byte_transmit_counter_0__bdd_4_lut_29330.LUT_INIT = 16'he4aa;
    SB_LUT4 i18050_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n22624));
    defparam i18050_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1285 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n5019));
    defparam i1_2_lut_3_lut_adj_1285.LUT_INIT = 16'h0202;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n18536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n18535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n18534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n18533));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n18532));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n18531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n18530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n18529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n18528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n18527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n18526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n18525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n18524));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n18523));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n18522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n18521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n18520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n18519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n18518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n18517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n18516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n18515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n18514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n18513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n18512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n18511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n18510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n18509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n18508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n18507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n18506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n18505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n18504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n18503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n18502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n18501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n18500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n18499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n18498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n18497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n18496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n18495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n18494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n18493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n18492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n18491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n18490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n18489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n18485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n18484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n18483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n18482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n18481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n18480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n18479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n18478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n18477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n18476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n18475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n18474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n18473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n18472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n18471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n18470));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n18469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n18468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n18467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n18466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n18465));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n18464));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n18463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n18462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n18461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n18460));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n18459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n18458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n18457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n18456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n18455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n18454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n18453));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n18452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n18451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n18450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5]_c [0]), .C(clk32MHz), 
           .D(n18449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5]_c [1]), .C(clk32MHz), 
           .D(n18448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n18447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n18446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n18445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n18444));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5][6] ), .C(clk32MHz), 
           .D(n18443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5][7] ), .C(clk32MHz), 
           .D(n18442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n18441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n18440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n18439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n18438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n18437));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1286 (.I0(control_mode_c[0]), .I1(\control_mode[5] ), 
            .I2(n10_adj_4166), .I3(control_mode[3]), .O(n21710));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1286.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_6 (.CI(n25557), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n25558));
    SB_LUT4 i17154_3_lut (.I0(control_mode_c[0]), .I1(\data_in_frame[1]_c [0]), 
            .I2(n32040), .I3(GND_net), .O(n18054));
    defparam i17154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1287 (.I0(n27737), .I1(\data_in_frame[6] [3]), 
            .I2(n30537), .I3(n31058), .O(n30840));
    defparam i1_2_lut_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n18436));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1288 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[1]_c [2]), .I3(GND_net), .O(n16999));
    defparam i1_2_lut_3_lut_adj_1288.LUT_INIT = 16'h9696;
    SB_LUT4 n35507_bdd_4_lut (.I0(n35507), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n35510));
    defparam n35507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1289 (.I0(\data_in_frame[1]_c [2]), .I1(\data_in_frame[1]_c [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n17265));   // verilog/coms.v(96[12:25])
    defparam i2_3_lut_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i17398_2_lut_3_lut (.I0(n63_adj_3958), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));   // verilog/coms.v(157[6] 159[9])
    defparam i17398_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\data_in_frame[6] [3]), .I1(n30537), 
            .I2(n31058), .I3(GND_net), .O(n17636));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1291 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n16840));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1291.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n18435));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n18434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n18433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n18432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n18431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n18430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n18429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n18428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n18427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n18426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n18425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n18424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n18423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n18422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n18421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n18420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n18419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n18418));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n18417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n18416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n18415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n18414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n18413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n18412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n18411));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n18410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n18409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n18408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n18407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n18406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n18405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n18404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n18403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n18402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n18401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n18400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n18399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n18398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n18397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n18396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n18395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n18394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n18393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n18392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n18391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n18390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n18389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n18388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n18387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n18386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n18385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n18384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n18383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n18382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n18381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n18380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n18379));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n18378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n18377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n18376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n18375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n18374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n18373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n18372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n18371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n18370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n18369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n18368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n18367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n18366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n18365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n18364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n18363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n18362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n18361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n18360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n18359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n18358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n18357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n18356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n18355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n18354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n18353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n18352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n18351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n18350));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n17277));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1293 (.I0(n16797), .I1(\data_in_frame[2] [1]), 
            .I2(n17290), .I3(GND_net), .O(n30926));
    defparam i1_2_lut_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1294 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n16797));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n18349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n18348));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1295 (.I0(n16797), .I1(n17290), .I2(\data_in_frame[6] [7]), 
            .I3(\data_in_frame[4] [5]), .O(n30537));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n30913));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(Kp_23__N_884), .I1(\data_in_frame[8] [1]), 
            .I2(n27737), .I3(GND_net), .O(n27776));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1298 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[3] [7]), .O(n6_adj_4088));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1299 (.I0(\data_in_frame[1]_c [0]), .I1(Kp_23__N_779), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n17134));
    defparam i1_2_lut_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i13531_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18111));
    defparam i13531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1300 (.I0(\data_in_frame[1][7] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[6] [4]), .I3(\data_in_frame[4] [2]), .O(n30496));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1301 (.I0(\data_in_frame[5] [4]), .I1(n30755), 
            .I2(\data_in_frame[5] [5]), .I3(\data_in_frame[7] [6]), .O(n30655));
    defparam i1_2_lut_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1302 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[6] [2]), .O(n6_adj_4072));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1]_c [3]), .I3(GND_net), .O(n6_adj_4065));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1304 (.I0(n17134), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_779), .I3(n30604), .O(n6_adj_4059));
    defparam i1_2_lut_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i13532_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18112));
    defparam i13532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1305 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(n10_adj_4058), .I3(\data_in_frame[4] [3]), .O(n8));   // verilog/coms.v(73[16:42])
    defparam i5_3_lut_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i13533_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18113));
    defparam i13533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13534_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18114));
    defparam i13534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1306 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(n30614), .O(n16954));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1307 (.I0(n63_adj_3958), .I1(n63_c), .I2(n63), 
            .I3(GND_net), .O(n13810));   // verilog/coms.v(157[6] 159[9])
    defparam i2_2_lut_3_lut_adj_1307.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(n16797), .I1(\data_in_frame[4] [6]), 
            .I2(n31067), .I3(GND_net), .O(n6_adj_4057));
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i13535_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18115));
    defparam i13535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n29947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n18347));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1309 (.I0(Kp_23__N_779), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1]_c [0]), .I3(\data_in_frame[3] [0]), .O(n17452));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n18346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n18345));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13536_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18116));
    defparam i13536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n18344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n18343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n18342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n18341));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13537_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18117));
    defparam i13537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13538_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30473), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18118));
    defparam i13538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13683_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n18263));
    defparam i13683_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13684_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n18264));
    defparam i13684_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13685_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n18265));
    defparam i13685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13686_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n18266));
    defparam i13686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13687_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n18267));
    defparam i13687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13688_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n18268));
    defparam i13688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1310 (.I0(n28697), .I1(\data_out_frame[23] [5]), 
            .I2(n16279), .I3(GND_net), .O(n30874));
    defparam i1_2_lut_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1311 (.I0(n30649), .I1(n30949), .I2(\data_out_frame[20] [7]), 
            .I3(n28699), .O(n31016));
    defparam i1_2_lut_4_lut_adj_1311.LUT_INIT = 16'h9669;
    SB_LUT4 i13689_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n18269));
    defparam i13689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_5_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n25556), .O(n2_adj_4159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n18055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n18340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n18339));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13473_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30455), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n18053));
    defparam i13473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_29325 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n35501));
    defparam byte_transmit_counter_0__bdd_4_lut_29325.LUT_INIT = 16'he4aa;
    SB_LUT4 equal_120_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4035));   // verilog/coms.v(154[7:23])
    defparam equal_120_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_130_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4179));   // verilog/coms.v(154[7:23])
    defparam equal_130_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13541_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18121));
    defparam i13541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n18338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n18337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n18336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n18335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n18334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n18333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n18332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n18331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n18330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n18329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n18328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n18327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n18326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n18325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n18324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n18323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n18317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n18316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n18315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n18314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n18313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n18312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n18311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n18310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n18309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n18308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n18307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n18306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n18305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n18304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n18303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n18302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n18301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n18300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode_c[0]), .C(clk32MHz), .D(n18054));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13542_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n18122));
    defparam i13542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n18053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n18052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n18051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n18050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n18049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n18299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n18298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n18297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n18296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n18295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n18294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n18293));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13543_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n18123));
    defparam i13543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n18040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n18292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n18291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n18290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n18289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n18288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n18287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n18286));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n18285));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n35501_bdd_4_lut (.I0(n35501), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n35504));
    defparam n35501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n18284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n18283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n18282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n18281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n18280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n18279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n18278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n18277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n18276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n18275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n18274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n18273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n18272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n18271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n18270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n18269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n18268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n18267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n18266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n18265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n18264));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13544_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n18124));
    defparam i13544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n18263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1]_c [0]), .C(clk32MHz), 
           .D(n18262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1]_c [1]), .C(clk32MHz), 
           .D(n18261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1]_c [2]), .C(clk32MHz), 
           .D(n18260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1]_c [3]), .C(clk32MHz), 
           .D(n18259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n18258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n18257));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1][6] ), .C(clk32MHz), 
           .D(n18256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1][7] ), .C(clk32MHz), 
           .D(n18255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n18254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n18253));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n18252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n18251));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n18250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n18249));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n18248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n18247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n18246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n18245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n18244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n18243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n18242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n18241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n18240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n18239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n18238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n18237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n18236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n18235));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n18234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n18233));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n18232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n18231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n18230));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n18229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n18228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n18227));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n18226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n18225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n18224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n18223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n18222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n18221));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13545_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n18125));
    defparam i13545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n18220));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n18219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n18218));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n18217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n18216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n18215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n18214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n18213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n18212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n18211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n18210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n18209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n18208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n18207));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13546_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n18126));
    defparam i13546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n18206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n18205));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1312 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [7]), .O(n29847));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1312.LUT_INIT = 16'hf400;
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18199));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1313 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [8]), .O(n29851));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1313.LUT_INIT = 16'hf400;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18187));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1314 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n32881));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_adj_1314.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n18179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18169));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1315 (.I0(n21861), .I1(n10_adj_4112), .I2(GND_net), 
            .I3(GND_net), .O(n30473));
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'hdddd;
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n18157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n18156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n18155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n18151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18144));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13539_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18119));
    defparam i13539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_5 (.CI(n25556), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n25557));
    SB_LUT4 i1_2_lut_4_lut_adj_1316 (.I0(n30649), .I1(n30949), .I2(\data_out_frame[20] [7]), 
            .I3(n16263), .O(n30863));
    defparam i1_2_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i13540_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30459), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18120));
    defparam i13540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18142));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18141));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1317 (.I0(n16882), .I1(n10_adj_4025), .I2(\data_in_frame[8] [2]), 
            .I3(\data_in_frame[8] [3]), .O(n28732));
    defparam i5_3_lut_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18140));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13675_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[7]), 
            .I3(\data_in_frame[1][7] ), .O(n18255));
    defparam i13675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18139));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18135));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13676_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[6]), 
            .I3(\data_in_frame[1][6] ), .O(n18256));
    defparam i13676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1318 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21861), .O(n30447));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1318.LUT_INIT = 16'hefff;
    SB_LUT4 i13677_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n18257));
    defparam i13677_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut (.I0(n16619), .I1(n13865), .I2(n13914), .I3(n16606), 
            .O(n4_adj_3951));   // verilog/coms.v(212[5:16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h44f4;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18130));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18129));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13678_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n18258));
    defparam i13678_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13679_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n18259));
    defparam i13679_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13680_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[2]), 
            .I3(\data_in_frame[1]_c [2]), .O(n18260));
    defparam i13680_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1319 (.I0(n27501), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[10] [2]), .I3(GND_net), .O(n30995));
    defparam i1_2_lut_3_lut_adj_1319.LUT_INIT = 16'h9696;
    SB_LUT4 i13681_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[1]), 
            .I3(\data_in_frame[1]_c [1]), .O(n18261));
    defparam i13681_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13682_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30447), .I2(rx_data[0]), 
            .I3(\data_in_frame[1]_c [0]), .O(n18262));
    defparam i13682_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n21861), .O(n30459));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_112_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3981));   // verilog/coms.v(154[7:23])
    defparam equal_112_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 add_43_2_lut (.I0(n2026), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18127));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29422 (.I0(byte_transmit_counter[1]), 
            .I1(n34086), .I2(n34087), .I3(byte_transmit_counter[2]), .O(n35495));
    defparam byte_transmit_counter_1__bdd_4_lut_29422.LUT_INIT = 16'he4aa;
    SB_LUT4 n35495_bdd_4_lut (.I0(n35495), .I1(n17_adj_4083), .I2(n16_adj_4080), 
            .I3(byte_transmit_counter[2]), .O(n35498));
    defparam n35495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13667_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n18247));
    defparam i13667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29316 (.I0(byte_transmit_counter[1]), 
            .I1(n34064), .I2(n34065), .I3(byte_transmit_counter[2]), .O(n35489));
    defparam byte_transmit_counter_1__bdd_4_lut_29316.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18126));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13668_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n18248));
    defparam i13668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13669_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n18249));
    defparam i13669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13670_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n18250));
    defparam i13670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18124));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13671_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n18251));
    defparam i13671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13672_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n18252));
    defparam i13672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13673_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n18253));
    defparam i13673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13674_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30459), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n18254));
    defparam i13674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n35489_bdd_4_lut (.I0(n35489), .I1(n17_adj_4063), .I2(n16_adj_4062), 
            .I3(byte_transmit_counter[2]), .O(n35492));
    defparam n35489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13659_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n18239));
    defparam i13659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1320 (.I0(\data_in_frame[1] [5]), .I1(n31055), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[6] [0]), .O(n30666));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i13660_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n18240));
    defparam i13660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18123));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13661_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n18241));
    defparam i13661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18121));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13662_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n18242));
    defparam i13662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(n16246), .I1(\data_out_frame[18] [0]), 
            .I2(\data_out_frame[18] [7]), .I3(GND_net), .O(n6_adj_3927));
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1322 (.I0(n16246), .I1(\data_out_frame[18] [0]), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n7));
    defparam i2_2_lut_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i13663_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n18243));
    defparam i13663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13664_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n18244));
    defparam i13664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13665_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n18245));
    defparam i13665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(tx_transmit_N_3304), .I1(n21830), 
            .I2(n13810), .I3(GND_net), .O(n13865));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'he0e0;
    SB_LUT4 i13666_3_lut_4_lut (.I0(n8_adj_3981), .I1(n30463), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n18246));
    defparam i13666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13651_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n18231));
    defparam i13651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(tx_transmit_N_3304), .I1(n21830), 
            .I2(n16619), .I3(GND_net), .O(n19));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'h0e0e;
    SB_LUT4 i13652_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n18232));
    defparam i13652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1325 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [9]), .O(n29855));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1325.LUT_INIT = 16'hf400;
    SB_LUT4 i13653_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n18233));
    defparam i13653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13654_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n18234));
    defparam i13654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13655_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n18235));
    defparam i13655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13656_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n18236));
    defparam i13656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29311 (.I0(byte_transmit_counter[1]), 
            .I1(n34068), .I2(n34069), .I3(byte_transmit_counter[2]), .O(n35483));
    defparam byte_transmit_counter_1__bdd_4_lut_29311.LUT_INIT = 16'he4aa;
    SB_LUT4 i13657_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n18237));
    defparam i13657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13658_3_lut_4_lut (.I0(n10_adj_4179), .I1(n30451), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n18238));
    defparam i13658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1326 (.I0(n21861), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n30451));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1326.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_4_lut_adj_1327 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n16954), .I3(n16963), .O(n27501));
    defparam i2_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1328 (.I0(\data_in_frame[14] [5]), .I1(n4_c), 
            .I2(n5_c), .I3(GND_net), .O(n10_adj_4023));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_3_lut_adj_1328.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1329 (.I0(n21861), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n30455));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1329.LUT_INIT = 16'hfffd;
    SB_LUT4 i13635_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n18215));
    defparam i13635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13636_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n18216));
    defparam i13636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13637_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n18217));
    defparam i13637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13638_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n18218));
    defparam i13638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13639_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n18219));
    defparam i13639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13640_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n18220));
    defparam i13640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13641_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n18221));
    defparam i13641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n35483_bdd_4_lut (.I0(n35483), .I1(n17_adj_4056), .I2(n16_adj_4055), 
            .I3(byte_transmit_counter[2]), .O(n35486));
    defparam n35483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13642_3_lut_4_lut (.I0(n8_adj_4068), .I1(n30463), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n18222));
    defparam i13642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1330 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [10]), .O(n29859));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1330.LUT_INIT = 16'hf400;
    SB_LUT4 i13627_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n18207));
    defparam i13627_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13628_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n18208));
    defparam i13628_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13629_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n18209));
    defparam i13629_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17421_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n21993));
    defparam i17421_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13630_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n18210));
    defparam i13630_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13631_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n18211));
    defparam i13631_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13632_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n18212));
    defparam i13632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13633_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n18213));
    defparam i13633_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13634_3_lut_4_lut (.I0(n21993), .I1(n30463), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n18214));
    defparam i13634_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[9] [6]), .I3(GND_net), .O(n30671));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 equal_117_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4068));
    defparam equal_117_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13619_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18199));
    defparam i13619_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1332 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [11]), .O(n29863));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1332.LUT_INIT = 16'hf400;
    SB_LUT4 i3_4_lut_adj_1333 (.I0(\data_out_frame[25] [6]), .I1(n28637), 
            .I2(n30870), .I3(n31034), .O(n32377));
    defparam i3_4_lut_adj_1333.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1334 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[25] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30870));
    defparam i1_2_lut_adj_1334.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1335 (.I0(\data_out_frame[18] [3]), .I1(n32847), 
            .I2(n30870), .I3(n30874), .O(n18_adj_4187));
    defparam i7_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1336 (.I0(n17262), .I1(n18_adj_4187), .I2(n28699), 
            .I3(n31078), .O(n20_adj_4188));
    defparam i9_4_lut_adj_1336.LUT_INIT = 16'h9669;
    SB_LUT4 i4_2_lut (.I0(n30949), .I1(n28404), .I2(GND_net), .I3(GND_net), 
            .O(n15_adj_4189));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1337 (.I0(n15_adj_4189), .I1(n20_adj_4188), .I2(n16671), 
            .I3(n31901), .O(n31747));
    defparam i10_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1338 (.I0(\data_out_frame[24] [1]), .I1(n28610), 
            .I2(n28379), .I3(n30778), .O(n32037));
    defparam i3_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1339 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [12]), .O(n29867));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1339.LUT_INIT = 16'hf400;
    SB_LUT4 i6_4_lut_adj_1340 (.I0(n31084), .I1(n27790), .I2(n30739), 
            .I3(\data_out_frame[23] [7]), .O(n14_adj_4190));
    defparam i6_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1341 (.I0(\data_out_frame[24] [2]), .I1(n14_adj_4190), 
            .I2(n10_adj_4180), .I3(n28725), .O(n31772));
    defparam i7_4_lut_adj_1341.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1342 (.I0(\data_out_frame[17] [4]), .I1(n31102), 
            .I2(n31022), .I3(n30806), .O(n28610));
    defparam i3_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1343 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [1]), .I3(\data_in_frame[9] [4]), .O(n30857));
    defparam i1_2_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1344 (.I0(\data_out_frame[24] [4]), .I1(n32847), 
            .I2(n27760), .I3(\data_out_frame[24] [3]), .O(n32412));
    defparam i3_4_lut_adj_1344.LUT_INIT = 16'h9669;
    SB_LUT4 i13620_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18200));
    defparam i13620_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_out_frame[19] [6]), .I1(n28723), 
            .I2(GND_net), .I3(GND_net), .O(n31022));
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1346 (.I0(n17226), .I1(n30969), .I2(n31022), 
            .I3(n31025), .O(n32564));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1347 (.I0(n2196), .I1(n30643), .I2(n32564), .I3(GND_net), 
            .O(n32219));
    defparam i2_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 i13621_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18201));
    defparam i13621_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[20] [1]), .I1(n31108), 
            .I2(GND_net), .I3(GND_net), .O(n30969));
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1349 (.I0(\data_in_frame[10] [3]), .I1(n17356), 
            .I2(n31132), .I3(GND_net), .O(n10_adj_4013));
    defparam i2_2_lut_3_lut_adj_1349.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1350 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_986), .I3(\data_in_frame[12] [6]), .O(n30620));
    defparam i2_3_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1351 (.I0(n32847), .I1(n28748), .I2(n30828), 
            .I3(n6_adj_4184), .O(n31697));
    defparam i4_4_lut_adj_1351.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29306 (.I0(byte_transmit_counter[1]), 
            .I1(n34071), .I2(n34072), .I3(byte_transmit_counter[2]), .O(n35477));
    defparam byte_transmit_counter_1__bdd_4_lut_29306.LUT_INIT = 16'he4aa;
    SB_LUT4 i13622_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18202));
    defparam i13622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13623_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18203));
    defparam i13623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1921_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_3963));
    defparam i1921_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i13624_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18204));
    defparam i13624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13625_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n18205));
    defparam i13625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_in_frame[9] [4]), .I1(n28088), 
            .I2(n17350), .I3(GND_net), .O(n28787));
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i13626_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30455), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n18206));
    defparam i13626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[11] [2]), 
            .I2(n30592), .I3(GND_net), .O(n31087));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_LUT4 n35477_bdd_4_lut (.I0(n35477), .I1(n17_adj_4053), .I2(n16_adj_4050), 
            .I3(byte_transmit_counter[2]), .O(n35480));
    defparam n35477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13611_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n18191));
    defparam i13611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1354 (.I0(n16246), .I1(n31052), .I2(n31712), 
            .I3(n28404), .O(n10_adj_4191));
    defparam i4_4_lut_adj_1354.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_out_frame[17] [5]), .I1(n28725), 
            .I2(GND_net), .I3(GND_net), .O(n31102));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i13612_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n18192));
    defparam i13612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1356 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [13]), .O(n29871));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1356.LUT_INIT = 16'hf400;
    SB_LUT4 i2_3_lut_4_lut_adj_1357 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(n8), .I3(Kp_23__N_986), .O(n30592));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1358 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [14]), .O(n29875));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1358.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [2]), 
            .I2(n28404), .I3(GND_net), .O(n28667));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1360 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [15]), .O(n29879));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1360.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(n28125), .I1(n30767), .I2(\data_in_frame[9] [6]), 
            .I3(GND_net), .O(n27688));
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_in_frame[10] [4]), .I1(n16954), 
            .I2(n30767), .I3(GND_net), .O(n31070));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1363 (.I0(\data_out_frame[24] [1]), .I1(n27760), 
            .I2(GND_net), .I3(GND_net), .O(n31084));
    defparam i1_2_lut_adj_1363.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(n28787), .I3(\data_in_frame[13] [6]), .O(n30809));
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1365 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30643));
    defparam i1_2_lut_adj_1365.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(\data_in_frame[10] [7]), .I1(n30787), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n31123));
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(Kp_23__N_1082), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[11] [6]), .I3(\data_in_frame[9] [5]), .O(n31117));
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1368 (.I0(n16895), .I1(\data_in_frame[9] [1]), 
            .I2(n8), .I3(n31129), .O(n30946));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut_adj_1369 (.I0(\data_in_frame[16] [2]), .I1(n17350), 
            .I2(n16895), .I3(n30638), .O(n11_adj_3985));   // verilog/coms.v(70[16:27])
    defparam i3_2_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(\data_in_frame[16] [2]), .I1(n17350), 
            .I2(n16895), .I3(GND_net), .O(n31075));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[24] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n30778));
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1372 (.I0(n16822), .I1(n30802), .I2(n8_adj_4185), 
            .I3(n30966), .O(n31078));
    defparam i1_4_lut_adj_1372.LUT_INIT = 16'h9669;
    SB_LUT4 i4_2_lut_4_lut_adj_1373 (.I0(\data_in[3] [4]), .I1(n10_adj_3972), 
            .I2(\data_in[2] [7]), .I3(\data_in[3] [0]), .O(n15_adj_3977));
    defparam i4_2_lut_4_lut_adj_1373.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_3_lut_4_lut_adj_1374 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n16594), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_3965));
    defparam i1_3_lut_4_lut_adj_1374.LUT_INIT = 16'hfefc;
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n16429), .O(n16607));   // verilog/coms.v(263[5:27])
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'hfffb;
    SB_LUT4 i28787_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n17937));
    defparam i28787_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut_adj_1376 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n1), .I3(\FRAME_MATCHER.state [1]), .O(n5_adj_3956));
    defparam i1_4_lut_4_lut_adj_1376.LUT_INIT = 16'h6273;
    SB_LUT4 i2_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state_31__N_2515 [3]), 
            .O(n6_adj_3957));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h8898;
    SB_LUT4 i2_3_lut_adj_1377 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(n28784), .I3(GND_net), .O(n30806));
    defparam i2_3_lut_adj_1377.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1378 (.I0(n31148), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n22632), .I3(n16614), .O(n16583));
    defparam i1_3_lut_4_lut_adj_1378.LUT_INIT = 16'haaae;
    SB_LUT4 i4_4_lut_adj_1379 (.I0(n30806), .I1(n28740), .I2(\data_out_frame[19] [2]), 
            .I3(n30823), .O(n10_adj_4178));
    defparam i4_4_lut_adj_1379.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1380 (.I0(n28725), .I1(n10_adj_4178), .I2(n28654), 
            .I3(GND_net), .O(n28379));
    defparam i5_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1381 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [16]), .O(n29883));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1381.LUT_INIT = 16'hf400;
    SB_LUT4 i2_3_lut_adj_1382 (.I0(n27790), .I1(n28740), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n17226));
    defparam i2_3_lut_adj_1382.LUT_INIT = 16'h6969;
    SB_LUT4 i13613_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n18193));
    defparam i13613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13614_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n18194));
    defparam i13614_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13615_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n18195));
    defparam i13615_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1383 (.I0(n30486), .I1(n31078), .I2(n28697), 
            .I3(n30778), .O(n30_adj_4192));
    defparam i11_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1384 (.I0(n28667), .I1(n30_adj_4192), .I2(n31016), 
            .I3(\data_out_frame[20] [3]), .O(n34_adj_4193));
    defparam i15_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i13616_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n18196));
    defparam i13616_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1385 (.I0(n17226), .I1(n30703), .I2(n31034), 
            .I3(n28748), .O(n32_adj_4194));
    defparam i13_4_lut_adj_1385.LUT_INIT = 16'h9669;
    SB_LUT4 i14_4_lut_adj_1386 (.I0(n31108), .I1(n28784), .I2(n30729), 
            .I3(n28622), .O(n33_adj_4195));
    defparam i14_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1387 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [1]), 
            .I2(n30617), .I3(n30843), .O(n6));
    defparam i1_2_lut_3_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29301 (.I0(byte_transmit_counter[1]), 
            .I1(n34074), .I2(n34075), .I3(byte_transmit_counter[2]), .O(n35471));
    defparam byte_transmit_counter_1__bdd_4_lut_29301.LUT_INIT = 16'he4aa;
    SB_LUT4 i13617_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n18197));
    defparam i13617_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13618_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30447), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n18198));
    defparam i13618_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1388 (.I0(\data_out_frame[23] [7]), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[23] [0]), .I3(n17457), .O(n31_adj_4196));
    defparam i12_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1389 (.I0(n2696), .I1(n13810), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state[3] ), .O(n29835));
    defparam i1_3_lut_4_lut_adj_1389.LUT_INIT = 16'hf800;
    SB_LUT4 i18_4_lut_adj_1390 (.I0(n31_adj_4196), .I1(n33_adj_4195), .I2(n32_adj_4194), 
            .I3(n34_adj_4193), .O(n31901));
    defparam i18_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i13603_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n18183));
    defparam i13603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1391 (.I0(n2696), .I1(n13810), .I2(n11_adj_3982), 
            .I3(n16604), .O(n9_adj_3953));
    defparam i1_3_lut_4_lut_adj_1391.LUT_INIT = 16'h88f8;
    SB_LUT4 i13604_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n18184));
    defparam i13604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1392 (.I0(n2483), .I1(n17440), .I2(n28631), .I3(n27784), 
            .O(n30860));
    defparam i3_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i13605_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n18185));
    defparam i13605_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13606_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n18186));
    defparam i13606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1393 (.I0(n30521), .I1(\data_out_frame[25] [7]), 
            .I2(n31901), .I3(n30541), .O(n10_adj_4183));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1393.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1394 (.I0(\FRAME_MATCHER.state [1]), .I1(n16429), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n16613));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_4_lut_adj_1394.LUT_INIT = 16'hfeff;
    SB_LUT4 i13607_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n18187));
    defparam i13607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16822));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1396 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [17]), .O(n29887));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1396.LUT_INIT = 16'hf400;
    SB_LUT4 i6_4_lut_adj_1397 (.I0(n30998), .I1(n31001), .I2(n28723), 
            .I3(n30992), .O(n15_adj_4197));
    defparam i6_4_lut_adj_1397.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1398 (.I0(n15_adj_4197), .I1(\data_out_frame[18] [0]), 
            .I2(n14_adj_4177), .I3(\data_out_frame[18] [1]), .O(n28622));
    defparam i8_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i13608_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n18188));
    defparam i13608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1399 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [18]), .O(n29891));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1399.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_adj_1400 (.I0(n2196), .I1(\data_out_frame[25] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n31061));
    defparam i1_2_lut_adj_1400.LUT_INIT = 16'h6666;
    SB_LUT4 i13609_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n18189));
    defparam i13609_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [31]), .O(n29939));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'hf400;
    SB_LUT4 i5_3_lut_4_lut_adj_1402 (.I0(n16246), .I1(\data_out_frame[18] [0]), 
            .I2(n27774), .I3(n10_adj_4191), .O(n31108));
    defparam i5_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i13610_3_lut_4_lut (.I0(n10_adj_4035), .I1(n30459), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n18190));
    defparam i13610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n35471_bdd_4_lut (.I0(n35471), .I1(n17_adj_4049), .I2(n16_adj_4048), 
            .I3(byte_transmit_counter[2]), .O(n35474));
    defparam n35471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1403 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [19]), .O(n29895));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1403.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(n16263), .I1(n27823), .I2(GND_net), 
            .I3(GND_net), .O(n30729));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1405 (.I0(n30714), .I1(\data_out_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n31001));
    defparam i1_2_lut_adj_1405.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1406 (.I0(n30770), .I1(n30737), .I2(\data_out_frame[17] [7]), 
            .I3(n31001), .O(n10_adj_4198));
    defparam i4_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1407 (.I0(n30758), .I1(n10_adj_4198), .I2(n28767), 
            .I3(GND_net), .O(n28404));
    defparam i5_3_lut_adj_1407.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1408 (.I0(\data_out_frame[23] [4]), .I1(n28697), 
            .I2(\data_out_frame[23] [5]), .I3(n16279), .O(n28631));
    defparam i1_2_lut_4_lut_adj_1408.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1409 (.I0(\data_out_frame[23] [3]), .I1(n28748), 
            .I2(\data_out_frame[23] [4]), .I3(GND_net), .O(n30966));
    defparam i1_2_lut_3_lut_adj_1409.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(\data_out_frame[19] [1]), .I1(n30515), 
            .I2(\data_out_frame[16] [5]), .I3(n17053), .O(n30834));
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1411 (.I0(\data_out_frame[24] [7]), .I1(n28667), 
            .I2(n30820), .I3(n6_adj_4182), .O(n2483));
    defparam i4_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_out_frame[25] [1]), .I1(n2483), 
            .I2(GND_net), .I3(GND_net), .O(n30575));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[14] [2]), 
            .I2(n16888), .I3(n30717), .O(n12_adj_3943));
    defparam i5_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1414 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5][6] ), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n6_adj_3941));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5][7] ), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n1241));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1416 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [20]), .O(n29899));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1416.LUT_INIT = 16'hf400;
    SB_LUT4 i17266_2_lut_4_lut (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [21]), .O(n21837));   // verilog/coms.v(212[5:16])
    defparam i17266_2_lut_4_lut.LUT_INIT = 16'hf400;
    SB_LUT4 i4_4_lut_adj_1417 (.I0(\data_out_frame[25] [2]), .I1(n17262), 
            .I2(n28702), .I3(n6_adj_4176), .O(n32125));
    defparam i4_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1418 (.I0(n2066), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[23] [0]), .I3(GND_net), .O(n30820));
    defparam i2_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n30992));
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(n17336), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n30998));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1421 (.I0(\data_out_frame[16] [1]), .I1(n1835), 
            .I2(n17057), .I3(n17336), .O(n30758));
    defparam i2_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1422 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[5][7] ), .O(n30899));
    defparam i2_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1423 (.I0(\data_out_frame[18] [2]), .I1(n30998), 
            .I2(n30992), .I3(n27850), .O(n12_adj_4199));
    defparam i5_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1424 (.I0(n30770), .I1(n12_adj_4199), .I2(n30758), 
            .I3(n31093), .O(n28699));
    defparam i6_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1425 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[13] [2]), .I3(n30837), .O(n6_adj_3940));
    defparam i1_2_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1426 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n30541));
    defparam i1_2_lut_adj_1426.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1427 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [22]), .O(n29903));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1427.LUT_INIT = 16'hf400;
    SB_LUT4 i4_4_lut_adj_1428 (.I0(\data_out_frame[20] [4]), .I1(n28730), 
            .I2(n30820), .I3(n6_adj_4175), .O(n17440));
    defparam i4_4_lut_adj_1428.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1429 (.I0(n17440), .I1(n30541), .I2(GND_net), 
            .I3(GND_net), .O(n30542));
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1430 (.I0(\data_out_frame[12] [0]), .I1(n30502), 
            .I2(\data_out_frame[13] [6]), .I3(n27850), .O(n12_adj_4200));
    defparam i5_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1431 (.I0(n17057), .I1(n12_adj_4200), .I2(n30887), 
            .I3(\data_out_frame[15] [7]), .O(n31712));
    defparam i6_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\data_out_frame[18] [4]), .I1(n14898), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4181));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1433 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [23]), .O(n29907));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1433.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17457));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1435 (.I0(n16697), .I1(n31049), .I2(n30562), 
            .I3(\data_out_frame[16] [3]), .O(n14898));
    defparam i3_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1436 (.I0(n14900), .I1(n30524), .I2(n14898), 
            .I3(GND_net), .O(n2066));
    defparam i2_3_lut_adj_1436.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1437 (.I0(\data_out_frame[18] [3]), .I1(n31712), 
            .I2(GND_net), .I3(GND_net), .O(n28730));
    defparam i1_2_lut_adj_1437.LUT_INIT = 16'h9999;
    SB_LUT4 i25081_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n22632));
    defparam i25081_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1438 (.I0(n30863), .I1(\data_out_frame[25] [3]), 
            .I2(n28730), .I3(n2066), .O(n14_adj_4201));
    defparam i6_4_lut_adj_1438.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [24]), .O(n29911));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'hf400;
    SB_LUT4 i7_4_lut_adj_1440 (.I0(n9_adj_4174), .I1(n14_adj_4201), .I2(n30802), 
            .I3(n32095), .O(n31607));
    defparam i7_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1441 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(n30846), .I3(n30617), .O(n28310));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1441.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1442 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [25]), .O(n29915));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1442.LUT_INIT = 16'hf400;
    SB_LUT4 i2_3_lut_4_lut_adj_1443 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[8] [4]), .O(n30929));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[8] [2]), .O(n31111));
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5]_c [1]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[7] [1]), .O(n30890));
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1446 (.I0(\data_out_frame[23] [2]), .I1(n27823), 
            .I2(GND_net), .I3(GND_net), .O(n30527));
    defparam i1_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1447 (.I0(\data_out_frame[23] [3]), .I1(n30527), 
            .I2(n16263), .I3(n16279), .O(n32095));
    defparam i3_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_4_lut (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[5] [4]), .O(n29));
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1448 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[25] [4]), 
            .I2(n27784), .I3(GND_net), .O(n32617));
    defparam i2_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [26]), .O(n29919));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'hf400;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29296 (.I0(byte_transmit_counter[1]), 
            .I1(n34077), .I2(n34078), .I3(byte_transmit_counter[2]), .O(n35465));
    defparam byte_transmit_counter_1__bdd_4_lut_29296.LUT_INIT = 16'he4aa;
    SB_LUT4 n35465_bdd_4_lut (.I0(n35465), .I1(n17_adj_4045), .I2(n16_adj_4042), 
            .I3(byte_transmit_counter[2]), .O(n35468));
    defparam n35465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n22));
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29291 (.I0(byte_transmit_counter[1]), 
            .I1(n34080), .I2(n34081), .I3(byte_transmit_counter[2]), .O(n35459));
    defparam byte_transmit_counter_1__bdd_4_lut_29291.LUT_INIT = 16'he4aa;
    SB_LUT4 n35459_bdd_4_lut (.I0(n35459), .I1(n17_adj_4041), .I2(n16_adj_4040), 
            .I3(byte_transmit_counter[2]), .O(n35462));
    defparam n35459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[14] [2]), 
            .I2(\data_out_frame[16] [7]), .I3(n28656), .O(n31004));
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_29286 (.I0(byte_transmit_counter[1]), 
            .I1(n34083), .I2(n34084), .I3(byte_transmit_counter[2]), .O(n35453));
    defparam byte_transmit_counter_1__bdd_4_lut_29286.LUT_INIT = 16'he4aa;
    SB_LUT4 n35453_bdd_4_lut (.I0(n35453), .I1(n17_adj_4039), .I2(n16_adj_4038), 
            .I3(byte_transmit_counter[2]), .O(n35456));
    defparam n35453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_56_i1_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[0] ), .I3(\encoder0_position_scaled[0] ), 
            .O(motor_state[0]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [27]), .O(n29923));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'hf400;
    SB_LUT4 i1_2_lut_4_lut_adj_1453 (.I0(n16619), .I1(n13865), .I2(n2_adj_3955), 
            .I3(\FRAME_MATCHER.state [28]), .O(n29927));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_4_lut_adj_1453.LUT_INIT = 16'hf400;
    SB_LUT4 mux_56_i2_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[1] ), .I3(\encoder0_position_scaled[1] ), 
            .O(motor_state[1]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i3_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[2] ), .I3(\encoder0_position_scaled[2] ), 
            .O(motor_state[2]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i4_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[3] ), .I3(\encoder0_position_scaled[3] ), 
            .O(motor_state[3]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i5_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[4] ), .I3(\encoder0_position_scaled[4] ), 
            .O(motor_state[4]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i6_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[5] ), .I3(\encoder0_position_scaled[5] ), 
            .O(motor_state[5]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i7_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[6] ), .I3(\encoder0_position_scaled[6] ), 
            .O(motor_state[6]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i8_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[7] ), .I3(\encoder0_position_scaled[7] ), 
            .O(motor_state[7]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i9_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[8] ), .I3(\encoder0_position_scaled[8] ), 
            .O(motor_state[8]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i10_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[9] ), .I3(\encoder0_position_scaled[9] ), 
            .O(motor_state[9]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i11_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[10] ), .I3(\encoder0_position_scaled[10] ), 
            .O(motor_state[10]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[14] [2]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n30783));
    defparam i1_2_lut_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 mux_56_i12_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[11] ), .I3(\encoder0_position_scaled[11] ), 
            .O(motor_state[11]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i13_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[12] ), .I3(\encoder0_position_scaled[12] ), 
            .O(motor_state[12]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i14_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[13] ), .I3(\encoder0_position_scaled[13] ), 
            .O(motor_state[13]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i15_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[14] ), .I3(\encoder0_position_scaled[14] ), 
            .O(motor_state[14]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i16_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[15] ), .I3(\encoder0_position_scaled[15] ), 
            .O(motor_state[15]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i17_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[16] ), .I3(\encoder0_position_scaled[16] ), 
            .O(motor_state[16]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i18_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[17] ), .I3(\encoder0_position_scaled[17] ), 
            .O(motor_state[17]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(n30863), .I1(n30966), .I2(n32095), 
            .I3(GND_net), .O(n27784));
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'h6969;
    SB_LUT4 mux_56_i19_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[18] ), .I3(\encoder0_position_scaled[18] ), 
            .O(motor_state[18]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i20_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[19] ), .I3(\encoder0_position_scaled[19] ), 
            .O(motor_state[19]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i2_3_lut_4_lut_adj_1456 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[10] [0]), .O(n30884));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 mux_56_i21_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[20] ), .I3(\encoder0_position_scaled[20] ), 
            .O(motor_state[20]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i2_3_lut_4_lut_adj_1457 (.I0(n30863), .I1(n30966), .I2(n28631), 
            .I3(n30521), .O(n32090));
    defparam i2_3_lut_4_lut_adj_1457.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[9] [3]), .O(n30711));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 mux_56_i22_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[21] ), .I3(\encoder0_position_scaled[22] ), 
            .O(motor_state[21]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i24_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[23] ), .I3(\encoder0_position_scaled[22] ), 
            .O(motor_state[23]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_56_i23_3_lut_4_lut (.I0(control_mode_c[1]), .I1(n21710), 
            .I2(\motor_state_23__N_74[22] ), .I3(\encoder0_position_scaled[22] ), 
            .O(motor_state[22]));   // verilog/coms.v(127[12] 300[6])
    defparam mux_56_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i5_3_lut_4_lut_adj_1459 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [4]), .I3(n10_adj_3936), .O(n16666));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[5]_c [0]), .I3(GND_net), .O(n4_adj_3938));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(n16878), .I1(\data_out_frame[14] [3]), 
            .I2(n32935), .I3(n17040), .O(n17053));
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1462 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [3]), 
            .I2(n30823), .I3(n28784), .O(n28697));
    defparam i2_3_lut_4_lut_adj_1462.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1463 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n30623));
    defparam i2_2_lut_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1464 (.I0(\data_out_frame[12] [1]), .I1(n30499), 
            .I2(n30884), .I3(\data_out_frame[5] [5]), .O(n30905));
    defparam i1_2_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1465 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[5] [2]), .O(n6_adj_3929));   // verilog/coms.v(71[16:27])
    defparam i1_3_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 i17146_3_lut (.I0(\data_out_frame[5]_c [1]), .I1(control_mode_c[1]), 
            .I2(n13933), .I3(GND_net), .O(n18448));
    defparam i17146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26960_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33129));
    defparam i26960_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1466 (.I0(\FRAME_MATCHER.state [1]), .I1(n30361), 
            .I2(n33129), .I3(\FRAME_MATCHER.state[0] ), .O(n13703));
    defparam i1_4_lut_adj_1466.LUT_INIT = 16'hccce;
    SB_LUT4 i3_4_lut_adj_1467 (.I0(n13703), .I1(n16614), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state_31__N_2515 [3]), .O(n13933));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1467.LUT_INIT = 16'h2000;
    SB_LUT4 i17147_3_lut (.I0(\data_out_frame[5]_c [0]), .I1(control_mode_c[0]), 
            .I2(n13933), .I3(GND_net), .O(n18449));
    defparam i17147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1468 (.I0(n17053), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [4]), .I3(n16702), .O(n14900));
    defparam i2_3_lut_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1469 (.I0(n27850), .I1(\data_out_frame[13] [4]), 
            .I2(n16666), .I3(n30714), .O(n30737));
    defparam i1_2_lut_4_lut_adj_1469.LUT_INIT = 16'h9669;
    SB_LUT4 i13523_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18103));
    defparam i13523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13524_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18104));
    defparam i13524_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13525_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18105));
    defparam i13525_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n30598));
    defparam i2_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i13526_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18106));
    defparam i13526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13527_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18107));
    defparam i13527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i17787_2_lut_4_lut (.I0(n31_adj_4007), .I1(n31_adj_3932), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n14151), .O(n1));
    defparam i17787_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 i3_2_lut_4_lut_adj_1471 (.I0(n31_adj_4007), .I1(n31_adj_3932), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[3] ), 
            .O(n11));
    defparam i3_2_lut_4_lut_adj_1471.LUT_INIT = 16'hffca;
    SB_LUT4 i13528_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18108));
    defparam i13528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13529_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18109));
    defparam i13529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13530_3_lut_4_lut (.I0(n10_adj_4112), .I1(n30451), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18110));
    defparam i13530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1472 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n30463), .I3(\FRAME_MATCHER.i [0]), .O(n30466));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1472.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_4_lut_adj_1473 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[12] [3]), .I3(n10_adj_3931), .O(n30515));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    uart_tx tx (.GND_net(GND_net), .VCC_net(VCC_net), .n17831(n17831), 
            .clk32MHz(clk32MHz), .n17982(n17982), .r_SM_Main({r_SM_Main}), 
            .\r_SM_Main_2__N_3404[1] (\r_SM_Main_2__N_3404[1] ), .tx_o(tx_o), 
            .tx_data({tx_data}), .\r_SM_Main_2__N_3407[0] (r_SM_Main_2__N_3407[0]), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n4(n4), .n18322(n18322), 
            .n18058(n18058), .tx_active(tx_active), .n35944(n35944), .n9799(n9799), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.GND_net(GND_net), .n17825(n17825), .clk32MHz(clk32MHz), 
            .n17980(n17980), .VCC_net(VCC_net), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_5 ), 
            .n16549(n16549), .n4(n4_adj_6), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), 
            .n18488(n18488), .rx_data_ready(rx_data_ready), .n21943(n21943), 
            .n4_adj_1(n4_adj_7), .n4_adj_2(n4_adj_8), .n16544(n16544), 
            .n18540(n18540), .rx_data({rx_data}), .n18048(n18048), .n18047(n18047), 
            .n18046(n18046), .n18045(n18045), .n18044(n18044), .n18043(n18043), 
            .n18042(n18042)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (GND_net, VCC_net, n17831, clk32MHz, n17982, r_SM_Main, 
            \r_SM_Main_2__N_3404[1] , tx_o, tx_data, \r_SM_Main_2__N_3407[0] , 
            \r_Bit_Index[0] , n4, n18322, n18058, tx_active, n35944, 
            n9799, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    output n17831;
    input clk32MHz;
    output n17982;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3404[1] ;
    output tx_o;
    input [7:0]tx_data;
    input \r_SM_Main_2__N_3407[0] ;
    output \r_Bit_Index[0] ;
    output n4;
    input n18322;
    input n18058;
    output tx_active;
    input n35944;
    output n9799;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n26322, n26321, n26320, n26319, n26318, n26317, n26316, 
        n26315;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n17963, n3, n1, n13923;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n11632, n22679, n11631, n35636, n35528, o_Tx_Serial_N_3435, 
        n10, n32075, n35633, n35525, n3_adj_3924;
    
    SB_LUT4 r_Clock_Count_1466_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n26322), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1466_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n26321), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_9 (.CI(n26321), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n26322));
    SB_LUT4 r_Clock_Count_1466_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n26320), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_8 (.CI(n26320), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n26321));
    SB_LUT4 r_Clock_Count_1466_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n26319), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_7 (.CI(n26319), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n26320));
    SB_LUT4 r_Clock_Count_1466_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n26318), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_6 (.CI(n26318), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n26319));
    SB_LUT4 r_Clock_Count_1466_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n26317), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_5 (.CI(n26317), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n26318));
    SB_LUT4 r_Clock_Count_1466_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n26316), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_4 (.CI(n26316), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n26317));
    SB_LUT4 r_Clock_Count_1466_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n26315), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_3 (.CI(n26315), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n26316));
    SB_LUT4 r_Clock_Count_1466_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1466_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1466_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n26315));
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n17831), 
            .D(n307[2]), .R(n17982));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n17831), 
            .D(n307[1]), .R(n17982));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i28809_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3404[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n17963));
    defparam i28809_4_lut.LUT_INIT = 16'h4445;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n11632), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i7130_4_lut (.I0(\r_SM_Main_2__N_3407[0] ), .I1(n22679), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3404[1] ), .O(n11631));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7130_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7131_3_lut (.I0(n11631), .I1(\r_SM_Main_2__N_3404[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n11632));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7131_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR r_Clock_Count_1466__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1858964_i1_3_lut (.I0(n35636), .I1(n35528), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3435));
    defparam i1858964_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3435), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_1466__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1569_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1569_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n32075));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n32075), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3404[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n22679));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13402_3_lut (.I0(n17831), .I1(n22679), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17982));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13402_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1576_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1576_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n35633));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n35633_bdd_4_lut (.I0(n35633), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n35636));
    defparam n35633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_29427 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n35525));
    defparam r_Bit_Index_0__bdd_4_lut_29427.LUT_INIT = 16'he4aa;
    SB_LUT4 n35525_bdd_4_lut (.I0(n35525), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n35528));
    defparam n35525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_1466__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1466__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1466__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1466__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1466__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1466__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13923), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3924), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1466__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n17963));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3404[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i9171_2_lut_3_lut (.I0(\r_SM_Main_2__N_3404[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3924));
    defparam i9171_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n18322));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n18058));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n35944));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3407[0] ), 
            .I3(r_SM_Main[1]), .O(n13923));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3404[1] ), .O(n17831));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i5306_2_lut (.I0(\r_SM_Main_2__N_3407[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n9799));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5306_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, n17825, clk32MHz, n17980, VCC_net, \r_Bit_Index[0] , 
            n16549, n4, r_Rx_Data, RX_N_2, n18488, rx_data_ready, 
            n21943, n4_adj_1, n4_adj_2, n16544, n18540, rx_data, 
            n18048, n18047, n18046, n18045, n18044, n18043, n18042) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n17825;
    input clk32MHz;
    output n17980;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n16549;
    output n4;
    output r_Rx_Data;
    input RX_N_2;
    input n18488;
    output rx_data_ready;
    output n21943;
    output n4_adj_1;
    output n4_adj_2;
    output n16544;
    input n18540;
    output [7:0]rx_data;
    input n18048;
    input n18047;
    input n18046;
    input n18045;
    input n18044;
    input n18043;
    input n18042;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n26314, n26313, n26312, n26311, n26310, n26309, n26308;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_2__N_3333;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n30433, n16447;
    wire [2:0]r_SM_Main_2__N_3339;
    
    wire n31284, n31286, n17961, n6, n17815, n22821, n3, r_Rx_Data_R, 
        n12, n8, n22665, n22751, n1, n10, n30081, n17758;
    
    SB_LUT4 r_Clock_Count_1464_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n26314), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1464_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n26313), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1464_add_4_8 (.CI(n26313), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n26314));
    SB_LUT4 r_Clock_Count_1464_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n26312), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1464_add_4_7 (.CI(n26312), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n26313));
    SB_LUT4 r_Clock_Count_1464_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n26311), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1464_add_4_6 (.CI(n26311), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n26312));
    SB_LUT4 r_Clock_Count_1464_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n26310), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1464_add_4_5 (.CI(n26310), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n26311));
    SB_LUT4 r_Clock_Count_1464_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n26309), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1464_add_4_4 (.CI(n26309), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n26310));
    SB_LUT4 r_Clock_Count_1464_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n26308), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n17825), 
            .D(n326[2]), .R(n17980));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n17825), 
            .D(n326[1]), .R(n17980));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY r_Clock_Count_1464_add_4_3 (.CI(n26308), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n26309));
    SB_LUT4 r_Clock_Count_1464_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1464_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3333[2]), 
            .R(n30433));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_3333[2]), .O(n16447));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(\r_Bit_Index[0] ), .I1(n16447), .I2(GND_net), 
            .I3(GND_net), .O(n16549));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_138_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_138_i4_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY r_Clock_Count_1464_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n26308));
    SB_LUT4 i25125_2_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3339[0]), .I2(GND_net), 
            .I3(GND_net), .O(n31284));
    defparam i25125_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n31286), .I2(r_SM_Main_2__N_3333[2]), 
            .I3(r_SM_Main[1]), .O(n17961));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main_2__N_3339[0]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i28769_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6), 
            .I3(r_Rx_Data), .O(n17815));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i28769_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3333[2]), 
            .I2(r_SM_Main[1]), .I3(n31284), .O(n22821));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h707a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_2));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1464__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n17815), .D(n37[0]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i5_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[0]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i6_4_lut (.I0(r_Clock_Count[2]), .I1(n12), .I2(r_Clock_Count[4]), 
            .I3(n8), .O(r_SM_Main_2__N_3339[0]));
    defparam i6_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n22665), .I1(r_SM_Main_2__N_3333[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n22751));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3339[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n22751), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1547_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1547_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_839 (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[7]), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(120[34:51])
    defparam i1_2_lut_adj_839.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[3]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i18103_4_lut (.I0(r_Clock_Count[5]), .I1(n8), .I2(n10), .I3(r_Clock_Count[1]), 
            .O(r_SM_Main_2__N_3333[2]));
    defparam i18103_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n22665));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13400_3_lut (.I0(n17825), .I1(n22665), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n17980));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13400_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3333[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n17825));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1554_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1554_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n22821), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1464__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n17815), .D(n37[7]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n18488));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n30081));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i17372_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n21943));
    defparam i17372_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_134_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_134_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_136_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_136_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_840 (.I0(n16447), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n16544));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_840.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18540));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1464__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n17815), .D(n37[6]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1464__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n17815), .D(n37[5]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1464__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n17815), .D(n37[4]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1464__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n17815), .D(n37[3]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1464__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n17815), .D(n37[2]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n18048));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n18047));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n18046));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n18045));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n18044));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n18043));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n18042));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Clock_Count_1464__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n17815), .D(n37[1]), .R(n17961));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i25127_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_Rx_Data), .I2(r_SM_Main_2__N_3339[0]), 
            .I3(GND_net), .O(n31286));
    defparam i25127_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3333[2]), 
            .I3(r_SM_Main[0]), .O(n17758));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n17758), 
            .I3(rx_data_ready), .O(n30081));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i28952_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n30433));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i28952_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    
endmodule
