// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Feb 17 14:44:31 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(116[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(117[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(126[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(223[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(225[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(226[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(227[22:30])
    
    wire n48687;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(228[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(229[22:24])
    
    wire n38453, n38682;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(231[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(232[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(233[22:35])
    
    wire n43821, n44589;
    wire [12:0]current;   // verilog/TinyFPGA_B.v(235[22:29])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(263[22:33])
    wire [7:0]data;   // verilog/TinyFPGA_B.v(326[14:18])
    
    wire data_ready, sda_out, n38681, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(350[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(358[15:20])
    
    wire pwm_setpoint_23__N_215;
    wire [23:0]pwm_setpoint_23__N_191;
    wire [23:0]pwm_setpoint_23__N_11;
    wire [7:0]commutation_state_7__N_216;
    
    wire commutation_state_7__N_224, n28235, n28234;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(222[11:28])
    
    wire n28233, n28232, n28231, n28230, n28229, n28228, GHA_N_367, 
        GLA_N_384, GHB_N_389, GLB_N_398, GHC_N_403, GLC_N_412, dti_N_416, 
        n28227, n28226, n28225, n28224, n28223, n28222, n28221, 
        RX_N_10, n1632;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_279;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        read_N_421, n731, n1195, n28220, n7, n38452, n1673;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(224[11:28])
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n38451, n28219, n48659, n26227, n38680, n38450;
    wire [3:0]state_3__N_528;
    
    wire n38679, n38678, n38677, n38676, n38675, n26367, n38449, 
        n5, n38198, n38674, n15, n48209, n38197, n38673, n38448, 
        n10, n38196, n38672, n28218, n4, n28217, n28216, n28215, 
        n28214, n38447, n38671, n28213, n6976, n28212, n28211, 
        n28210, n38446, n38670, n38669, n28209, n38668, n652, 
        n38445, n38667, \neo_pixel_transmitter.done_N_742 , n4_adj_5161, 
        n38666, n28208, n28207, n38444, n28206, n28205, n38665, 
        n28204, n38664, n28203, n38443, n38663, n38442, n38662, 
        n28202, n28200, n38661, n625;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n38660, n28199, n623, n3, n4_adj_5162, n5_adj_5163, n6, 
        n7_adj_5164, n8, n9, n10_adj_5165, n11, n12, n13, n14, 
        n15_adj_5166, n16, n17, n18, n19, n20, n21, n22, n23, 
        n24, n25, n622, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire n621, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n38659, n15_adj_5167, n38658, n14_adj_5168, n38657, n38922, 
        n122, n38921, n38656, n38920, n38655, n43900, n42022, 
        n25_adj_5169, n17_adj_5170, n38654, n38919, n38653, n38918, 
        n38917, n38916, n38915, n38652, n34453, n38651, n38914, 
        n38913, n38650, n38912, n38911, n38910, n38909, n38649, 
        n7_adj_5171, n38908, n26226, n38907, n38906, n38905, n38904, 
        n38903, n38902, n38901, n38900, n38899, n43911, n38648, 
        n38647, n38898, n38646, n38645, n38644, n38897, n34562, 
        n38896, n38643, n14_adj_5172, n38642, n38895, n38195, n38894, 
        n38641, n38640, n38639, n38638, n38637, n34566, n38636, 
        n38635, n38893, n38634, n38633, n38194, n38892, n38891, 
        n38890, n38889, n38888, n38887, n34688, n33899, n38632, 
        n38631, n38886, n38630, n38885, n34634, n33894, n38884, 
        n38883, n38882, n38881, n38425, n38880, n38424, n41744, 
        n38629, n38879, n38423, n34684, n38628, n38627, n38878, 
        n38877, n38876, n38875, n38626, n38625, n38624, n38623, 
        n49229, n38874, n38622, n34678, n38873, n38872, n38621, 
        n38620, n38871, n34676, n38870, n38619, n38869, n38422, 
        n38868, n38421, n38618, n38867, n38420, n34672, n36539, 
        n38866, n38865, n38864, n38617, n38616, n38863, n38862, 
        n48634, n38861, n34662, n38860, n38615, n38859, n34658, 
        n38858, n38857, n38614, n38613, n34654, n38193, n38612, 
        n38611, n38610, n34646, n34644, n38609, n38419, n34642, 
        n38192, n38608, n38418, n38607, n38606, n38856, n38417, 
        n38605, n38416, n38191, n38415, n38604, n38855, n38190, 
        n38854, n38189, n38603, n38602, n38414, n38853, n38601, 
        n38413, n38412, n38188, n38600, n38852, n38411, n38599, 
        n38598, n38597, n38596, n38851, n34616, n38850, n38410, 
        n38187, n38114, n38595, n38849, n38186, n38848, n38185, 
        n38847, n34610, n38409, n38594, n38593, n38408, n38592, 
        n38407, n38113, n34608, n38591, n38184, n38183, n38590, 
        n38846, n38589, n38182, n38406, n33869, n38845, n34602, 
        n44948, n38588, n38181, n38405, n38180, n38179, n38178, 
        n38844, n38177, n38404, n38587, n38403, n34598, n38843, 
        n34596, n38586, n38842, n38841, n38840, n34594, n38176, 
        n33855, n38839, n38112, n38585, n38838, n38837, n38111, 
        n38584, n38110, n2, n15_adj_5173, n38836, n12_adj_5174, 
        n38583, n38582, n38835, n3303, n38834, n43969, n38581, 
        n38580, n48746, n38833, n38579, n38578, n34588, n38832, 
        n7_adj_5175, n38098, n48719, n4452, n38577, n38576, n38831, 
        n38575, n122_adj_5176, n38830, n38829, n38574, n38828, n43926, 
        n43941, n4_adj_5177, n38827, n38573, n29908, n38572, n38571, 
        n38826, n38570, n38825, n38824, n38823, n2_adj_5178, n23755, 
        n5_adj_5179, n26211, n25_adj_5180, n24_adj_5181, n38569, n38568, 
        n38822, \FRAME_MATCHER.i_31__N_2622 , \FRAME_MATCHER.i_31__N_2624 , 
        n38567, \FRAME_MATCHER.i_31__N_2626 , n5_adj_5182, n45208, n48309, 
        n405, n23_adj_5183, n22_adj_5184, n21_adj_5185, n20_adj_5186, 
        n19_adj_5187, n18_adj_5188, n17_adj_5189, n16_adj_5190, n15_adj_5191, 
        n14_adj_5192, n13_adj_5193, n12_adj_5194, n11_adj_5195, n10_adj_5196, 
        n9_adj_5197, n8_adj_5198, n7_adj_5199, n6_adj_5200, n5_adj_5201, 
        n4_adj_5202, n3_adj_5203, n46038, n14_adj_5204, n46036, n5615, 
        n46032, n38821, n10_adj_5205, n43826, n46026, n38820, n38566, 
        n38565, n38819, n38818, n38564, n38563, n28715, n46020, 
        n38817, n38562, n38561, n38816, n38560, n38815, n38559, 
        n38814, n38558, n46014, n48601, n43846, n28714, n46008, 
        n28713, n28712, n28711, n28710, n28709, n46004, n46002, 
        n28708, n28707, n28706, n28705, n28704, n28703, n28702, 
        n28701, n28700, n28699, n28698, n28697, n38109, n38813, 
        n45990, n38557, n34584, n8_adj_5206, n49000, n28696, n28695, 
        n28694, n28693, n28692, n28691, n28690, n28689, n45984;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n28688, n28687, n28686, n28685, n28684, n28683, 
        n28682, n28681, n28680, direction_N_3907, n45978, n28662, 
        n28661, n5_adj_5207, n38812, n45972, n28198, n38556, n28638, 
        n28637, n38811, n45970, n28636, n28635, n28634, n28633, 
        n28632;
    wire [1:0]a_new_adj_5349;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5209, n38097, n1973, n1964, n38555, n28630, 
        n28629, n38554, n38553, n38552, n4_adj_5210, n45964, n45962, 
        direction_N_3907_adj_5211, n45960, n28623, n28622, n28621, 
        n28620, n28619, n28618, n28617, n28616, n28615, n28614, 
        n28613, n28612, n34578, n38551, n43883, n5_adj_5212, n28577, 
        rw;
    wire [7:0]state_adj_5373;   // verilog/eeprom.v(23[11:16])
    
    wire n45944, n28576, n28575, n28574, n28573, n28572, n28571, 
        n28570, n28569, n28568, n33, n28567, n45938, n28566, n28565;
    wire [15:0]data_adj_5377;   // verilog/tli4970.v(27[14:18])
    
    wire n45932, n38550, n34576, n28564, n28563, n28562, n28561, 
        n28560, n32, n31, n28559, n28558, n28197, n28196, n28195, 
        n28194, n28193, n28192, n28191, n28190, n28189, n28188, 
        n28187, n28186, n28185, n28184, n28183, n28182, n28557, 
        n48571, n28556, n28555, n45926, n4_adj_5222, n28554, n28553, 
        n28552, n38108, n38549, n27804, n28551, n28550, n28549, 
        n28548, n28547, n28545, n28544, n28542, n28541, n28540, 
        n28539, n28538, n28537, n28536, n45920, n38548, n38810, 
        n28534, n30, n45918, n28529, state_7__N_4293, n7072, n38809, 
        n38144, n28181, n28180, n38096, n28516, n28515, n28514, 
        n28513, n28512, n28511, n28510, n38547, n28509, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n38143, n4_adj_5223, n3813, n45916, n38808, n38546, n38545, 
        n38807, n38806, n38544, n27767, n28015, n34568, n27763;
    wire [2:0]r_SM_Main_2__N_3542;
    
    wire n28179;
    wire [2:0]r_SM_Main_adj_5388;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5390;   // verilog/uart_tx.v(33[16:27])
    
    wire n38142, n38543, n38542, n38541, n38805;
    wire [2:0]r_SM_Main_2__N_3613;
    
    wire n38804, n38141, n38540, n38803, n28452, n28451, n28450;
    wire [7:0]state_adj_5401;   // verilog/i2c_controller.v(33[12:17])
    
    wire n28449, n38802, n28448;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n28056, n28054, n28447, n28446, n6_adj_5229, n7233, n38539, 
        n9_adj_5230, n38538, n38537, n38801, n38107;
    wire [7:0]state_7__N_4087;
    
    wire n28445, n28178, n38536, n38800, n38799, n38535, n38798, 
        n38095, n11_adj_5231, n28438, n28437;
    wire [7:0]state_7__N_4103;
    
    wire n38534, n38533, n38532, n28433, n38531, n28432, n28431, 
        n28430, n28429, n28428, n28427, n28426, n38530, n38797, 
        n38796, n28425, n28424, n45896, n28423, n28177, n28176, 
        n28175, n28174, n28173, n28172, n28171, n28170, n29, n28169, 
        n28422, n28168, n28167, n28421, n38795, n4_adj_5232, n28420, 
        n28419, n28, n27, n26, n25_adj_5233, n24_adj_5234, n23_adj_5235, 
        n22_adj_5236, n21_adj_5237, n20_adj_5238, n19_adj_5239, n18_adj_5240, 
        n17_adj_5241, n16_adj_5242, n15_adj_5243, n14_adj_5244, n13_adj_5245, 
        n12_adj_5246, n11_adj_5247, n10_adj_5248, n9_adj_5249, n8_adj_5250, 
        n28417, n28166, n28165, n28164, n28163, n28162, n28161, 
        n28160, n28159, n28156, n28155, n28153, n28152, n28151, 
        n28149, n28148, n28146, n28145, n28144, n28143, n28142, 
        n28141, n28140, n28139, n28138, n28137, n28135, n28134, 
        n28133, n28132, n28131, n28130, n28129, n28416, n28415, 
        n38140, n28414, n38139, n38794, n28413, n38529, n28412, 
        n28411, n28410, n28409, n27713, n28128, n28127, n28408, 
        n28407, n3_adj_5251, n28406, n28405, n28404, n828, n829, 
        n830, n831, n832, n833, n834, n861, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n934, n935, n936, n937, n938, n939, n940, n941, 
        n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n960, n995, 
        n996, n997, n998, n999, n1000, n1001, n6_adj_5252, n1026, 
        n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1059, 
        n48540, n1093_adj_5253, n1094_adj_5254, n1095_adj_5255, n1096_adj_5256, 
        n1097_adj_5257, n1098_adj_5258, n1099_adj_5259, n1100_adj_5260, 
        n1101_adj_5261, n45890, n1125, n1126, n1127, n1128, n1129, 
        n1130, n1131, n1132, n1133, n1158, n45884, n1193, n1194, 
        n1195_adj_5262, n1196, n1197, n1198, n1199, n1200, n1201, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n42504, n42634, n28125, n28087, n1257, n38528, 
        n48291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
        n1299, n1300, n1301, n38793, n45878, n45876, n38792, n1323, 
        n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
        n1332, n1333, n38527, n45868, n1356, n45858, n1391, n1392, 
        n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
        n1401, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
        n1429, n1430, n1431, n1432, n1433, n48330, n1455, n45852, 
        n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
        n1497, n1498, n1499, n1500, n1501, n43868, n45846, n1521, 
        n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
        n1530, n1531, n1532, n1533, n1554, n1589, n1590, n1591, 
        n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
        n1600, n1601, n45840, n1620, n1621, n1622, n1623, n1624, 
        n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632_adj_5263, 
        n1633, n1653, n45838, n1688, n1689, n1690, n1691, n1692, 
        n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
        n1701, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
        n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
        n1752, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
        n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
        n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
        n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
        n45830, n1851, n1886, n1887, n1888, n1889, n1890, n1891, 
        n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
        n1900, n1901, n23568, n45820, n1917, n1918, n1919, n1920, 
        n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
        n1929, n1930, n1931, n1932, n1933, n1950, n45814, n45808, 
        n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
        n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
        n2001, n48507, n2016, n2017, n2018, n2019, n2020, n2021, 
        n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n45804, n2049, n28403, n38106, 
        n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, 
        n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
        n2100, n2101, n38791, n2115, n2116, n2117, n2118, n2119, 
        n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
        n2128, n2129, n2130, n2131, n2132, n2133, n2148, n38138, 
        n45796, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
        n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
        n2198, n2199, n2200, n2201, n2214, n2215, n2216, n2217, 
        n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
        n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
        n26390, n26385, n2247, n28402, n2282, n2283, n2284, n2285, 
        n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
        n45786, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
        n2320, n2321, n2322, n2323, n2327, n2329, n2330, n2331, 
        n2332, n2333, n2346, n5_adj_5264, n2381, n2382, n2383, 
        n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, 
        n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
        n2400, n2401, n2412, n2413, n2414, n2415, n2416, n2417, 
        n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, 
        n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
        n2445, n42843, n42836, n2480, n2481, n2482, n2483, n2484, 
        n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
        n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
        n2501, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
        n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
        n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
        n45780, n2544, n44891, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2643, n45774, n2678, n2679, n2680, n2681, 
        n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
        n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, 
        n2698, n2699, n2700, n2701, n45770, n2709, n2710, n2711, 
        n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
        n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
        n2728, n2729, n2730, n2731, n2732, n2733, n2742, n42422, 
        n28401, n42822, n2777, n2778, n2779, n2780, n2781, n2782, 
        n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
        n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
        n2799, n2800, n2801, n2808, n2809, n2810, n2811, n2812, 
        n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
        n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
        n2829, n2830, n2831, n2832, n2833, n2841, n45766, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
        n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
        n2930, n2931, n2932, n2933, n2940, n2975, n2976, n2977, 
        n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
        n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
        n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
        n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
        n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
        n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
        n3030, n3031, n3032, n3033, n3039, n26380, n26377, n3074, 
        n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
        n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
        n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
        n3099, n3100, n3101, n3105, n3106, n3107, n3108, n3109, 
        n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
        n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
        n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3138, n45760, n26372, n3173, n3174, n3175, n3176, n3177, 
        n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
        n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
        n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
        n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
        n3228, n3229, n3230, n3231, n3232, n3233, n3237, n28124, 
        n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
        n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
        n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
        n3295, n3296, n3298, n3299, n3300, n3301, n45750, n48475, 
        n45746, n23534, n38790, n28400, n27636, n24_adj_5265, n28399, 
        n44756, n28398, n48271, n28397, n62, n28396, n27596, n27595, 
        n26240, n45738, n28395, n34636, n26243, n28394, n44743, 
        n28393, n28392, n38789, n7650, n28391, n45732, n27564, 
        n28390, n28389, n27904, n28388, n28387, n28123, n28386, 
        n48186, n28385, n27540, n28384, n45726, n45718, n7648, 
        n47237, n45712, n63, n7647, n7646, n45702, n47230, n45698, 
        n45696, n45341, n7645, n6_adj_5266, n45686, n45678, n4_adj_5267, 
        n48440, n38137, n43904, n46240, n47224, n8_adj_5268, n7_adj_5269, 
        n4_adj_5270, n14_adj_5271, n10_adj_5272, n38788, n45668, n48248, 
        n46237, n45658, n45320, n45656, n28122, n38136, n28121, 
        n46236, n6_adj_5273, n46235, n45650, n45644, n48394, n28120, 
        n28119, n26334, n38526, n38525, n38787, n38524, n38786, 
        n38785, n38523, n38784, n38522, n38783, n38521, n42180, 
        n38782, n38520, n38781, n45211, n38780, n38519, n38094, 
        n38518, n45636, n38517, n38779, n38778, n44588, n28118, 
        n28117, n45628, n38777, n38776, n45622, n38135, n38775, 
        n38774, n45616, n26879, n38516, n38515, n38514, n38513, 
        n5_adj_5274, n28116, n28115, n28114, n28113, n45606, n38134, 
        n48, n49, n50, n51, n52, n53, n54, n55, n38773, n45600, 
        n48986, n45596, n38133, n26237, n48230, n45590, n45588, 
        n38512, n28383, n28382, n28381, n28380, n28379, n28378, 
        n28377, n28376, n28373, n28372, n28368, n28365, n28362, 
        n28361, n28360, n28109, n45576, n28359, n28358, n28357, 
        n28356, n28355, n28354, n28353, n28352, n28351, n28350, 
        n28107, n28106, n28105, n28349, n28348, n28347, n28346, 
        n28345, n28344, n28343, n28342, n45570, n45568, n45562, 
        n45556, n45550, n28341, n28340, n28339, n28338, n28337, 
        n28336, n28335, n28329, n28328, n28327, n28326, n28325, 
        n28324, n28323, n28322, n28321, n28320, n28319, n28318, 
        n28317, n28316, n28315, n28314, n28313, n28312, n28311, 
        n28310, n47200, n28309, n28308, n28307, n28306, n28305, 
        n28304, n28303, n28302, n28301, n28300, n28299, n28298, 
        n28297, n28296, n38772, n38771, n38511, n38770, n28295, 
        n28294, n28293, n28292, n28291, n48384, n38132, n38769, 
        n38510, n28104, n28103, n28102, n28101, n28100, n28099, 
        n28098, n28097, n28290, n28289, n28288, n28287, n28286, 
        n28285, n28284, n28283, n38509, n38508, n38768, n28096, 
        n28095, n28094, n28093, n28092, n28091, n28090, n28089, 
        n28088, n28282, n28281, n28280, n28279, n28278, n28277, 
        n28276, n28275, n28274, n46265, n38767, n38766, n45544, 
        n38765, n38764, n45538, n45536, n38131, n38130, n38129, 
        n38763, n28273, n28272, n28271, n28270, n28269, n28268, 
        n28267, n28266, n28262, n28261, n28260, n28259, n28258, 
        n28257, n28256, n28255, n28254, n28253, n28252, n28251, 
        n28250, n28249, n28248, n28247, n28246, n28245, n28244, 
        n28243, n28242, n38507, n38762, n38506, n28241, n28240, 
        n28239, n28238, n28237, n28236, n38505, n38128, n38504, 
        n38761, n45522, n48371, n45518, n38760, n45512, n45504, 
        n10_adj_5275, n45498, n38105, n38127, n38759, n38503, n47188, 
        n47187, n38758, n26344, n47186, n45492, n26339, n38502, 
        n46211, n38501, n38500, n38757, n38499, n38126, n38756, 
        n38755, n45488, n38754, n38498, n42722, n47185, n38104, 
        n45482, n38753, n38752, n38751, n47184, n2_adj_5276, n3_adj_5277, 
        n4_adj_5278, n5_adj_5279, n6_adj_5280, n7_adj_5281, n8_adj_5282, 
        n9_adj_5283, n10_adj_5284, n11_adj_5285, n12_adj_5286, n13_adj_5287, 
        n14_adj_5288, n15_adj_5289, n16_adj_5290, n17_adj_5291, n18_adj_5292, 
        n19_adj_5293, n20_adj_5294, n21_adj_5295, n22_adj_5296, n23_adj_5297, 
        n24_adj_5298, n25_adj_5299, n26_adj_5300, n27_adj_5301, n28_adj_5302, 
        n29_adj_5303, n30_adj_5304, n31_adj_5305, n32_adj_5306, n33_adj_5307, 
        n45480, n38497, n45478, n48357, n38496, n38495, n38093, 
        n47183, n38750, n38494, n38493, n38492, n38491, n38749, 
        n45462, n47182, n38748, n38747, n45458, n39132, n38490, 
        n39131, n38746, n38489, n38745, n38744, n38488, n45454, 
        n39130, n39129, n43638, n38743, n45450, n39128, n39127, 
        n39126, n39125, n39124, n38487, n38742, n38125, n38741, 
        n39123, n39122, n39121, n38740, n39120, n39119, n38739, 
        n38486, n38092, n38738, n38737, n12_adj_5308, n39118, n45442, 
        n9_adj_5309, n38736, n39117, n4_adj_5310, n39116, n38735, 
        n39115, n39114, n39113, n38485, n39112, n38124, n39111, 
        n38734, n38733, n38123, n39110, n39109, n38732, n38484, 
        n39108, n39107, n45440, n38483, n39106, n39105, n39104, 
        n39103, n39102, n45438, n38731, n38730, n38482, n38481, 
        n38480, n38729, n45436, n38479, n38728, n38727, n45434, 
        n38726, n38725, n45432, n45430, n38724, n38723, n38722, 
        n38721, n45428, n38720, n45426, n43929, n38719, n38718, 
        n42830, n38122, n38717, n38716, n43608, n45424, n38715, 
        n38714, n45422, n38713, n38712, n45418, n38711, n38478, 
        n38477, n38476, n38475, n38710, n38709, n45416, n38708, 
        n38474, n38473, n38121, n38707, n38706, n45412, n38705, 
        n38704, n38472, n45261, n43584, n38471, n38470, n38703, 
        n38469, n38702, n38103, n38468, n38467, n45404, n38466, 
        n38465, n38102, n45402, n45400, n38701, n38101, n38120, 
        n38464, n47173, n45398, n45396, n45394, n38700, n38699, 
        n38698, n38100, n45388, n38119, n38118, n38697, n38203, 
        n38099, n38696, n45382, n43558, n38117, n43556, n38695, 
        n38091, n43554, n38694, n47171, n38693, n48326, n38463, 
        n38462, n38461, n38692, n38691, n38460, n43552, n38459, 
        n38202, n38201, n43549, n43818, n38200, n45376, n38690, 
        n34750, n18940, n38199, n45374, n38689, n38688, n38458, 
        n38457, n38116, n45368, n38687, n45366, n38115, n38456, 
        n45364, n13_adj_5311, n15_adj_5312, n19_adj_5313, n38455, 
        n21_adj_5314, n25_adj_5315, n38686, n27_adj_5316, n38685, 
        n37, n38454, n41, n38684, n7649, n38683;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5288));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5287));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5286));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_DFF dir_175 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5285));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33210_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48291));
    defparam i33210_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE dti_177 (.Q(dti), .C(CLK_c), .E(n27540), .D(dti_N_416));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i21094_3_lut (.I0(n941), .I1(n1632_adj_5263), .I2(n1633), 
            .I3(GND_net), .O(n34602));
    defparam i21094_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n45726));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n1629), .I1(n34602), .I2(n1630), .I3(n1631), 
            .O(n43846));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1582 (.I0(n1623), .I1(n43846), .I2(n1624), .I3(n45726), 
            .O(n45732));
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i33213_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n45732), 
            .O(n1653));
    defparam i33213_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i969_3_lut (.I0(n1422), .I1(n1489), 
            .I2(n1455), .I3(GND_net), .O(n1521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5284));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i4_4_lut (.I0(n7_adj_5171), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n26240), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5283));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4103[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 mux_236_i2_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20477_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_421));   // verilog/TinyFPGA_B.v(363[12:35])
    defparam i20477_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5282));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15200_3_lut (.I0(\data_out_frame[27] [1]), .I1(n26879), .I2(n27804), 
            .I3(GND_net), .O(n28711));   // verilog/coms.v(127[12] 300[6])
    defparam i15200_3_lut.LUT_INIT = 16'hcaca;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_10_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16), 
            .I3(n38184), .O(pwm_setpoint_23__N_191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_11_lut.LUT_INIT = 16'hC33C;
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .CLK_c(CLK_c), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .\state_3__N_528[1] (state_3__N_528[1]), 
            .start(start), .LED_c(LED_c), .\state[1] (state[1]), .n44588(n44588), 
            .timer({timer}), .VCC_net(VCC_net), .neopxl_color({neopxl_color}), 
            .n28137(n28137), .n27713(n27713), .n43584(n43584), .n41744(n41744), 
            .n28096(n28096), .n14(n14_adj_5172), .n28577(n28577), .n28576(n28576), 
            .n28575(n28575), .n28574(n28574), .n28573(n28573), .n28572(n28572), 
            .n28571(n28571), .n28570(n28570), .n28569(n28569), .n28568(n28568), 
            .n28567(n28567), .n28566(n28566), .n28565(n28565), .n28564(n28564), 
            .n28563(n28563), .n28562(n28562), .n28561(n28561), .n28560(n28560), 
            .n28559(n28559), .n28558(n28558), .n28557(n28557), .n28556(n28556), 
            .n28555(n28555), .n28554(n28554), .n28553(n28553), .n28552(n28552), 
            .n28551(n28551), .n28550(n28550), .n28549(n28549), .n28548(n28548), 
            .n28547(n28547), .\neo_pixel_transmitter.done_N_742 (\neo_pixel_transmitter.done_N_742 ), 
            .NEOPXL_c(NEOPXL_c), .n47171(n47171)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_LUT4 i15201_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n23568), .I3(GND_net), .O(n28712));   // verilog/coms.v(127[12] 300[6])
    defparam i15201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5281));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5243), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15202_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n23568), .I3(GND_net), .O(n28713));   // verilog/coms.v(127[12] 300[6])
    defparam i15202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5280));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5279));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33249_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48330));
    defparam i33249_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5278));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14710_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n23568), 
            .I3(GND_net), .O(n28221));   // verilog/coms.v(127[12] 300[6])
    defparam i14710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14711_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n23568), 
            .I3(GND_net), .O(n28222));   // verilog/coms.v(127[12] 300[6])
    defparam i14711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n45678));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i3_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i15203_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n23568), .I3(GND_net), .O(n28714));   // verilog/coms.v(127[12] 300[6])
    defparam i15203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15204_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n23568), .I3(GND_net), .O(n28715));   // verilog/coms.v(127[12] 300[6])
    defparam i15204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33228_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48309));
    defparam i33228_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n45650));
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'heeee;
    SB_LUT4 i21167_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n34676));
    defparam i21167_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5277));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5276));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i4_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1584 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n42634));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'hd054;
    SB_LUT4 mux_236_i5_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1585 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n45650), 
            .O(n45656));
    defparam i1_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n1529), .I1(n45656), .I2(n34676), .I3(n1530), 
            .O(n45658));
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'heccc;
    SB_LUT4 i33231_4_lut (.I0(n1522), .I1(n1521), .I2(n45658), .I3(n1523), 
            .O(n1554));
    defparam i33231_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i20257_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i20257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20256_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i20256_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20552_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i20552_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_10_add_3_11 (.CI(n38184), .I0(GND_net), .I1(n16), 
            .CO(n38185));
    SB_LUT4 unary_minus_10_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17), 
            .I3(n38183), .O(pwm_setpoint_23__N_191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n38495), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5272));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i491_2_lut (.I0(n1195), .I1(n26226), .I2(GND_net), .I3(GND_net), 
            .O(n1973));   // verilog/TinyFPGA_B.v(376[9] 382[12])
    defparam i491_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_236_i6_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i7_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32238_4_lut (.I0(n5_adj_5179), .I1(n6_adj_5266), .I2(n6976), 
            .I3(n1973), .O(n47230));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i32238_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33245_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48326));
    defparam i33245_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n38495), .I0(n1431), 
            .I1(VCC_net), .CO(n38496));
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n38494), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n38494), .I0(n1432), 
            .I1(GND_net), .CO(n38495));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n38493), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n38493), .I0(n1433), 
            .I1(VCC_net), .CO(n38494));
    SB_LUT4 i21169_4_lut (.I0(n939), .I1(n1431), .I2(n1432), .I3(n1433), 
            .O(n34678));
    defparam i21169_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n45696));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut (.I0(n1424), .I1(n1425), .I2(n1426), .I3(GND_net), 
            .O(n45702));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(n1429), .I1(n45696), .I2(n34678), .I3(n1430), 
            .O(n45698));
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'heccc;
    SB_LUT4 i33248_4_lut (.I0(n1422), .I1(n45698), .I2(n45702), .I3(n1423), 
            .O(n1455));
    defparam i33248_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i33276_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48357));
    defparam i33276_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14857_3_lut (.I0(n28056), .I1(r_Bit_Index[0]), .I2(n27767), 
            .I3(GND_net), .O(n28368));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14857_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i33290_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48371));
    defparam i33290_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14854_3_lut (.I0(n28054), .I1(r_Bit_Index_adj_5390[0]), .I2(n27763), 
            .I3(GND_net), .O(n28365));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14854_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i33303_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48384));
    defparam i33303_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i8_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20364_2_lut (.I0(n23755), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n33855));
    defparam i20364_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15171_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n27596), .I3(GND_net), .O(n28682));   // verilog/coms.v(127[12] 300[6])
    defparam i15171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14664_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n23568), .I3(GND_net), .O(n28175));   // verilog/coms.v(127[12] 300[6])
    defparam i14664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14669_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n23568), .I3(GND_net), .O(n28180));   // verilog/coms.v(127[12] 300[6])
    defparam i14669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14670_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n23568), .I3(GND_net), .O(n28181));   // verilog/coms.v(127[12] 300[6])
    defparam i14670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14671_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n23568), .I3(GND_net), .O(n28182));   // verilog/coms.v(127[12] 300[6])
    defparam i14671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14672_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n23568), .I3(GND_net), .O(n28183));   // verilog/coms.v(127[12] 300[6])
    defparam i14672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14673_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n23568), .I3(GND_net), .O(n28184));   // verilog/coms.v(127[12] 300[6])
    defparam i14673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33459_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48540));
    defparam i33459_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14665_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n23568), .I3(GND_net), .O(n28176));   // verilog/coms.v(127[12] 300[6])
    defparam i14665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14666_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n23568), .I3(GND_net), .O(n28177));   // verilog/coms.v(127[12] 300[6])
    defparam i14666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14674_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n23568), .I3(GND_net), .O(n28185));   // verilog/coms.v(127[12] 300[6])
    defparam i14674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14630_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n33899), 
            .I3(n26339), .O(n28141));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14630_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5196));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14675_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n23568), .I3(GND_net), .O(n28186));   // verilog/coms.v(127[12] 300[6])
    defparam i14675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14676_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n23568), .I3(GND_net), .O(n28187));   // verilog/coms.v(127[12] 300[6])
    defparam i14676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14677_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n23568), .I3(GND_net), .O(n28188));   // verilog/coms.v(127[12] 300[6])
    defparam i14677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14678_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n23568), .I3(GND_net), .O(n28189));   // verilog/coms.v(127[12] 300[6])
    defparam i14678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14679_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n23568), .I3(GND_net), .O(n28190));   // verilog/coms.v(127[12] 300[6])
    defparam i14679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5197));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14680_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n23568), .I3(GND_net), .O(n28191));   // verilog/coms.v(127[12] 300[6])
    defparam i14680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14681_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28192));   // verilog/coms.v(127[12] 300[6])
    defparam i14681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5198));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14682_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n23568), .I3(GND_net), .O(n28193));   // verilog/coms.v(127[12] 300[6])
    defparam i14682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14683_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28194));   // verilog/coms.v(127[12] 300[6])
    defparam i14683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14684_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28195));   // verilog/coms.v(127[12] 300[6])
    defparam i14684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14685_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28196));   // verilog/coms.v(127[12] 300[6])
    defparam i14685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14686_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28197));   // verilog/coms.v(127[12] 300[6])
    defparam i14686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33606_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48687));
    defparam i33606_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14631_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n33899), 
            .I3(n26334), .O(n28142));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14631_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5199));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14687_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n23568), .I3(GND_net), .O(n28198));   // verilog/coms.v(127[12] 300[6])
    defparam i14687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14688_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n23568), .I3(GND_net), .O(n28199));   // verilog/coms.v(127[12] 300[6])
    defparam i14688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14689_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n23568), 
            .I3(GND_net), .O(n28200));   // verilog/coms.v(127[12] 300[6])
    defparam i14689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5200));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5201));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33490_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48571));
    defparam i33490_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33426_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48507));
    defparam i33426_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14632_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28143));   // verilog/coms.v(127[12] 300[6])
    defparam i14632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14633_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n27595), 
            .I3(GND_net), .O(n28144));   // verilog/coms.v(127[12] 300[6])
    defparam i14633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14634_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n27595), 
            .I3(GND_net), .O(n28145));   // verilog/coms.v(127[12] 300[6])
    defparam i14634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14635_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n27596), .I3(GND_net), .O(n28146));   // verilog/coms.v(127[12] 300[6])
    defparam i14635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_10_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_279));   // verilog/TinyFPGA_B.v(321[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 mux_236_i9_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_238_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_10_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i10_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i33394_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48475));
    defparam i33394_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n7072), 
            .D(n1083), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n7072), 
            .D(n1082), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n7072), 
            .D(n1081), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n7072), 
            .D(n1080), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n7072), 
            .D(n1079), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n7072), 
            .D(n1078), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n7072), 
            .D(n1077), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5244), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14712_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n23568), 
            .I3(GND_net), .O(n28223));   // verilog/coms.v(127[12] 300[6])
    defparam i14712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5271));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_5271), .I2(n10_adj_5272), 
            .I3(ID[6]), .O(n26226));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i11_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i12_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14637_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28148));   // verilog/coms.v(127[12] 300[6])
    defparam i14637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \ID_READOUT_FSM.state_2__I_0_i5_2_lut  (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_5179));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam \ID_READOUT_FSM.state_2__I_0_i5_2_lut .LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33313_1_lut (.I0(n34750), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48394));
    defparam i33313_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i13_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14638_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28149));   // verilog/coms.v(127[12] 300[6])
    defparam i14638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5311));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5313));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1589 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5270));
    defparam i1_2_lut_adj_1589.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5270), .I2(delay_counter[10]), 
            .I3(n26243), .O(n44743));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5312));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_4_lut_adj_1590 (.I0(n44743), .I1(n26237), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n45211));
    defparam i2_4_lut_adj_1590.LUT_INIT = 16'hffec;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(n3220), .I1(n27_adj_5316), .I2(n3287), 
            .I3(n3237), .O(n45394));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n3227), .I1(n19_adj_5313), .I2(n3294), 
            .I3(n3237), .O(n45396));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'heefc;
    SB_LUT4 mux_238_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5268));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1593 (.I0(delay_counter[22]), .I1(n45211), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5269));
    defparam i2_4_lut_adj_1593.LUT_INIT = 16'ha8a0;
    SB_LUT4 i20478_4_lut (.I0(n7_adj_5269), .I1(delay_counter[31]), .I2(n26240), 
            .I3(n8_adj_5268), .O(n1195));   // verilog/TinyFPGA_B.v(378[14:38])
    defparam i20478_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5174));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1594 (.I0(delay_counter[28]), .I1(n12_adj_5174), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n26240));
    defparam i6_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n26237));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5168));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1595 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5167));
    defparam i6_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5167), .I1(delay_counter[2]), .I2(n14_adj_5168), 
            .I3(delay_counter[6]), .O(n26243));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4511_4_lut (.I0(n26243), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5265));
    defparam i4511_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1596 (.I0(n24_adj_5265), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n44756));
    defparam i2_4_lut_adj_1596.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1597 (.I0(n44756), .I1(delay_counter[18]), .I2(n26237), 
            .I3(GND_net), .O(n45208));
    defparam i2_3_lut_adj_1597.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1598 (.I0(delay_counter[23]), .I1(n45208), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5171));
    defparam i2_4_lut_adj_1598.LUT_INIT = 16'heaaa;
    SB_LUT4 i2_4_lut_adj_1599 (.I0(n9_adj_5309), .I1(n4_adj_5310), .I2(\FRAME_MATCHER.i_31__N_2624 ), 
            .I3(n3303), .O(n44891));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1599.LUT_INIT = 16'heefe;
    SB_LUT4 i1_4_lut_adj_1600 (.I0(n3224), .I1(n21_adj_5314), .I2(n3291), 
            .I3(n3237), .O(n45398));
    defparam i1_4_lut_adj_1600.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(n3219), .I1(n15_adj_5312), .I2(n3286), 
            .I3(n3237), .O(n45402));
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(n3221), .I1(n13_adj_5311), .I2(n3288), 
            .I3(n3237), .O(n45400));
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'heefc;
    SB_LUT4 mux_238_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(\FRAME_MATCHER.state [0]), .I1(n42830), 
            .I2(n23534), .I3(n44891), .O(n12_adj_5308));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'haf8c;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n3218), .I1(n25_adj_5315), .I2(n3285), 
            .I3(n3237), .O(n45404));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33293_4_lut (.I0(n45678), .I1(n1125), .I2(n45636), .I3(n34684), 
            .O(n1158));
    defparam i33293_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i1_4_lut_adj_1605 (.I0(\FRAME_MATCHER.state [3]), .I1(n12_adj_5308), 
            .I2(n43608), .I3(\FRAME_MATCHER.state [1]), .O(n42180));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1605.LUT_INIT = 16'hccce;
    SB_LUT4 i1_4_lut_adj_1606 (.I0(n45402), .I1(n45398), .I2(n45396), 
            .I3(n45394), .O(n45412));
    defparam i1_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n45412), .I1(n37), .I2(n45404), .I3(n45400), 
            .O(n45416));
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_236_i14_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20947_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n34453));
    defparam i20947_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i21054_4_lut (.I0(n34453), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n34562));
    defparam i21054_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 mux_236_i15_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14640_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n23568), .I3(GND_net), .O(n28151));   // verilog/coms.v(127[12] 300[6])
    defparam i14640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n47200), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5264));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n3216), .I1(n45416), .I2(n3283), .I3(n3237), 
            .O(n45418));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'heefc;
    SB_LUT4 i14641_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n23568), .I3(GND_net), .O(n28152));   // verilog/coms.v(127[12] 300[6])
    defparam i14641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21125_4_lut (.I0(n34562), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n34634));
    defparam i21125_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_i2186_3_lut (.I0(n3215), .I1(n3282), 
            .I2(n3237), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(n41), .I1(n34634), .I2(n45418), .I3(n5_adj_5264), 
            .O(n45422));
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1610 (.I0(n3214), .I1(n45422), .I2(n3281), .I3(n3237), 
            .O(n45424));
    defparam i1_4_lut_adj_1610.LUT_INIT = 16'heefc;
    SB_LUT4 i14642_3_lut (.I0(current[0]), .I1(data_adj_5377[0]), .I2(n44589), 
            .I3(GND_net), .O(n28153));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1611 (.I0(n3213), .I1(n45424), .I2(n3280), .I3(n3237), 
            .O(n45426));
    defparam i1_4_lut_adj_1611.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(n3212), .I1(n45426), .I2(n3279), .I3(n3237), 
            .O(n45428));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1613 (.I0(n3211), .I1(n45428), .I2(n3278), .I3(n3237), 
            .O(n45430));
    defparam i1_4_lut_adj_1613.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(n3210), .I1(n45430), .I2(n3277), .I3(n3237), 
            .O(n45432));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(n122_adj_5176), .I1(data_ready), .I2(state_adj_5373[1]), 
            .I3(state_adj_5373[0]), .O(n42504));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'hccd0;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n3209), .I1(n45432), .I2(n3276), .I3(n3237), 
            .O(n45434));
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(n3208), .I1(n45434), .I2(n3275), .I3(n3237), 
            .O(n45436));
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1618 (.I0(n3207), .I1(n45436), .I2(n3274), .I3(n3237), 
            .O(n45438));
    defparam i1_4_lut_adj_1618.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1619 (.I0(n3206), .I1(n45438), .I2(n3273), .I3(n3237), 
            .O(n45440));
    defparam i1_4_lut_adj_1619.LUT_INIT = 16'heefc;
    SB_LUT4 mux_236_i16_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14644_4_lut (.I0(rw), .I1(state_adj_5373[0]), .I2(state_adj_5373[1]), 
            .I3(n5615), .O(n28155));   // verilog/eeprom.v(26[8] 58[4])
    defparam i14644_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5276), .I3(n39132), .O(n2_adj_5178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(n3205), .I1(n45440), .I2(n3272), .I3(n3237), 
            .O(n45442));
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'heefc;
    SB_LUT4 i33316_4_lut (.I0(n45442), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n34750));
    defparam i33316_4_lut.LUT_INIT = 16'h1105;
    SB_CARRY add_224_14 (.CI(n38133), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n38134));
    SB_LUT4 i14645_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n23568), .I3(GND_net), .O(n28156));   // verilog/coms.v(127[12] 300[6])
    defparam i14645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5277), .I3(n39131), .O(n3_adj_5251)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n39131), 
            .I0(GND_net), .I1(n3_adj_5277), .CO(n39132));
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5278), .I3(n39130), .O(n4_adj_5222)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n38493));
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n39130), 
            .I0(GND_net), .I1(n4_adj_5278), .CO(n39131));
    SB_LUT4 i14648_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5388[1]), .I2(n18940), 
            .I3(n4_adj_5177), .O(n28159));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14648_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n48330), .I1(n1323), 
            .I2(VCC_net), .I3(n38492), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5279), .I3(n39129), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n39129), 
            .I0(GND_net), .I1(n5_adj_5279), .CO(n39130));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5280), .I3(n39128), .O(n6_adj_5229)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n39128), 
            .I0(GND_net), .I1(n6_adj_5280), .CO(n39129));
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5281), .I3(n39127), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n39127), 
            .I0(GND_net), .I1(n7_adj_5281), .CO(n39128));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5282), .I3(n39126), .O(n8_adj_5250)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n39126), 
            .I0(GND_net), .I1(n8_adj_5282), .CO(n39127));
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n38491), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14649_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n23568), .I3(GND_net), .O(n28160));   // verilog/coms.v(127[12] 300[6])
    defparam i14649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14691_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n23568), 
            .I3(GND_net), .O(n28202));   // verilog/coms.v(127[12] 300[6])
    defparam i14691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14692_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n23568), 
            .I3(GND_net), .O(n28203));   // verilog/coms.v(127[12] 300[6])
    defparam i14692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5283), .I3(n39125), .O(n9_adj_5249)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5252));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1621 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_216[0]));   // verilog/TinyFPGA_B.v(148[4] 150[7])
    defparam i1_3_lut_adj_1621.LUT_INIT = 16'h1414;
    SB_LUT4 i14650_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n23568), .I3(GND_net), .O(n28161));   // verilog/coms.v(127[12] 300[6])
    defparam i14650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n39125), 
            .I0(GND_net), .I1(n9_adj_5283), .CO(n39126));
    SB_LUT4 unary_minus_10_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5284), .I3(n39124), .O(n10_adj_5248)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n39124), 
            .I0(GND_net), .I1(n10_adj_5284), .CO(n39125));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5285), .I3(n39123), .O(n11_adj_5247)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i17_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i18_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14651_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n23568), .I3(GND_net), .O(n28162));   // verilog/coms.v(127[12] 300[6])
    defparam i14651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14652_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n23568), .I3(GND_net), .O(n28163));   // verilog/coms.v(127[12] 300[6])
    defparam i14652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14580_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n23568), .I3(GND_net), .O(n28091));   // verilog/coms.v(127[12] 300[6])
    defparam i14580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i19_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i20_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14653_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n23568), .I3(GND_net), .O(n28164));   // verilog/coms.v(127[12] 300[6])
    defparam i14653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14693_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n23568), 
            .I3(GND_net), .O(n28204));   // verilog/coms.v(127[12] 300[6])
    defparam i14693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n39123), 
            .I0(GND_net), .I1(n11_adj_5285), .CO(n39124));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5286), .I3(n39122), .O(n12_adj_5246)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14533_4_lut (.I0(n7072), .I1(n1195), .I2(n47237), .I3(n26227), 
            .O(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i14533_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14654_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n23568), .I3(GND_net), .O(n28165));   // verilog/coms.v(127[12] 300[6])
    defparam i14654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33359_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48440));
    defparam i33359_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14655_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[12]), 
            .I2(n23568), .I3(GND_net), .O(n28166));   // verilog/coms.v(127[12] 300[6])
    defparam i14655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1622 (.I0(n3228), .I1(n3218), .I2(n3219), .I3(GND_net), 
            .O(n46002));
    defparam i1_3_lut_adj_1622.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(n3224), .I1(n3227), .I2(n3226), .I3(n3220), 
            .O(n46004));
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1624 (.I0(n46004), .I1(n46002), .I2(n3222), .I3(n3223), 
            .O(n46008));
    defparam i1_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14656_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n23568), .I3(GND_net), .O(n28167));   // verilog/coms.v(127[12] 300[6])
    defparam i14656_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n39122), 
            .I0(GND_net), .I1(n12_adj_5286), .CO(n39123));
    SB_LUT4 i1_4_lut_adj_1625 (.I0(n3215), .I1(n3216), .I2(n46008), .I3(n3217), 
            .O(n46014));
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n3212), .I1(n3213), .I2(n3214), .I3(n46014), 
            .O(n46020));
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 i14694_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n23568), 
            .I3(GND_net), .O(n28205));   // verilog/coms.v(127[12] 300[6])
    defparam i14694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1627 (.I0(n3209), .I1(n3210), .I2(n3211), .I3(n46020), 
            .O(n46026));
    defparam i1_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5287), .I3(n39121), .O(n13_adj_5245)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n38491), .I0(n1324), 
            .I1(VCC_net), .CO(n38492));
    SB_LUT4 i14657_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n23568), .I3(GND_net), .O(n28168));   // verilog/coms.v(127[12] 300[6])
    defparam i14657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21127_4_lut (.I0(n957), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n34636));
    defparam i21127_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1628 (.I0(n3221), .I1(n3225), .I2(GND_net), .I3(GND_net), 
            .O(n46036));
    defparam i1_2_lut_adj_1628.LUT_INIT = 16'heeee;
    SB_LUT4 i14695_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n23568), 
            .I3(GND_net), .O(n28206));   // verilog/coms.v(127[12] 300[6])
    defparam i14695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14658_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n23568), .I3(GND_net), .O(n28169));   // verilog/coms.v(127[12] 300[6])
    defparam i14658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1629 (.I0(n3206), .I1(n3207), .I2(n3208), .I3(n46026), 
            .O(n46032));
    defparam i1_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n39121), 
            .I0(GND_net), .I1(n13_adj_5287), .CO(n39122));
    SB_LUT4 i1_4_lut_adj_1630 (.I0(n3229), .I1(n46036), .I2(n34636), .I3(n3230), 
            .O(n46038));
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5288), .I3(n39120), .O(n14_adj_5244)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5202));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5203));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i21_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i33363_4_lut (.I0(n3204), .I1(n46038), .I2(n46032), .I3(n3205), 
            .O(n3237));
    defparam i33363_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_238_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_236_i22_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14659_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n23568), .I3(GND_net), .O(n28170));   // verilog/coms.v(127[12] 300[6])
    defparam i14659_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n39120), 
            .I0(GND_net), .I1(n14_adj_5288), .CO(n39121));
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14660_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n23568), .I3(GND_net), .O(n28171));   // verilog/coms.v(127[12] 300[6])
    defparam i14660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14661_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n23568), .I3(GND_net), .O(n28172));   // verilog/coms.v(127[12] 300[6])
    defparam i14661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14662_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n23568), .I3(GND_net), .O(n28173));   // verilog/coms.v(127[12] 300[6])
    defparam i14662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14663_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n23568), .I3(GND_net), .O(n28174));   // verilog/coms.v(127[12] 300[6])
    defparam i14663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15172_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n27596), .I3(GND_net), .O(n28683));   // verilog/coms.v(127[12] 300[6])
    defparam i15172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14696_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n23568), 
            .I3(GND_net), .O(n28207));   // verilog/coms.v(127[12] 300[6])
    defparam i14696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15173_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n27596), .I3(GND_net), .O(n28684));   // verilog/coms.v(127[12] 300[6])
    defparam i15173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15174_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28685));   // verilog/coms.v(127[12] 300[6])
    defparam i15174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15175_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28686));   // verilog/coms.v(127[12] 300[6])
    defparam i15175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15176_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n27596), .I3(GND_net), .O(n28687));   // verilog/coms.v(127[12] 300[6])
    defparam i15176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15177_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n27596), .I3(GND_net), .O(n28688));   // verilog/coms.v(127[12] 300[6])
    defparam i15177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14697_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n23568), 
            .I3(GND_net), .O(n28208));   // verilog/coms.v(127[12] 300[6])
    defparam i14697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33638_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48719));
    defparam i33638_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15178_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n27596), .I3(GND_net), .O(n28689));   // verilog/coms.v(127[12] 300[6])
    defparam i15178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15179_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n27596), .I3(GND_net), .O(n28690));   // verilog/coms.v(127[12] 300[6])
    defparam i15179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1631 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam i4_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1632 (.I0(control_mode[6]), .I1(n10), .I2(control_mode[2]), 
            .I3(GND_net), .O(n26344));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam i5_3_lut_adj_1632.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5289), .I3(n39119), .O(n15_adj_5243)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n39119), 
            .I0(GND_net), .I1(n15_adj_5289), .CO(n39120));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5290), .I3(n39118), .O(n16_adj_5242)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n39118), 
            .I0(GND_net), .I1(n16_adj_5290), .CO(n39119));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5291), .I3(n39117), .O(n17_adj_5241)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n39117), 
            .I0(GND_net), .I1(n17_adj_5291), .CO(n39118));
    SB_LUT4 i15180_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28691));   // verilog/coms.v(127[12] 300[6])
    defparam i15180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5292), .I3(n39116), .O(n18_adj_5240)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_236_i23_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n39116), 
            .I0(GND_net), .I1(n18_adj_5292), .CO(n39117));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5293), .I3(n39115), .O(n19_adj_5239)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1633 (.I0(n26211), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5173));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_adj_1633.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_adj_1634 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n26344), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i2_3_lut_adj_1634.LUT_INIT = 16'hfdfd;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_5173), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n39115), 
            .I0(GND_net), .I1(n19_adj_5293), .CO(n39116));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5294), .I3(n39114), .O(n20_adj_5238)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n39114), 
            .I0(GND_net), .I1(n20_adj_5294), .CO(n39115));
    SB_CARRY unary_minus_10_add_3_10 (.CI(n38183), .I0(GND_net), .I1(n17), 
            .CO(n38184));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5295), .I3(n39113), .O(n21_adj_5237)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15181_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n27596), .I3(GND_net), .O(n28692));   // verilog/coms.v(127[12] 300[6])
    defparam i15181_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n39113), 
            .I0(GND_net), .I1(n21_adj_5295), .CO(n39114));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5296), .I3(n39112), .O(n22_adj_5236)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n39112), 
            .I0(GND_net), .I1(n22_adj_5296), .CO(n39113));
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5297), .I3(n39111), .O(n23_adj_5235)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15182_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28693));   // verilog/coms.v(127[12] 300[6])
    defparam i15182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n38490), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n39111), 
            .I0(GND_net), .I1(n23_adj_5297), .CO(n39112));
    SB_LUT4 add_145_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n38093), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5298), .I3(n39110), .O(n24_adj_5234)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n39110), 
            .I0(GND_net), .I1(n24_adj_5298), .CO(n39111));
    SB_LUT4 mux_236_i24_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5299), .I3(n39109), .O(n25_adj_5233)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n39109), 
            .I0(GND_net), .I1(n25_adj_5299), .CO(n39110));
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n38490), .I0(n1325), 
            .I1(VCC_net), .CO(n38491));
    SB_LUT4 add_224_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n38132), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5300), .I3(n39108), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15183_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n27596), .I3(GND_net), .O(n28694));   // verilog/coms.v(127[12] 300[6])
    defparam i15183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21058_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n34566));
    defparam i21058_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15184_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n27596), .I3(GND_net), .O(n28695));   // verilog/coms.v(127[12] 300[6])
    defparam i15184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n38489), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15185_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n27596), .I3(GND_net), .O(n28696));   // verilog/coms.v(127[12] 300[6])
    defparam i15185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(n3129), .I1(n34566), .I2(n3130), .I3(n3131), 
            .O(n43929));
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'ha080;
    SB_LUT4 i15186_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n27596), .I3(GND_net), .O(n28697));   // verilog/coms.v(127[12] 300[6])
    defparam i15186_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n7072), 
            .D(n1086), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n39108), 
            .I0(GND_net), .I1(n26_adj_5300), .CO(n39109));
    SB_LUT4 i1_4_lut_adj_1636 (.I0(n3121), .I1(n3124), .I2(n3127), .I3(n3128), 
            .O(n45450));
    defparam i1_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i33578_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48659));
    defparam i33578_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15187_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28698));   // verilog/coms.v(127[12] 300[6])
    defparam i15187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5301), .I3(n39107), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15188_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28699));   // verilog/coms.v(127[12] 300[6])
    defparam i15188_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n39107), 
            .I0(GND_net), .I1(n27_adj_5301), .CO(n39108));
    SB_LUT4 i15189_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n27596), .I3(GND_net), .O(n28700));   // verilog/coms.v(127[12] 300[6])
    defparam i15189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1637 (.I0(n3117), .I1(n45450), .I2(n3118), .I3(n3122), 
            .O(n45454));
    defparam i1_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1638 (.I0(n43929), .I1(n3115), .I2(n3120), .I3(n3119), 
            .O(n45766));
    defparam i1_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5302), .I3(n39106), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n39106), 
            .I0(GND_net), .I1(n28_adj_5302), .CO(n39107));
    SB_LUT4 i1_4_lut_adj_1639 (.I0(n3116), .I1(n3125), .I2(n3123), .I3(n3126), 
            .O(n45712));
    defparam i1_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5303), .I3(n39105), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n45766), .I1(n3112), .I2(n3111), .I3(n45454), 
            .O(n45458));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n39105), 
            .I0(GND_net), .I1(n29_adj_5303), .CO(n39106));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5304), .I3(n39104), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n38489), .I0(n1326), 
            .I1(VCC_net), .CO(n38490));
    SB_CARRY add_224_13 (.CI(n38132), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n38133));
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n7072), 
            .D(n1093), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n39104), 
            .I0(GND_net), .I1(n30_adj_5304), .CO(n39105));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5305), .I3(n39103), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n38488), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n38488), .I0(n1327), 
            .I1(VCC_net), .CO(n38489));
    SB_LUT4 i15190_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n27596), .I3(GND_net), .O(n28701));   // verilog/coms.v(127[12] 300[6])
    defparam i15190_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n39103), 
            .I0(GND_net), .I1(n31_adj_5305), .CO(n39104));
    SB_LUT4 i1_4_lut_adj_1641 (.I0(n3110), .I1(n3113), .I2(n3114), .I3(n45712), 
            .O(n45718));
    defparam i1_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5306), .I3(n39102), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(n3108), .I1(n45718), .I2(n45458), .I3(n3109), 
            .O(n45462));
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n39102), 
            .I0(GND_net), .I1(n32_adj_5306), .CO(n39103));
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n7072), 
            .D(n1092), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5307), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5307), .CO(n39102));
    SB_LUT4 i33397_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n45462), 
            .O(n3138));
    defparam i33397_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i14387_2_lut (.I0(n27564), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i14387_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14698_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n23568), 
            .I3(GND_net), .O(n28209));   // verilog/coms.v(127[12] 300[6])
    defparam i14698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n38487), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14699_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n23568), 
            .I3(GND_net), .O(n28210));   // verilog/coms.v(127[12] 300[6])
    defparam i14699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14700_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n23568), 
            .I3(GND_net), .O(n28211));   // verilog/coms.v(127[12] 300[6])
    defparam i14700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15191_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n27596), .I3(GND_net), .O(n28702));   // verilog/coms.v(127[12] 300[6])
    defparam i15191_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n38487), .I0(n1328), 
            .I1(VCC_net), .CO(n38488));
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32988_4_lut (.I0(commutation_state[1]), .I1(n23755), .I2(dti), 
            .I3(commutation_state[2]), .O(n27564));
    defparam i32988_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i14701_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n23568), 
            .I3(GND_net), .O(n28212));   // verilog/coms.v(127[12] 300[6])
    defparam i14701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n38486), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15192_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n27596), .I3(GND_net), .O(n28703));   // verilog/coms.v(127[12] 300[6])
    defparam i15192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14702_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n23568), 
            .I3(GND_net), .O(n28213));   // verilog/coms.v(127[12] 300[6])
    defparam i14702_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n38486), .I0(n1329), 
            .I1(GND_net), .CO(n38487));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n38485), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n38131), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15193_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28704));   // verilog/coms.v(127[12] 300[6])
    defparam i15193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15194_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28705));   // verilog/coms.v(127[12] 300[6])
    defparam i15194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n38485), .I0(n1330), 
            .I1(GND_net), .CO(n38486));
    SB_LUT4 i15195_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n27596), .I3(GND_net), .O(n28706));   // verilog/coms.v(127[12] 300[6])
    defparam i15195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33553_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48634));
    defparam i33553_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14703_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n23568), 
            .I3(GND_net), .O(n28214));   // verilog/coms.v(127[12] 300[6])
    defparam i14703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14704_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n23568), 
            .I3(GND_net), .O(n28215));   // verilog/coms.v(127[12] 300[6])
    defparam i14704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14705_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n23568), 
            .I3(GND_net), .O(n28216));   // verilog/coms.v(127[12] 300[6])
    defparam i14705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n38484), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n38484), .I0(n1331), 
            .I1(VCC_net), .CO(n38485));
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096_adj_5256), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_8 (.CI(n38127), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n38128));
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n7072), 
            .D(n1085), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i15196_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n27596), .I3(GND_net), .O(n28707));   // verilog/coms.v(127[12] 300[6])
    defparam i15196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i15197_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n27596), .I3(GND_net), .O(n28708));   // verilog/coms.v(127[12] 300[6])
    defparam i15197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195_adj_5262), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n38101), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14581_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n23568), .I3(GND_net), .O(n28092));   // verilog/coms.v(127[12] 300[6])
    defparam i14581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15198_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n27596), .I3(GND_net), .O(n28709));   // verilog/coms.v(127[12] 300[6])
    defparam i15198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n38483), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n7072), 
            .D(n1108), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n38483), .I0(n1332), 
            .I1(GND_net), .CO(n38484));
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n38482), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14714_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n23568), .I3(GND_net), .O(n28225));   // verilog/coms.v(127[12] 300[6])
    defparam i14714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14706_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n23568), 
            .I3(GND_net), .O(n28217));   // verilog/coms.v(127[12] 300[6])
    defparam i14706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15199_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n27596), .I3(GND_net), .O(n28710));   // verilog/coms.v(127[12] 300[6])
    defparam i15199_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n38482), .I0(n1333), 
            .I1(VCC_net), .CO(n38483));
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n7072), 
            .D(n1084), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n38482));
    SB_LUT4 unary_minus_10_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n38182), .O(pwm_setpoint_23__N_191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n38126), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n48357), .I1(n1224), 
            .I2(VCC_net), .I3(n38481), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n38480), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n38480), .I0(n1225), 
            .I1(VCC_net), .CO(n38481));
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(n3026), .I1(n3019), .I2(n3027), .I3(n3023), 
            .O(n45918));
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1644 (.I0(n3020), .I1(n3025), .I2(n3022), .I3(n3024), 
            .O(n45916));
    defparam i1_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n38479), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n38479), .I0(n1226), 
            .I1(VCC_net), .CO(n38480));
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n38478), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n38478), .I0(n1227), 
            .I1(VCC_net), .CO(n38479));
    SB_CARRY unary_minus_10_add_3_9 (.CI(n38182), .I0(GND_net), .I1(n18), 
            .CO(n38183));
    SB_LUT4 i1_3_lut_adj_1645 (.I0(n45918), .I1(n3021), .I2(n3028), .I3(GND_net), 
            .O(n45920));
    defparam i1_3_lut_adj_1645.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n38477), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21060_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n34568));
    defparam i21060_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n38477), .I0(n1228), 
            .I1(VCC_net), .CO(n38478));
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n38476), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n38476), .I0(n1229), 
            .I1(GND_net), .CO(n38477));
    SB_LUT4 unary_minus_10_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19), 
            .I3(n38181), .O(pwm_setpoint_23__N_191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n3017), .I1(n3018), .I2(n45920), .I3(n45916), 
            .O(n45926));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n3029), .I1(n34568), .I2(n3030), .I3(n3031), 
            .O(n43969));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n38475), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_8 (.CI(n38181), .I0(GND_net), .I1(n19), 
            .CO(n38182));
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n3015), .I1(n43969), .I2(n3016), .I3(n45926), 
            .O(n45932));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n45932), 
            .O(n45938));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n45938), 
            .O(n45944));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i33430_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n45944), 
            .O(n3039));
    defparam i33430_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n38475), .I0(n1230), 
            .I1(GND_net), .CO(n38476));
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n38474), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n38474), .I0(n1231), 
            .I1(VCC_net), .CO(n38475));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n38473), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14724_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n23568), .I3(GND_net), .O(n28235));   // verilog/coms.v(127[12] 300[6])
    defparam i14724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14725_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28236));   // verilog/coms.v(127[12] 300[6])
    defparam i14725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14726_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n23568), .I3(GND_net), .O(n28237));   // verilog/coms.v(127[12] 300[6])
    defparam i14726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14727_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28238));   // verilog/coms.v(127[12] 300[6])
    defparam i14727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33520_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48601));
    defparam i33520_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n38180), .O(pwm_setpoint_23__N_191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n38473), .I0(n1232), 
            .I1(GND_net), .CO(n38474));
    SB_LUT4 i14576_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n23568), .I3(GND_net), .O(n28087));   // verilog/coms.v(127[12] 300[6])
    defparam i14576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n38472), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14728_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28239));   // verilog/coms.v(127[12] 300[6])
    defparam i14728_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n38472), .I0(n1233), 
            .I1(VCC_net), .CO(n38473));
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14729_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28240));   // verilog/coms.v(127[12] 300[6])
    defparam i14729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5166));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14582_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n23568), .I3(GND_net), .O(n28093));   // verilog/coms.v(127[12] 300[6])
    defparam i14582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14583_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n23568), .I3(GND_net), .O(n28094));   // verilog/coms.v(127[12] 300[6])
    defparam i14583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14730_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n23568), .I3(GND_net), .O(n28241));   // verilog/coms.v(127[12] 300[6])
    defparam i14730_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n38472));
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n48371), .I1(n1125), 
            .I2(VCC_net), .I3(n38471), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14584_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n23568), .I3(GND_net), .O(n28095));   // verilog/coms.v(127[12] 300[6])
    defparam i14584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14731_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n23568), .I3(GND_net), .O(n28242));   // verilog/coms.v(127[12] 300[6])
    defparam i14731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14732_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28243));   // verilog/coms.v(127[12] 300[6])
    defparam i14732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14733_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4087[0]), 
            .I3(n122_adj_5176), .O(n28244));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14733_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14585_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n44588), .I3(GND_net), .O(n28096));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14586_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n23568), .I3(GND_net), .O(n28097));   // verilog/coms.v(127[12] 300[6])
    defparam i14586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n38470), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14587_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n23568), .I3(GND_net), .O(n28098));   // verilog/coms.v(127[12] 300[6])
    defparam i14587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14734_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28245));   // verilog/coms.v(127[12] 300[6])
    defparam i14734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14588_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n23568), .I3(GND_net), .O(n28099));   // verilog/coms.v(127[12] 300[6])
    defparam i14588_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_12 (.CI(n38131), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n38132));
    SB_LUT4 i14589_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n23568), .I3(GND_net), .O(n28100));   // verilog/coms.v(127[12] 300[6])
    defparam i14589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n38470), .I0(n1126), 
            .I1(VCC_net), .CO(n38471));
    SB_CARRY unary_minus_10_add_3_7 (.CI(n38180), .I0(GND_net), .I1(n20), 
            .CO(n38181));
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14735_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28246));   // verilog/coms.v(127[12] 300[6])
    defparam i14735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14736_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n23568), .I3(GND_net), .O(n28247));   // verilog/coms.v(127[12] 300[6])
    defparam i14736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n38469), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14590_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n23568), .I3(GND_net), .O(n28101));   // verilog/coms.v(127[12] 300[6])
    defparam i14590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_224_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n38130), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n38469), .I0(n1127), 
            .I1(VCC_net), .CO(n38470));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n38468), .O(n1195_adj_5262)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14715_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n23568), .I3(GND_net), .O(n28226));   // verilog/coms.v(127[12] 300[6])
    defparam i14715_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_11 (.CI(n38130), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n38131));
    SB_LUT4 unary_minus_10_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n38179), .O(pwm_setpoint_23__N_191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14591_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n23568), .I3(GND_net), .O(n28102));   // verilog/coms.v(127[12] 300[6])
    defparam i14591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14592_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n23568), .I3(GND_net), .O(n28103));   // verilog/coms.v(127[12] 300[6])
    defparam i14592_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n38468), .I0(n1128), 
            .I1(VCC_net), .CO(n38469));
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n38467), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14593_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n23568), .I3(GND_net), .O(n28104));   // verilog/coms.v(127[12] 300[6])
    defparam i14593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14737_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28248));   // verilog/coms.v(127[12] 300[6])
    defparam i14737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14738_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28249));   // verilog/coms.v(127[12] 300[6])
    defparam i14738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14739_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28250));   // verilog/coms.v(127[12] 300[6])
    defparam i14739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14594_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n23568), .I3(GND_net), .O(n28105));   // verilog/coms.v(127[12] 300[6])
    defparam i14594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14595_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n23568), .I3(GND_net), .O(n28106));   // verilog/coms.v(127[12] 300[6])
    defparam i14595_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n38467), .I0(n1129), 
            .I1(GND_net), .CO(n38468));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n38466), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_6 (.CI(n38179), .I0(GND_net), .I1(n21), 
            .CO(n38180));
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n38466), .I0(n1130), 
            .I1(GND_net), .CO(n38467));
    SB_LUT4 i14596_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n45341), .I3(GND_net), 
            .O(n28107));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14596_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n38465), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n38465), .I0(n1131), 
            .I1(VCC_net), .CO(n38466));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n38464), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14740_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28251));   // verilog/coms.v(127[12] 300[6])
    defparam i14740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14707_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n23568), 
            .I3(GND_net), .O(n28218));   // verilog/coms.v(127[12] 300[6])
    defparam i14707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n38129), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32208_2_lut (.I0(start), .I1(n14_adj_5172), .I2(GND_net), 
            .I3(GND_net), .O(n47173));   // verilog/neopixel.v(35[12] 117[6])
    defparam i32208_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31_4_lut (.I0(n47173), .I1(n47171), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n41744));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_10 (.CI(n38129), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n38130));
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n38464), .I0(n1132), 
            .I1(GND_net), .CO(n38465));
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n38463), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n38463), .I0(n1133), 
            .I1(VCC_net), .CO(n38464));
    SB_LUT4 unary_minus_10_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n38178), .O(pwm_setpoint_23__N_191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_5 (.CI(n38178), .I0(GND_net), .I1(n22), 
            .CO(n38179));
    SB_LUT4 unary_minus_10_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23), 
            .I3(n38177), .O(pwm_setpoint_23__N_191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14598_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28109));   // verilog/coms.v(127[12] 300[6])
    defparam i14598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14708_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n23568), 
            .I3(GND_net), .O(n28219));   // verilog/coms.v(127[12] 300[6])
    defparam i14708_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n38463));
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n38462), .O(n1093_adj_5253)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_742 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14602_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[1]), .I2(n5_adj_5212), 
            .I3(n26390), .O(n28113));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14602_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14603_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[2]), .I2(n5_adj_5207), 
            .I3(n26390), .O(n28114));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14603_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14604_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[3]), .I2(n33894), 
            .I3(n26390), .O(n28115));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14604_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14605_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[4]), .I2(n9_adj_5230), 
            .I3(n26385), .O(n28116));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14605_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14741_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n23568), .I3(GND_net), .O(n28252));   // verilog/coms.v(127[12] 300[6])
    defparam i14741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n38128), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n38461), .O(n1094_adj_5254)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14606_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[5]), .I2(n5_adj_5212), 
            .I3(n26385), .O(n28117));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14606_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_224_9 (.CI(n38128), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n38129));
    SB_CARRY unary_minus_10_add_3_4 (.CI(n38177), .I0(GND_net), .I1(n23), 
            .CO(n38178));
    SB_LUT4 i14607_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[6]), .I2(n5_adj_5207), 
            .I3(n26385), .O(n28118));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14607_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_10_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n38176), .O(pwm_setpoint_23__N_191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14608_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[7]), .I2(n33894), 
            .I3(n26385), .O(n28119));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14608_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n38461), .I0(n1027), 
            .I1(VCC_net), .CO(n38462));
    SB_CARRY add_145_13 (.CI(n38101), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n38102));
    SB_LUT4 i14742_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n23568), .I3(GND_net), .O(n28253));   // verilog/coms.v(127[12] 300[6])
    defparam i14742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14743_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n23568), .I3(GND_net), .O(n28254));   // verilog/coms.v(127[12] 300[6])
    defparam i14743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14609_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[8]), .I2(n9_adj_5230), 
            .I3(n26380), .O(n28120));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14744_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n23568), .I3(GND_net), .O(n28255));   // verilog/coms.v(127[12] 300[6])
    defparam i14744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14745_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n23568), .I3(GND_net), .O(n28256));   // verilog/coms.v(127[12] 300[6])
    defparam i14745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14610_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[9]), .I2(n5_adj_5212), 
            .I3(n26380), .O(n28121));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14610_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14611_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[10]), .I2(n5_adj_5207), 
            .I3(n26380), .O(n28122));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14746_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n23568), .I3(GND_net), .O(n28257));   // verilog/coms.v(127[12] 300[6])
    defparam i14746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14747_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n23568), .I3(GND_net), .O(n28258));   // verilog/coms.v(127[12] 300[6])
    defparam i14747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14612_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[11]), .I2(n33894), 
            .I3(n26380), .O(n28123));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14612_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14748_4_lut (.I0(state_7__N_4103[3]), .I1(data[0]), .I2(n10_adj_5275), 
            .I3(n26372), .O(n28259));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14748_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n38460), .O(n1095_adj_5255)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14749_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n23568), .I3(GND_net), .O(n28260));   // verilog/coms.v(127[12] 300[6])
    defparam i14749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14750_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n23568), .I3(GND_net), .O(n28261));   // verilog/coms.v(127[12] 300[6])
    defparam i14750_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n38460), .I0(n1028), 
            .I1(VCC_net), .CO(n38461));
    SB_CARRY add_224_7 (.CI(n38126), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n38127));
    SB_CARRY add_145_5 (.CI(n38093), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n38094));
    SB_LUT4 i14751_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n23568), .I3(GND_net), .O(n28262));   // verilog/coms.v(127[12] 300[6])
    defparam i14751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n2922), .I1(n2926), .I2(n2921), .I3(n2928), 
            .O(n45480));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_145_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n38100), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14755_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28266));   // verilog/coms.v(127[12] 300[6])
    defparam i14755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n5_adj_5179), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n1973), .I3(read_N_421), .O(n25_adj_5169));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'h7350;
    SB_LUT4 i14756_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28267));   // verilog/coms.v(127[12] 300[6])
    defparam i14756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n2924), .I1(n2920), .I2(n2927), .I3(n2925), 
            .O(n45478));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1654 (.I0(n45480), .I1(n2919), .I2(n2923), .I3(GND_net), 
            .O(n45482));
    defparam i1_3_lut_adj_1654.LUT_INIT = 16'hfefe;
    SB_LUT4 i14757_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28268));   // verilog/coms.v(127[12] 300[6])
    defparam i14757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31188_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n46211));
    defparam i31188_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_10_add_3_3 (.CI(n38176), .I0(GND_net), .I1(n24), 
            .CO(n38177));
    SB_LUT4 i21133_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n34642));
    defparam i21133_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_224_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n38125), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33325_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6976), .I2(n46211), 
            .I3(n25_adj_5169), .O(n17_adj_5170));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i33325_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i14758_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28269));   // verilog/coms.v(127[12] 300[6])
    defparam i14758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14759_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28270));   // verilog/coms.v(127[12] 300[6])
    defparam i14759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14760_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28271));   // verilog/coms.v(127[12] 300[6])
    defparam i14760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14761_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28272));   // verilog/coms.v(127[12] 300[6])
    defparam i14761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14762_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28273));   // verilog/coms.v(127[12] 300[6])
    defparam i14762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n2917), .I1(n2918), .I2(n45482), .I3(n45478), 
            .O(n45488));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(n2929), .I1(n2930), .I2(GND_net), .I3(GND_net), 
            .O(n45990));
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'h8888;
    SB_LUT4 i14763_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28274));   // verilog/coms.v(127[12] 300[6])
    defparam i14763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14613_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[12]), .I2(n9_adj_5230), 
            .I3(n26377), .O(n28124));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14613_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14764_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28275));   // verilog/coms.v(127[12] 300[6])
    defparam i14764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14765_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28276));   // verilog/coms.v(127[12] 300[6])
    defparam i14765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14766_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28277));   // verilog/coms.v(127[12] 300[6])
    defparam i14766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14767_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28278));   // verilog/coms.v(127[12] 300[6])
    defparam i14767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14768_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28279));   // verilog/coms.v(127[12] 300[6])
    defparam i14768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14769_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28280));   // verilog/coms.v(127[12] 300[6])
    defparam i14769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14770_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28281));   // verilog/coms.v(127[12] 300[6])
    defparam i14770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14771_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28282));   // verilog/coms.v(127[12] 300[6])
    defparam i14771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14772_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28283));   // verilog/coms.v(127[12] 300[6])
    defparam i14772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14773_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28284));   // verilog/coms.v(127[12] 300[6])
    defparam i14773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14774_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28285));   // verilog/coms.v(127[12] 300[6])
    defparam i14774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n45990), .I1(n2916), .I2(n45488), .I3(n34642), 
            .O(n45492));
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1658 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n45492), 
            .O(n45498));
    defparam i1_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n45498), 
            .O(n45504));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i14775_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28286));   // verilog/coms.v(127[12] 300[6])
    defparam i14775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14776_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28287));   // verilog/coms.v(127[12] 300[6])
    defparam i14776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33462_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n45504), 
            .O(n2940));
    defparam i33462_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5307));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14777_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28288));   // verilog/coms.v(127[12] 300[6])
    defparam i14777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5306));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14778_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n23568), .I3(GND_net), .O(n28289));   // verilog/coms.v(127[12] 300[6])
    defparam i14778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14779_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n23568), .I3(GND_net), .O(n28290));   // verilog/coms.v(127[12] 300[6])
    defparam i14779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(pwm_setpoint_23__N_191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14780_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n23568), .I3(GND_net), .O(n28291));   // verilog/coms.v(127[12] 300[6])
    defparam i14780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14781_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n23568), .I3(GND_net), .O(n28292));   // verilog/coms.v(127[12] 300[6])
    defparam i14781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n38459), .O(n1096_adj_5256)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(244[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14782_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n23568), .I3(GND_net), .O(n28293));   // verilog/coms.v(127[12] 300[6])
    defparam i14782_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n7072), 
            .D(n1107), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14783_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n23568), .I3(GND_net), .O(n28294));   // verilog/coms.v(127[12] 300[6])
    defparam i14783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14784_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n23568), .I3(GND_net), .O(n28295));   // verilog/coms.v(127[12] 300[6])
    defparam i14784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14785_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n23568), .I3(GND_net), .O(n28296));   // verilog/coms.v(127[12] 300[6])
    defparam i14785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5305));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14786_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n23568), .I3(GND_net), .O(n28297));   // verilog/coms.v(127[12] 300[6])
    defparam i14786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14787_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n23568), .I3(GND_net), .O(n28298));   // verilog/coms.v(127[12] 300[6])
    defparam i14787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14788_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n23568), .I3(GND_net), .O(n28299));   // verilog/coms.v(127[12] 300[6])
    defparam i14788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5304));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14789_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n23568), .I3(GND_net), .O(n28300));   // verilog/coms.v(127[12] 300[6])
    defparam i14789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_10_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n38176));
    SB_LUT4 i14790_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n23568), .I3(GND_net), .O(n28301));   // verilog/coms.v(127[12] 300[6])
    defparam i14790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14791_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n23568), .I3(GND_net), .O(n28302));   // verilog/coms.v(127[12] 300[6])
    defparam i14791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14792_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n23568), .I3(GND_net), .O(n28303));   // verilog/coms.v(127[12] 300[6])
    defparam i14792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14793_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n23568), .I3(GND_net), .O(n28304));   // verilog/coms.v(127[12] 300[6])
    defparam i14793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14794_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n23568), .I3(GND_net), .O(n28305));   // verilog/coms.v(127[12] 300[6])
    defparam i14794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14795_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n23568), .I3(GND_net), .O(n28306));   // verilog/coms.v(127[12] 300[6])
    defparam i14795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14796_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n23568), .I3(GND_net), .O(n28307));   // verilog/coms.v(127[12] 300[6])
    defparam i14796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14797_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n23568), .I3(GND_net), .O(n28308));   // verilog/coms.v(127[12] 300[6])
    defparam i14797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14709_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n23568), 
            .I3(GND_net), .O(n28220));   // verilog/coms.v(127[12] 300[6])
    defparam i14709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5303));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14798_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n23568), .I3(GND_net), .O(n28309));   // verilog/coms.v(127[12] 300[6])
    defparam i14798_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_12 (.CI(n38100), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n38101));
    SB_LUT4 i14799_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n23568), .I3(GND_net), .O(n28310));   // verilog/coms.v(127[12] 300[6])
    defparam i14799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14800_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n23568), .I3(GND_net), .O(n28311));   // verilog/coms.v(127[12] 300[6])
    defparam i14800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14801_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n23568), .I3(GND_net), .O(n28312));   // verilog/coms.v(127[12] 300[6])
    defparam i14801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14802_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n23568), .I3(GND_net), .O(n28313));   // verilog/coms.v(127[12] 300[6])
    defparam i14802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5302));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14803_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n23568), .I3(GND_net), .O(n28314));   // verilog/coms.v(127[12] 300[6])
    defparam i14803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14804_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n23568), .I3(GND_net), .O(n28315));   // verilog/coms.v(127[12] 300[6])
    defparam i14804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14805_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n23568), .I3(GND_net), .O(n28316));   // verilog/coms.v(127[12] 300[6])
    defparam i14805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5301));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14806_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n23568), .I3(GND_net), .O(n28317));   // verilog/coms.v(127[12] 300[6])
    defparam i14806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14807_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n23568), .I3(GND_net), .O(n28318));   // verilog/coms.v(127[12] 300[6])
    defparam i14807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14808_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n23568), .I3(GND_net), .O(n28319));   // verilog/coms.v(127[12] 300[6])
    defparam i14808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14809_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n23568), .I3(GND_net), .O(n28320));   // verilog/coms.v(127[12] 300[6])
    defparam i14809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14810_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n23568), .I3(GND_net), .O(n28321));   // verilog/coms.v(127[12] 300[6])
    defparam i14810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14811_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n23568), .I3(GND_net), .O(n28322));   // verilog/coms.v(127[12] 300[6])
    defparam i14811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14812_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n23568), .I3(GND_net), .O(n28323));   // verilog/coms.v(127[12] 300[6])
    defparam i14812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14813_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n23568), .I3(GND_net), .O(n28324));   // verilog/coms.v(127[12] 300[6])
    defparam i14813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14814_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n23568), .I3(GND_net), .O(n28325));   // verilog/coms.v(127[12] 300[6])
    defparam i14814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32716_3_lut (.I0(n2627), .I1(n2694), .I2(n2643), .I3(GND_net), 
            .O(n2726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32717_3_lut (.I0(n2726), .I1(n2793), .I2(n2742), .I3(GND_net), 
            .O(n2825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14815_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28326));   // verilog/coms.v(127[12] 300[6])
    defparam i14815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5300));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14816_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n23568), .I3(GND_net), .O(n28327));   // verilog/coms.v(127[12] 300[6])
    defparam i14816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14817_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28328));   // verilog/coms.v(127[12] 300[6])
    defparam i14817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14713_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n23568), 
            .I3(GND_net), .O(n28224));   // verilog/coms.v(127[12] 300[6])
    defparam i14713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14818_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28329));   // verilog/coms.v(127[12] 300[6])
    defparam i14818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n45320));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32714_3_lut (.I0(n2624), .I1(n2691), .I2(n2643), .I3(GND_net), 
            .O(n2723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14824_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n23568), .I3(GND_net), .O(n28335));   // verilog/coms.v(127[12] 300[6])
    defparam i14824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14825_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n23568), .I3(GND_net), .O(n28336));   // verilog/coms.v(127[12] 300[6])
    defparam i14825_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dti_counter_2188__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n7072), 
            .D(n1106), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14614_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[15]), .I2(n33894), 
            .I3(n26377), .O(n28125));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14614_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14826_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n23568), .I3(GND_net), .O(n28337));   // verilog/coms.v(127[12] 300[6])
    defparam i14826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15101_3_lut (.I0(current[12]), .I1(data_adj_5377[12]), .I2(n44589), 
            .I3(GND_net), .O(n28612));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14827_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n23568), .I3(GND_net), .O(n28338));   // verilog/coms.v(127[12] 300[6])
    defparam i14827_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n7072), 
            .D(n1091), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14828_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n23568), .I3(GND_net), .O(n28339));   // verilog/coms.v(127[12] 300[6])
    defparam i14828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14829_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n23568), .I3(GND_net), .O(n28340));   // verilog/coms.v(127[12] 300[6])
    defparam i14829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32715_3_lut (.I0(n2723), .I1(n2790), .I2(n2742), .I3(GND_net), 
            .O(n2822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14830_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n23568), .I3(GND_net), .O(n28341));   // verilog/coms.v(127[12] 300[6])
    defparam i14830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14831_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n23568), .I3(GND_net), .O(n28342));   // verilog/coms.v(127[12] 300[6])
    defparam i14831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14832_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n23568), .I3(GND_net), .O(n28343));   // verilog/coms.v(127[12] 300[6])
    defparam i14832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14833_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n23568), .I3(GND_net), .O(n28344));   // verilog/coms.v(127[12] 300[6])
    defparam i14833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14834_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n23568), .I3(GND_net), .O(n28345));   // verilog/coms.v(127[12] 300[6])
    defparam i14834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5299));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15102_3_lut (.I0(current[11]), .I1(data_adj_5377[11]), .I2(n44589), 
            .I3(GND_net), .O(n28613));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15103_3_lut (.I0(current[10]), .I1(data_adj_5377[10]), .I2(n44589), 
            .I3(GND_net), .O(n28614));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15104_3_lut (.I0(current[9]), .I1(data_adj_5377[9]), .I2(n44589), 
            .I3(GND_net), .O(n28615));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14835_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n23568), .I3(GND_net), .O(n28346));   // verilog/coms.v(127[12] 300[6])
    defparam i14835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14836_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n23568), .I3(GND_net), .O(n28347));   // verilog/coms.v(127[12] 300[6])
    defparam i14836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14837_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n23568), .I3(GND_net), .O(n28348));   // verilog/coms.v(127[12] 300[6])
    defparam i14837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14838_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n23568), .I3(GND_net), .O(n28349));   // verilog/coms.v(127[12] 300[6])
    defparam i14838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15105_3_lut (.I0(current[8]), .I1(data_adj_5377[8]), .I2(n44589), 
            .I3(GND_net), .O(n28616));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14839_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n23568), .I3(GND_net), .O(n28350));   // verilog/coms.v(127[12] 300[6])
    defparam i14839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15106_3_lut (.I0(current[7]), .I1(data_adj_5377[7]), .I2(n44589), 
            .I3(GND_net), .O(n28617));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14840_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n23568), .I3(GND_net), .O(n28351));   // verilog/coms.v(127[12] 300[6])
    defparam i14840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14841_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n23568), 
            .I3(GND_net), .O(n28352));   // verilog/coms.v(127[12] 300[6])
    defparam i14841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14842_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n23568), 
            .I3(GND_net), .O(n28353));   // verilog/coms.v(127[12] 300[6])
    defparam i14842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14843_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n23568), 
            .I3(GND_net), .O(n28354));   // verilog/coms.v(127[12] 300[6])
    defparam i14843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14844_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n23568), 
            .I3(GND_net), .O(n28355));   // verilog/coms.v(127[12] 300[6])
    defparam i14844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15107_3_lut (.I0(current[6]), .I1(data_adj_5377[6]), .I2(n44589), 
            .I3(GND_net), .O(n28618));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14845_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n23568), 
            .I3(GND_net), .O(n28356));   // verilog/coms.v(127[12] 300[6])
    defparam i14845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14846_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n23568), 
            .I3(GND_net), .O(n28357));   // verilog/coms.v(127[12] 300[6])
    defparam i14846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14847_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n23568), 
            .I3(GND_net), .O(n28358));   // verilog/coms.v(127[12] 300[6])
    defparam i14847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32712_3_lut (.I0(n2622), .I1(n2689), .I2(n2643), .I3(GND_net), 
            .O(n2721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14848_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n23568), 
            .I3(GND_net), .O(n28359));   // verilog/coms.v(127[12] 300[6])
    defparam i14848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14849_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28360));   // verilog/coms.v(127[12] 300[6])
    defparam i14849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32713_3_lut (.I0(n2721), .I1(n2788), .I2(n2742), .I3(GND_net), 
            .O(n2820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14850_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28361));   // verilog/coms.v(127[12] 300[6])
    defparam i14850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15108_3_lut (.I0(current[5]), .I1(data_adj_5377[5]), .I2(n44589), 
            .I3(GND_net), .O(n28619));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14716_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n23568), .I3(GND_net), .O(n28227));   // verilog/coms.v(127[12] 300[6])
    defparam i14716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14717_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n23568), .I3(GND_net), .O(n28228));   // verilog/coms.v(127[12] 300[6])
    defparam i14717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14851_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n45261), .I3(GND_net), 
            .O(n28362));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i14851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14861_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5223), 
            .I3(n26339), .O(n28372));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14861_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14862_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28373));   // verilog/coms.v(127[12] 300[6])
    defparam i14862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14718_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n23568), .I3(GND_net), .O(n28229));   // verilog/coms.v(127[12] 300[6])
    defparam i14718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2188_add_4_9_lut (.I0(n47182), .I1(n33855), .I2(dti_counter[7]), 
            .I3(n38922), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i15109_3_lut (.I0(current[4]), .I1(data_adj_5377[4]), .I2(n44589), 
            .I3(GND_net), .O(n28620));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 dti_counter_2188_add_4_8_lut (.I0(n47183), .I1(n33855), .I2(dti_counter[6]), 
            .I3(n38921), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_8 (.CI(n38921), .I0(n33855), .I1(dti_counter[6]), 
            .CO(n38922));
    SB_LUT4 dti_counter_2188_add_4_7_lut (.I0(n47184), .I1(n33855), .I2(dti_counter[5]), 
            .I3(n38920), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_7 (.CI(n38920), .I0(n33855), .I1(dti_counter[5]), 
            .CO(n38921));
    SB_LUT4 dti_counter_2188_add_4_6_lut (.I0(n47185), .I1(n33855), .I2(dti_counter[4]), 
            .I3(n38919), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_6 (.CI(n38919), .I0(n33855), .I1(dti_counter[4]), 
            .CO(n38920));
    SB_LUT4 dti_counter_2188_add_4_5_lut (.I0(n47186), .I1(n33855), .I2(dti_counter[3]), 
            .I3(n38918), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_5 (.CI(n38918), .I0(n33855), .I1(dti_counter[3]), 
            .CO(n38919));
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n38459), .I0(n1029), 
            .I1(GND_net), .CO(n38460));
    SB_LUT4 dti_counter_2188_add_4_4_lut (.I0(n47187), .I1(n33855), .I2(dti_counter[2]), 
            .I3(n38917), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_4 (.CI(n38917), .I0(n33855), .I1(dti_counter[2]), 
            .CO(n38918));
    SB_LUT4 dti_counter_2188_add_4_3_lut (.I0(n47188), .I1(n33855), .I2(dti_counter[1]), 
            .I3(n38916), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2188_add_4_3 (.CI(n38916), .I0(n33855), .I1(dti_counter[1]), 
            .CO(n38917));
    SB_LUT4 dti_counter_2188_add_4_2_lut (.I0(n47224), .I1(n1964), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_2188_add_4_2 (.CI(VCC_net), .I0(n1964), .I1(dti_counter[0]), 
            .CO(n38916));
    SB_LUT4 add_2693_25_lut (.I0(n48384), .I1(n2_adj_5276), .I2(n1059), 
            .I3(n38915), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2693_24_lut (.I0(n48371), .I1(n2_adj_5276), .I2(n1158), 
            .I3(n38914), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_24 (.CI(n38914), .I0(n2_adj_5276), .I1(n1158), .CO(n38915));
    SB_LUT4 add_2693_23_lut (.I0(n48357), .I1(n2_adj_5276), .I2(n1257), 
            .I3(n38913), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_23 (.CI(n38913), .I0(n2_adj_5276), .I1(n1257), .CO(n38914));
    SB_LUT4 i15110_3_lut (.I0(current[3]), .I1(data_adj_5377[3]), .I2(n44589), 
            .I3(GND_net), .O(n28621));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_22_lut (.I0(n48330), .I1(n2_adj_5276), .I2(n1356), 
            .I3(n38912), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_224_6 (.CI(n38125), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n38126));
    SB_CARRY add_2693_22 (.CI(n38912), .I0(n2_adj_5276), .I1(n1356), .CO(n38913));
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_21_lut (.I0(n48326), .I1(n2_adj_5276), .I2(n1455), 
            .I3(n38911), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_21 (.CI(n38911), .I0(n2_adj_5276), .I1(n1455), .CO(n38912));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_145_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n38092), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n38099), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n38124), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2693_20_lut (.I0(n48309), .I1(n2_adj_5276), .I2(n1554), 
            .I3(n38910), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_20 (.CI(n38910), .I0(n2_adj_5276), .I1(n1554), .CO(n38911));
    SB_LUT4 add_2693_19_lut (.I0(n48291), .I1(n2_adj_5276), .I2(n1653), 
            .I3(n38909), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n38458), .O(n1097_adj_5257)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_5 (.CI(n38124), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n38125));
    SB_CARRY add_2693_19 (.CI(n38909), .I0(n2_adj_5276), .I1(n1653), .CO(n38910));
    SB_LUT4 add_2693_18_lut (.I0(n48271), .I1(n2_adj_5276), .I2(n1752), 
            .I3(n38908), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_18 (.CI(n38908), .I0(n2_adj_5276), .I1(n1752), .CO(n38909));
    SB_LUT4 add_2693_17_lut (.I0(n48248), .I1(n2_adj_5276), .I2(n1851), 
            .I3(n38907), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_17 (.CI(n38907), .I0(n2_adj_5276), .I1(n1851), .CO(n38908));
    SB_LUT4 add_2693_16_lut (.I0(n48230), .I1(n2_adj_5276), .I2(n1950), 
            .I3(n38906), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_16 (.CI(n38906), .I0(n2_adj_5276), .I1(n1950), .CO(n38907));
    SB_LUT4 pwm_setpoint_23__I_0_i1_3_lut (.I0(duty[0]), .I1(pwm_setpoint_23__N_191[0]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2693_15_lut (.I0(n48209), .I1(n2_adj_5276), .I2(n2049), 
            .I3(n38905), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_15 (.CI(n38905), .I0(n2_adj_5276), .I1(n2049), .CO(n38906));
    SB_LUT4 i14866_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28377));   // verilog/coms.v(127[12] 300[6])
    defparam i14866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1660 (.I0(n2826), .I1(n2822), .I2(n2827), .I3(n2825), 
            .O(n45960));
    defparam i1_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1661 (.I0(n45960), .I1(n2821), .I2(n2828), .I3(GND_net), 
            .O(n45962));
    defparam i1_3_lut_adj_1661.LUT_INIT = 16'hfefe;
    SB_LUT4 i15111_3_lut (.I0(current[2]), .I1(data_adj_5377[2]), .I2(n44589), 
            .I3(GND_net), .O(n28622));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15111_3_lut.LUT_INIT = 16'hacac;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_224_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n38123), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2693_14_lut (.I0(n48186), .I1(n2_adj_5276), .I2(n2148), 
            .I3(n38904), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_14 (.CI(n38904), .I0(n2_adj_5276), .I1(n2148), .CO(n38905));
    SB_LUT4 add_2693_13_lut (.I0(n48746), .I1(n2_adj_5276), .I2(n2247), 
            .I3(n38903), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_13 (.CI(n38903), .I0(n2_adj_5276), .I1(n2247), .CO(n38904));
    SB_LUT4 i14867_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28378));   // verilog/coms.v(127[12] 300[6])
    defparam i14867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14868_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28379));   // verilog/coms.v(127[12] 300[6])
    defparam i14868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14869_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28380));   // verilog/coms.v(127[12] 300[6])
    defparam i14869_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i15112_3_lut (.I0(current[1]), .I1(data_adj_5377[1]), .I2(n44589), 
            .I3(GND_net), .O(n28623));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14870_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28381));   // verilog/coms.v(127[12] 300[6])
    defparam i14870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14871_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28382));   // verilog/coms.v(127[12] 300[6])
    defparam i14871_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n38458), .I0(n1030), 
            .I1(GND_net), .CO(n38459));
    SB_LUT4 i14872_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28383));   // verilog/coms.v(127[12] 300[6])
    defparam i14872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2693_12_lut (.I0(n48687), .I1(n2_adj_5276), .I2(n2346), 
            .I3(n38902), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_12 (.CI(n38902), .I0(n2_adj_5276), .I1(n2346), .CO(n38903));
    SB_LUT4 add_2693_11_lut (.I0(n48719), .I1(n2_adj_5276), .I2(n2445), 
            .I3(n38901), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_11 (.CI(n38901), .I0(n2_adj_5276), .I1(n2445), .CO(n38902));
    SB_LUT4 add_2693_10_lut (.I0(n48659), .I1(n2_adj_5276), .I2(n2544), 
            .I3(n38900), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_10 (.CI(n38900), .I0(n2_adj_5276), .I1(n2544), .CO(n38901));
    SB_LUT4 add_2693_9_lut (.I0(n48634), .I1(n2_adj_5276), .I2(n2643), 
            .I3(n38899), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_9 (.CI(n38899), .I0(n2_adj_5276), .I1(n2643), .CO(n38900));
    SB_LUT4 add_2693_8_lut (.I0(n48601), .I1(n2_adj_5276), .I2(n2742), 
            .I3(n38898), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_8 (.CI(n38898), .I0(n2_adj_5276), .I1(n2742), .CO(n38899));
    SB_LUT4 add_2693_7_lut (.I0(n48571), .I1(n2_adj_5276), .I2(n2841), 
            .I3(n38897), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_7 (.CI(n38897), .I0(n2_adj_5276), .I1(n2841), .CO(n38898));
    SB_LUT4 add_2693_6_lut (.I0(n48540), .I1(n2_adj_5276), .I2(n2940), 
            .I3(n38896), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n38457), .O(n1098_adj_5258)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14873_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n27595), 
            .I3(GND_net), .O(n28384));   // verilog/coms.v(127[12] 300[6])
    defparam i14873_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2693_6 (.CI(n38896), .I0(n2_adj_5276), .I1(n2940), .CO(n38897));
    SB_LUT4 i14874_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n27595), 
            .I3(GND_net), .O(n28385));   // verilog/coms.v(127[12] 300[6])
    defparam i14874_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n38457), .I0(n1031), 
            .I1(VCC_net), .CO(n38458));
    SB_LUT4 add_2693_5_lut (.I0(n48507), .I1(n2_adj_5276), .I2(n3039), 
            .I3(n38895), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14875_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n27595), 
            .I3(GND_net), .O(n28386));   // verilog/coms.v(127[12] 300[6])
    defparam i14875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14876_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n27595), 
            .I3(GND_net), .O(n28387));   // verilog/coms.v(127[12] 300[6])
    defparam i14876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n2819), .I1(n2820), .I2(n2824), .I3(n2823), 
            .O(n45964));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i14877_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n27595), 
            .I3(GND_net), .O(n28388));   // verilog/coms.v(127[12] 300[6])
    defparam i14877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21135_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n34644));
    defparam i21135_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n38456), .O(n1099_adj_5259)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2693_5 (.CI(n38895), .I0(n2_adj_5276), .I1(n3039), .CO(n38896));
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n38456), .I0(n1032), 
            .I1(GND_net), .CO(n38457));
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n38455), .O(n1100_adj_5260)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14878_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n27595), 
            .I3(GND_net), .O(n28389));   // verilog/coms.v(127[12] 300[6])
    defparam i14878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2693_4_lut (.I0(n48475), .I1(n2_adj_5276), .I2(n3138), 
            .I3(n38894), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_4 (.CI(n38894), .I0(n2_adj_5276), .I1(n3138), .CO(n38895));
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n38455), .I0(n1033), 
            .I1(VCC_net), .CO(n38456));
    SB_LUT4 i14879_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n27595), 
            .I3(GND_net), .O(n28390));   // verilog/coms.v(127[12] 300[6])
    defparam i14879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14880_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n27595), 
            .I3(GND_net), .O(n28391));   // verilog/coms.v(127[12] 300[6])
    defparam i14880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14881_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n27595), 
            .I3(GND_net), .O(n28392));   // verilog/coms.v(127[12] 300[6])
    defparam i14881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14882_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n27595), 
            .I3(GND_net), .O(n28393));   // verilog/coms.v(127[12] 300[6])
    defparam i14882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2693_3_lut (.I0(n48440), .I1(n2_adj_5276), .I2(n3237), 
            .I3(n38893), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14883_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n27595), 
            .I3(GND_net), .O(n28394));   // verilog/coms.v(127[12] 300[6])
    defparam i14883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14884_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n27595), 
            .I3(GND_net), .O(n28395));   // verilog/coms.v(127[12] 300[6])
    defparam i14884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14885_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n27595), 
            .I3(GND_net), .O(n28396));   // verilog/coms.v(127[12] 300[6])
    defparam i14885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1663 (.I0(n2817), .I1(n2818), .I2(n45964), .I3(n45962), 
            .O(n45970));
    defparam i1_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_CARRY add_2693_3 (.CI(n38893), .I0(n2_adj_5276), .I1(n3237), .CO(n38894));
    SB_LUT4 i1_4_lut_adj_1664 (.I0(n2829), .I1(n45970), .I2(n34644), .I3(n2830), 
            .O(n45972));
    defparam i1_4_lut_adj_1664.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1665 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n45972), 
            .O(n45978));
    defparam i1_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_10_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2693_2_lut (.I0(n48394), .I1(n2_adj_5276), .I2(n34750), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14886_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n27595), 
            .I3(GND_net), .O(n28397));   // verilog/coms.v(127[12] 300[6])
    defparam i14886_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2693_2 (.CI(VCC_net), .I0(n2_adj_5276), .I1(n34750), 
            .CO(n38893));
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(GND_net), .I1(n3204), 
            .I2(VCC_net), .I3(n38892), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n38891), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n38891), .I0(n3205), 
            .I1(VCC_net), .CO(n38892));
    SB_LUT4 i1_4_lut_adj_1666 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n45978), 
            .O(n45984));
    defparam i1_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n38890), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n38890), .I0(n3206), 
            .I1(VCC_net), .CO(n38891));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n38889), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n38889), .I0(n3207), 
            .I1(VCC_net), .CO(n38890));
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n38888), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n38888), .I0(n3208), 
            .I1(VCC_net), .CO(n38889));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n38887), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14887_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n27595), 
            .I3(GND_net), .O(n28398));   // verilog/coms.v(127[12] 300[6])
    defparam i14887_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n38887), .I0(n3209), 
            .I1(VCC_net), .CO(n38888));
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n38886), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n38886), .I0(n3210), 
            .I1(VCC_net), .CO(n38887));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n38885), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n38885), .I0(n3211), 
            .I1(VCC_net), .CO(n38886));
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101_adj_5261)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n38455));
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n38884), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14888_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n27595), 
            .I3(GND_net), .O(n28399));   // verilog/coms.v(127[12] 300[6])
    defparam i14888_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n38884), .I0(n3212), 
            .I1(VCC_net), .CO(n38885));
    SB_LUT4 i14889_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n27595), 
            .I3(GND_net), .O(n28400));   // verilog/coms.v(127[12] 300[6])
    defparam i14889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n38883), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n38883), .I0(n3213), 
            .I1(VCC_net), .CO(n38884));
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n38882), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n38882), .I0(n3214), 
            .I1(VCC_net), .CO(n38883));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n38881), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15118_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n42822), 
            .I3(GND_net), .O(n28629));   // verilog/coms.v(127[12] 300[6])
    defparam i15118_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n38881), .I0(n3215), 
            .I1(VCC_net), .CO(n38882));
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n38880), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n38880), .I0(n3216), 
            .I1(VCC_net), .CO(n38881));
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n38879), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n38879), .I0(n3217), 
            .I1(VCC_net), .CO(n38880));
    SB_LUT4 i14890_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n27595), 
            .I3(GND_net), .O(n28401));   // verilog/coms.v(127[12] 300[6])
    defparam i14890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_5245), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n38878), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n38878), .I0(n3218), 
            .I1(VCC_net), .CO(n38879));
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n38454), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n38877), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n38877), .I0(n3219), 
            .I1(VCC_net), .CO(n38878));
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n38453), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n38876), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14891_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n27595), 
            .I3(GND_net), .O(n28402));   // verilog/coms.v(127[12] 300[6])
    defparam i14891_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n38876), .I0(n3220), 
            .I1(VCC_net), .CO(n38877));
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n38453), .I0(n928), 
            .I1(VCC_net), .CO(n38454));
    SB_LUT4 i14892_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n27595), 
            .I3(GND_net), .O(n28403));   // verilog/coms.v(127[12] 300[6])
    defparam i14892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n38875), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n38875), .I0(n3221), 
            .I1(VCC_net), .CO(n38876));
    SB_LUT4 i14893_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n27595), 
            .I3(GND_net), .O(n28404));   // verilog/coms.v(127[12] 300[6])
    defparam i14893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n38874), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n38452), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n38874), .I0(n3222), 
            .I1(VCC_net), .CO(n38875));
    SB_LUT4 i14894_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n27595), 
            .I3(GND_net), .O(n28405));   // verilog/coms.v(127[12] 300[6])
    defparam i14894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n38873), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33494_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n45984), 
            .O(n2841));
    defparam i33494_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n38873), .I0(n3223), 
            .I1(VCC_net), .CO(n38874));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n38872), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n38872), .I0(n3224), 
            .I1(VCC_net), .CO(n38873));
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n38871), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n38871), .I0(n3225), 
            .I1(VCC_net), .CO(n38872));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n38870), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n38870), .I0(n3226), 
            .I1(VCC_net), .CO(n38871));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n38869), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n38869), .I0(n3227), 
            .I1(VCC_net), .CO(n38870));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n38868), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n38868), .I0(n3228), 
            .I1(VCC_net), .CO(n38869));
    SB_LUT4 i15119_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n42822), 
            .I3(GND_net), .O(n28630));   // verilog/coms.v(127[12] 300[6])
    defparam i15119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n38867), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n38867), .I0(n3229), 
            .I1(GND_net), .CO(n38868));
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n38866), .O(n47200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n38866), .I0(n3230), 
            .I1(GND_net), .CO(n38867));
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n38865), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n38865), .I0(n3231), 
            .I1(VCC_net), .CO(n38866));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n38864), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n38864), .I0(n3232), 
            .I1(GND_net), .CO(n38865));
    SB_LUT4 i14895_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n27595), 
            .I3(GND_net), .O(n28406));   // verilog/coms.v(127[12] 300[6])
    defparam i14895_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n38452), .I0(n929), 
            .I1(GND_net), .CO(n38453));
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n38863), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n38863), .I0(n3233), 
            .I1(VCC_net), .CO(n38864));
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n38451), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14896_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n27595), 
            .I3(GND_net), .O(n28407));   // verilog/coms.v(127[12] 300[6])
    defparam i14896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14897_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28408));   // verilog/coms.v(127[12] 300[6])
    defparam i14897_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n38451), .I0(n930), 
            .I1(GND_net), .CO(n38452));
    SB_LUT4 i1_4_lut_adj_1667 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5267));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'h7bde;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n38862), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n38862), .I0(n957), 
            .I1(GND_net), .CO(n38863));
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n38862));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n48475), .I1(n3105), 
            .I2(VCC_net), .I3(n38861), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n38860), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n38860), .I0(n3106), 
            .I1(VCC_net), .CO(n38861));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n38859), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n38859), .I0(n3107), 
            .I1(VCC_net), .CO(n38860));
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n38858), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n38858), .I0(n3108), 
            .I1(VCC_net), .CO(n38859));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n38857), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n38857), .I0(n3109), 
            .I1(VCC_net), .CO(n38858));
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n38856), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n38856), .I0(n3110), 
            .I1(VCC_net), .CO(n38857));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n38855), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n38450), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n38450), .I0(n931), 
            .I1(VCC_net), .CO(n38451));
    SB_LUT4 i14898_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28409));   // verilog/coms.v(127[12] 300[6])
    defparam i14898_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n38855), .I0(n3111), 
            .I1(VCC_net), .CO(n38856));
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n38854), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n38854), .I0(n3112), 
            .I1(VCC_net), .CO(n38855));
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n38449), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n38853), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n38853), .I0(n3113), 
            .I1(VCC_net), .CO(n38854));
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n38852), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n38852), .I0(n3114), 
            .I1(VCC_net), .CO(n38853));
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14899_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28410));   // verilog/coms.v(127[12] 300[6])
    defparam i14899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14900_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28411));   // verilog/coms.v(127[12] 300[6])
    defparam i14900_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_4 (.CI(n38123), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n38124));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n38851), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n38851), .I0(n3115), 
            .I1(VCC_net), .CO(n38852));
    SB_LUT4 i1_4_lut_adj_1668 (.I0(n5_adj_5274), .I1(n122), .I2(n3813), 
            .I3(n63), .O(n6_adj_5273));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'heaaa;
    SB_LUT4 unary_minus_10_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5165));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1669 (.I0(n49229), .I1(n6_adj_5273), .I2(\FRAME_MATCHER.i_31__N_2626 ), 
            .I3(n4452), .O(n8_adj_5206));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1669.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1670 (.I0(n122), .I1(n8_adj_5206), .I2(\FRAME_MATCHER.i_31__N_2622 ), 
            .I3(n7_adj_5175), .O(n49000));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1670.LUT_INIT = 16'hfefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n38850), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n38850), .I0(n3116), 
            .I1(VCC_net), .CO(n38851));
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n38849), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n38122), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n38449), .I0(n932), 
            .I1(GND_net), .CO(n38450));
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n38849), .I0(n3117), 
            .I1(VCC_net), .CO(n38850));
    SB_LUT4 unary_minus_10_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n38848), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n38848), .I0(n3118), 
            .I1(VCC_net), .CO(n38849));
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_11 (.CI(n38099), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n38100));
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n38847), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_3 (.CI(n38122), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n38123));
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n38847), .I0(n3119), 
            .I1(VCC_net), .CO(n38848));
    SB_LUT4 i14901_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28412));   // verilog/coms.v(127[12] 300[6])
    defparam i14901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14902_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28413));   // verilog/coms.v(127[12] 300[6])
    defparam i14902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15121_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n42822), 
            .I3(GND_net), .O(n28632));   // verilog/coms.v(127[12] 300[6])
    defparam i15121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n38846), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15122_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n42822), 
            .I3(GND_net), .O(n28633));   // verilog/coms.v(127[12] 300[6])
    defparam i15122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_279), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14903_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28414));   // verilog/coms.v(127[12] 300[6])
    defparam i14903_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_279), 
            .CO(n38122));
    SB_LUT4 add_145_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n38121), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n38846), .I0(n3120), 
            .I1(VCC_net), .CO(n38847));
    SB_LUT4 i14904_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28415));   // verilog/coms.v(127[12] 300[6])
    defparam i14904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n38845), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n38845), .I0(n3121), 
            .I1(VCC_net), .CO(n38846));
    SB_LUT4 i15123_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n42822), 
            .I3(GND_net), .O(n28634));   // verilog/coms.v(127[12] 300[6])
    defparam i15123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14905_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n27595), 
            .I3(GND_net), .O(n28416));   // verilog/coms.v(127[12] 300[6])
    defparam i14905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n38844), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n38844), .I0(n3122), 
            .I1(VCC_net), .CO(n38845));
    SB_LUT4 i15124_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n27595), 
            .I3(GND_net), .O(n28635));   // verilog/coms.v(127[12] 300[6])
    defparam i15124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n38843), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_adj_1671 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5205));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i2_2_lut_adj_1671.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n38843), .I0(n3123), 
            .I1(VCC_net), .CO(n38844));
    SB_LUT4 i14908_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n45341), .I3(GND_net), 
            .O(n28419));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15125_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n42822), 
            .I3(GND_net), .O(n28636));   // verilog/coms.v(127[12] 300[6])
    defparam i15125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14909_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n27595), .I3(GND_net), .O(n28420));   // verilog/coms.v(127[12] 300[6])
    defparam i14909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14910_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28421));   // verilog/coms.v(127[12] 300[6])
    defparam i14910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n38842), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n38842), .I0(n3124), 
            .I1(VCC_net), .CO(n38843));
    SB_CARRY add_145_4 (.CI(n38092), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n38093));
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n38841), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n38841), .I0(n3125), 
            .I1(VCC_net), .CO(n38842));
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n38840), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n38840), .I0(n3126), 
            .I1(VCC_net), .CO(n38841));
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n38839), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n38839), .I0(n3127), 
            .I1(VCC_net), .CO(n38840));
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n38448), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n38838), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n38448), .I0(n933), 
            .I1(VCC_net), .CO(n38449));
    SB_LUT4 add_145_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n38098), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n38838), .I0(n3128), 
            .I1(VCC_net), .CO(n38839));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n38837), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n38837), .I0(n3129), 
            .I1(GND_net), .CO(n38838));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n38836), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14911_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28422));   // verilog/coms.v(127[12] 300[6])
    defparam i14911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15126_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n42822), 
            .I3(GND_net), .O(n28637));   // verilog/coms.v(127[12] 300[6])
    defparam i15126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14912_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28423));   // verilog/coms.v(127[12] 300[6])
    defparam i14912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14913_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28424));   // verilog/coms.v(127[12] 300[6])
    defparam i14913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14914_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28425));   // verilog/coms.v(127[12] 300[6])
    defparam i14914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n38120), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n38836), .I0(n3130), 
            .I1(GND_net), .CO(n38837));
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n38835), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n38835), .I0(n3131), 
            .I1(VCC_net), .CO(n38836));
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n38834), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n38834), .I0(n3132), 
            .I1(GND_net), .CO(n38835));
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n38833), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n38833), .I0(n3133), 
            .I1(VCC_net), .CO(n38834));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n38833));
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(n48507), .I1(n3006), 
            .I2(VCC_net), .I3(n38832), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n38448));
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n38831), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n38831), .I0(n3007), 
            .I1(VCC_net), .CO(n38832));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n38830), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n38830), .I0(n3008), 
            .I1(VCC_net), .CO(n38831));
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n38829), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n38829), .I0(n3009), 
            .I1(VCC_net), .CO(n38830));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n38828), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n38828), .I0(n3010), 
            .I1(VCC_net), .CO(n38829));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n38827), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n38827), .I0(n3011), 
            .I1(VCC_net), .CO(n38828));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n38826), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n38826), .I0(n3012), 
            .I1(VCC_net), .CO(n38827));
    SB_LUT4 i6_4_lut_adj_1672 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5204));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i6_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n38825), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33264_4_lut (.I0(n43818), .I1(n1323), .I2(n1324), .I3(n45644), 
            .O(n1356));
    defparam i33264_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n1329), .I1(n34608), .I2(n1330), .I3(n1331), 
            .O(n43818));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n45644));
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i21100_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n34608));
    defparam i21100_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33279_4_lut (.I0(n1225), .I1(n1224), .I2(n43821), .I3(n45686), 
            .O(n1257));
    defparam i33279_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(n1229), .I1(n34610), .I2(n1230), .I3(n1231), 
            .O(n43821));
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n38825), .I0(n3013), 
            .I1(VCC_net), .CO(n38826));
    SB_LUT4 i15127_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n42822), 
            .I3(GND_net), .O(n28638));   // verilog/coms.v(127[12] 300[6])
    defparam i15127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14915_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28426));   // verilog/coms.v(127[12] 300[6])
    defparam i14915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14916_4_lut (.I0(CS_MISO_c), .I1(data_adj_5377[0]), .I2(n11_adj_5231), 
            .I3(state_7__N_4293), .O(n28427));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14916_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14917_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28428));   // verilog/coms.v(127[12] 300[6])
    defparam i14917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14918_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n27595), .I3(GND_net), .O(n28429));   // verilog/coms.v(127[12] 300[6])
    defparam i14918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14919_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n27595), .I3(GND_net), .O(n28430));   // verilog/coms.v(127[12] 300[6])
    defparam i14919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n38824), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n38824), .I0(n3014), 
            .I1(VCC_net), .CO(n38825));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n38823), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n38823), .I0(n3015), 
            .I1(VCC_net), .CO(n38824));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n38822), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n38822), .I0(n3016), 
            .I1(VCC_net), .CO(n38823));
    SB_LUT4 i14920_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n27595), .I3(GND_net), .O(n28431));   // verilog/coms.v(127[12] 300[6])
    defparam i14920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n38821), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n38447), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14921_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n27595), .I3(GND_net), .O(n28432));   // verilog/coms.v(127[12] 300[6])
    defparam i14921_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n38821), .I0(n3017), 
            .I1(VCC_net), .CO(n38822));
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14922_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n27595), .I3(GND_net), .O(n28433));   // verilog/coms.v(127[12] 300[6])
    defparam i14922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14926_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n27595), .I3(GND_net), .O(n28437));   // verilog/coms.v(127[12] 300[6])
    defparam i14926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n2723), .I1(n2721), .I2(n2726), .I3(n2728), 
            .O(n45366));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1677 (.I0(n2725), .I1(n2720), .I2(n2727), .I3(GND_net), 
            .O(n45364));
    defparam i1_3_lut_adj_1677.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1678 (.I0(n45366), .I1(n2722), .I2(n2724), .I3(GND_net), 
            .O(n45368));
    defparam i1_3_lut_adj_1678.LUT_INIT = 16'hfefe;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n38446), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n38446), .I0(n829), 
            .I1(GND_net), .CO(n38447));
    SB_CARRY add_145_32 (.CI(n38120), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n38121));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n38820), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n38820), .I0(n3018), 
            .I1(VCC_net), .CO(n38821));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n38819), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n38119), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21137_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n34646));
    defparam i21137_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i14927_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n27595), .I3(GND_net), .O(n28438));   // verilog/coms.v(127[12] 300[6])
    defparam i14927_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14934_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n42836), .I3(GND_net), .O(n28445));   // verilog/coms.v(127[12] 300[6])
    defparam i14934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1679 (.I0(n2718), .I1(n2719), .I2(n45368), .I3(n45364), 
            .O(n45374));
    defparam i1_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14935_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n42836), .I3(GND_net), .O(n28446));   // verilog/coms.v(127[12] 300[6])
    defparam i14935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n2729), .I1(n45374), .I2(n34646), .I3(n2730), 
            .O(n45376));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'heccc;
    SB_LUT4 i14936_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n42836), .I3(GND_net), .O(n28447));   // verilog/coms.v(127[12] 300[6])
    defparam i14936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n2715), .I1(n2716), .I2(n45376), .I3(n2717), 
            .O(n45382));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i14937_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n42836), .I3(GND_net), .O(n28448));   // verilog/coms.v(127[12] 300[6])
    defparam i14937_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n38819), .I0(n3019), 
            .I1(VCC_net), .CO(n38820));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n38818), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n38818), .I0(n3020), 
            .I1(VCC_net), .CO(n38819));
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n38817), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n38817), .I0(n3021), 
            .I1(VCC_net), .CO(n38818));
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n38816), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n38816), .I0(n3022), 
            .I1(VCC_net), .CO(n38817));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n38815), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n38815), .I0(n3023), 
            .I1(VCC_net), .CO(n38816));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n38814), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n38814), .I0(n3024), 
            .I1(VCC_net), .CO(n38815));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n38813), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n38813), .I0(n3025), 
            .I1(VCC_net), .CO(n38814));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n38812), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n38812), .I0(n3026), 
            .I1(VCC_net), .CO(n38813));
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n38811), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n38811), .I0(n3027), 
            .I1(VCC_net), .CO(n38812));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n38810), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n38445), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n38810), .I0(n3028), 
            .I1(VCC_net), .CO(n38811));
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14938_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n42836), .I3(GND_net), .O(n28449));   // verilog/coms.v(127[12] 300[6])
    defparam i14938_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n7072), 
            .D(n1105), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n38809), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n38809), .I0(n3029), 
            .I1(GND_net), .CO(n38810));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n38808), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n38808), .I0(n3030), 
            .I1(GND_net), .CO(n38809));
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n38807), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n38807), .I0(n3031), 
            .I1(VCC_net), .CO(n38808));
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n38806), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n38806), .I0(n3032), 
            .I1(GND_net), .CO(n38807));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n38805), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n38805), .I0(n3033), 
            .I1(VCC_net), .CO(n38806));
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n38805));
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n48540), .I1(n2907), 
            .I2(VCC_net), .I3(n38804), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n38803), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n38803), .I0(n2908), 
            .I1(VCC_net), .CO(n38804));
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n38802), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n38802), .I0(n2909), 
            .I1(VCC_net), .CO(n38803));
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n38801), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n38801), .I0(n2910), 
            .I1(VCC_net), .CO(n38802));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n38800), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n38800), .I0(n2911), 
            .I1(VCC_net), .CO(n38801));
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n38799), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n38799), .I0(n2912), 
            .I1(VCC_net), .CO(n38800));
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n38798), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n38798), .I0(n2913), 
            .I1(VCC_net), .CO(n38799));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n38797), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n38797), .I0(n2914), 
            .I1(VCC_net), .CO(n38798));
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n38796), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n38796), .I0(n2915), 
            .I1(VCC_net), .CO(n38797));
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n38795), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n38795), .I0(n2916), 
            .I1(VCC_net), .CO(n38796));
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n45382), 
            .O(n45388));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n38794), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n38794), .I0(n2917), 
            .I1(VCC_net), .CO(n38795));
    SB_LUT4 i14939_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n42836), .I3(GND_net), .O(n28450));   // verilog/coms.v(127[12] 300[6])
    defparam i14939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n38793), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n7072), 
            .D(n1104), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n38793), .I0(n2918), 
            .I1(VCC_net), .CO(n38794));
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n38792), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n38792), .I0(n2919), 
            .I1(VCC_net), .CO(n38793));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n38791), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33524_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n45388), 
            .O(n2742));
    defparam i33524_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n38791), .I0(n2920), 
            .I1(VCC_net), .CO(n38792));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n38790), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n38790), .I0(n2921), 
            .I1(VCC_net), .CO(n38791));
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n38445), .I0(n830), 
            .I1(GND_net), .CO(n38446));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n38789), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n38789), .I0(n2922), 
            .I1(VCC_net), .CO(n38790));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n38444), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n7072), 
            .D(n1103), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n38444), .I0(n831), 
            .I1(VCC_net), .CO(n38445));
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n38443), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n7072), 
            .D(n1102), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n38443), .I0(n832), 
            .I1(GND_net), .CO(n38444));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n38442), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14940_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n42836), .I3(GND_net), .O(n28451));   // verilog/coms.v(127[12] 300[6])
    defparam i14940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1683 (.I0(dti_counter[0]), .I1(n14_adj_5204), .I2(n10_adj_5205), 
            .I3(dti_counter[3]), .O(n23755));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i7_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n38788), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14941_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n42836), .I3(GND_net), .O(n28452));   // verilog/coms.v(127[12] 300[6])
    defparam i14941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5246), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n38788), .I0(n2923), 
            .I1(VCC_net), .CO(n38789));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n38787), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n42022));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n42634));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n38787), .I0(n2924), 
            .I1(VCC_net), .CO(n38788));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n38786), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n38786), .I0(n2925), 
            .I1(VCC_net), .CO(n38787));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n38785), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n38785), .I0(n2926), 
            .I1(VCC_net), .CO(n38786));
    SB_CARRY add_145_31 (.CI(n38119), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n38120));
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n38784), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n38784), .I0(n2927), 
            .I1(VCC_net), .CO(n38785));
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n38783), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n38783), .I0(n2928), 
            .I1(VCC_net), .CO(n38784));
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n38442), .I0(n833), 
            .I1(VCC_net), .CO(n38443));
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n38782), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n38782), .I0(n2929), 
            .I1(GND_net), .CO(n38783));
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n38781), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n38781), .I0(n2930), 
            .I1(GND_net), .CO(n38782));
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n38780), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n38780), .I0(n2931), 
            .I1(VCC_net), .CO(n38781));
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n38779), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n38779), .I0(n2932), 
            .I1(GND_net), .CO(n38780));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n38778), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n38778), .I0(n2933), 
            .I1(VCC_net), .CO(n38779));
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n38778));
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n48571), .I1(n2808), 
            .I2(VCC_net), .I3(n38777), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n38776), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n38776), .I0(n2809), 
            .I1(VCC_net), .CO(n38777));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n38775), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n38775), .I0(n2810), 
            .I1(VCC_net), .CO(n38776));
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n38774), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n38774), .I0(n2811), 
            .I1(VCC_net), .CO(n38775));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n38773), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n38773), .I0(n2812), 
            .I1(VCC_net), .CO(n38774));
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n38772), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093_adj_5253), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n38442));
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n38772), .I0(n2813), 
            .I1(VCC_net), .CO(n38773));
    SB_DFF dti_counter_2188__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n38771), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n38771), .I0(n2814), 
            .I1(VCC_net), .CO(n38772));
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n38118), .O(n1080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1722_rep_15_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1722_rep_15_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n38770), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n38770), .I0(n2815), 
            .I1(VCC_net), .CO(n38771));
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098_adj_5258), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY add_145_30 (.CI(n38118), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n38119));
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n38769), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_191[23]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n7072), 
            .D(n1101), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097_adj_5257), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n38769), .I0(n2816), 
            .I1(VCC_net), .CO(n38770));
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n38768), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n38768), .I0(n2817), 
            .I1(VCC_net), .CO(n38769));
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n935), .I1(n1101_adj_5261), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n38767), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n7072), 
            .D(n1090), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n7072), 
            .D(n1100), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n7072), 
            .D(n1099), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i2_3_lut (.I0(duty[1]), .I1(pwm_setpoint_23__N_191[1]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1724_rep_22_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1724_rep_22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100_adj_5260), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i3_3_lut (.I0(duty[2]), .I1(pwm_setpoint_23__N_191[2]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i4_3_lut (.I0(duty[3]), .I1(pwm_setpoint_23__N_191[3]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i5_3_lut (.I0(duty[4]), .I1(pwm_setpoint_23__N_191[4]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1719_rep_23_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1719_rep_23_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1721_rep_20_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1721_rep_20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i6_3_lut (.I0(duty[5]), .I1(pwm_setpoint_23__N_191[5]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i7_3_lut (.I0(duty[6]), .I1(pwm_setpoint_23__N_191[6]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i8_3_lut (.I0(duty[7]), .I1(pwm_setpoint_23__N_191[7]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i9_3_lut (.I0(duty[8]), .I1(pwm_setpoint_23__N_191[8]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1717_rep_21_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1717_rep_21_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i10_3_lut (.I0(duty[9]), .I1(pwm_setpoint_23__N_191[9]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i11_3_lut (.I0(duty[10]), .I1(pwm_setpoint_23__N_191[10]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33027_2_lut (.I0(n23755), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_416));
    defparam i33027_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1684 (.I0(n2621), .I1(n2625), .I2(GND_net), .I3(GND_net), 
            .O(n45868));
    defparam i1_2_lut_adj_1684.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n2624), .I1(n2623), .I2(n2622), .I3(n2628), 
            .O(n45876));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_setpoint_23__I_0_i12_3_lut (.I0(duty[11]), .I1(pwm_setpoint_23__N_191[11]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i13_3_lut (.I0(duty[12]), .I1(pwm_setpoint_23__N_191[12]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i14_3_lut (.I0(duty[13]), .I1(pwm_setpoint_23__N_191[13]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n2627), .I1(n45876), .I2(n45868), .I3(n2626), 
            .O(n45878));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_setpoint_23__I_0_i15_3_lut (.I0(duty[14]), .I1(pwm_setpoint_23__N_191[14]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14719_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n23568), .I3(GND_net), .O(n28230));   // verilog/coms.v(127[12] 300[6])
    defparam i14719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21068_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n34576));
    defparam i21068_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n2618), .I1(n2619), .I2(n45878), .I3(n2620), 
            .O(n45884));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_setpoint_23__I_0_i16_3_lut (.I0(duty[15]), .I1(pwm_setpoint_23__N_191[15]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i17_3_lut (.I0(duty[16]), .I1(pwm_setpoint_23__N_191[16]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i18_3_lut (.I0(duty[17]), .I1(pwm_setpoint_23__N_191[17]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099_adj_5259), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i19_3_lut (.I0(duty[18]), .I1(pwm_setpoint_23__N_191[18]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5247), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n2629), .I1(n34576), .I2(n2630), .I3(n2631), 
            .O(n43941));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n2616), .I1(n2617), .I2(n43941), .I3(n45884), 
            .O(n45890));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_setpoint_23__I_0_i20_3_lut (.I0(duty[19]), .I1(pwm_setpoint_23__N_191[19]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n45890), 
            .O(n45896));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n38767), .I0(n2818), 
            .I1(VCC_net), .CO(n38768));
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33557_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n45896), 
            .O(n2643));
    defparam i33557_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i21_3_lut (.I0(duty[20]), .I1(pwm_setpoint_23__N_191[20]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i22_3_lut (.I0(duty[21]), .I1(pwm_setpoint_23__N_191[21]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n38766), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n38766), .I0(n2819), 
            .I1(VCC_net), .CO(n38767));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n38765), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_setpoint_23__I_0_i23_3_lut (.I0(duty[22]), .I1(pwm_setpoint_23__N_191[22]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n38765), .I0(n2820), 
            .I1(VCC_net), .CO(n38766));
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n7072), 
            .D(n1089), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n38764), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n7072), 
            .D(n1088), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n38764), .I0(n2821), 
            .I1(VCC_net), .CO(n38765));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n38763), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n38763), .I0(n2822), 
            .I1(VCC_net), .CO(n38764));
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n38762), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n38762), .I0(n2823), 
            .I1(VCC_net), .CO(n38763));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n38761), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n38761), .I0(n2824), 
            .I1(VCC_net), .CO(n38762));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n38760), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n38760), .I0(n2825), 
            .I1(VCC_net), .CO(n38761));
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n38759), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n38759), .I0(n2826), 
            .I1(VCC_net), .CO(n38760));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n38758), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n38758), .I0(n2827), 
            .I1(VCC_net), .CO(n38759));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n38757), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n7072), 
            .D(n1098), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n17_adj_5170));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n7072), 
            .D(n1087), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14720_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n23568), .I3(GND_net), .O(n28231));   // verilog/coms.v(127[12] 300[6])
    defparam i14720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14616_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5223), 
            .I3(n26334), .O(n28127));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14616_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14617_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5210), 
            .I3(n26339), .O(n28128));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14617_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14618_4_lut (.I0(state_7__N_4103[3]), .I1(data[1]), .I2(n10_adj_5275), 
            .I3(n26367), .O(n28129));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14618_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n38757), .I0(n2828), 
            .I1(VCC_net), .CO(n38758));
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n38756), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14619_4_lut (.I0(state_7__N_4103[3]), .I1(data[2]), .I2(n4_adj_5232), 
            .I3(n26372), .O(n28130));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14619_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n38756), .I0(n2829), 
            .I1(GND_net), .CO(n38757));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n38755), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n38755), .I0(n2830), 
            .I1(GND_net), .CO(n38756));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n38754), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n38754), .I0(n2831), 
            .I1(VCC_net), .CO(n38755));
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n38753), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n38753), .I0(n2832), 
            .I1(GND_net), .CO(n38754));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n38752), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n38752), .I0(n2833), 
            .I1(VCC_net), .CO(n38753));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n38752));
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n48601), .I1(n2709), 
            .I2(VCC_net), .I3(n38751), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n38750), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n38750), .I0(n2710), 
            .I1(VCC_net), .CO(n38751));
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14620_4_lut (.I0(state_7__N_4103[3]), .I1(data[3]), .I2(n4_adj_5232), 
            .I3(n26367), .O(n28131));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14620_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14621_4_lut (.I0(state_7__N_4103[3]), .I1(data[4]), .I2(n4_adj_5161), 
            .I3(n26372), .O(n28132));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14621_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14622_4_lut (.I0(state_7__N_4103[3]), .I1(data[5]), .I2(n4_adj_5161), 
            .I3(n26367), .O(n28133));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14622_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n38749), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n38749), .I0(n2711), 
            .I1(VCC_net), .CO(n38750));
    SB_LUT4 encoder0_position_31__I_0_i1649_rep_24_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1649_rep_24_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n38748), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n38748), .I0(n2712), 
            .I1(VCC_net), .CO(n38749));
    SB_LUT4 i14623_4_lut (.I0(state_7__N_4103[3]), .I1(data[6]), .I2(n33869), 
            .I3(n26372), .O(n28134));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14623_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n38747), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n38747), .I0(n2713), 
            .I1(VCC_net), .CO(n38748));
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n38746), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n38746), .I0(n2714), 
            .I1(VCC_net), .CO(n38747));
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n38745), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14624_4_lut (.I0(state_7__N_4103[3]), .I1(data[7]), .I2(n33869), 
            .I3(n26367), .O(n28135));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14624_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n38745), .I0(n2715), 
            .I1(VCC_net), .CO(n38746));
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n38744), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n38744), .I0(n2716), 
            .I1(VCC_net), .CO(n38745));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n38743), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n38743), .I0(n2717), 
            .I1(VCC_net), .CO(n38744));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n38742), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n38742), .I0(n2718), 
            .I1(VCC_net), .CO(n38743));
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n38741), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n38741), .I0(n2719), 
            .I1(VCC_net), .CO(n38742));
    SB_LUT4 encoder0_position_31__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n38740), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n38740), .I0(n2720), 
            .I1(VCC_net), .CO(n38741));
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n38739), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n38739), .I0(n2721), 
            .I1(VCC_net), .CO(n38740));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n38738), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n38738), .I0(n2722), 
            .I1(VCC_net), .CO(n38739));
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n38737), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n38737), .I0(n2723), 
            .I1(VCC_net), .CO(n38738));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n38736), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n38736), .I0(n2724), 
            .I1(VCC_net), .CO(n38737));
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n38735), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5362_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_389));
    defparam i5362_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n38735), .I0(n2725), 
            .I1(VCC_net), .CO(n38736));
    SB_LUT4 i14626_4_lut (.I0(n43584), .I1(state[1]), .I2(state_3__N_528[1]), 
            .I3(n27713), .O(n28137));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14626_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i5364_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_398));
    defparam i5364_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n38734), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n38734), .I0(n2726), 
            .I1(VCC_net), .CO(n38735));
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n38733), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n38733), .I0(n2727), 
            .I1(VCC_net), .CO(n38734));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n38732), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n38732), .I0(n2728), 
            .I1(VCC_net), .CO(n38733));
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n38731), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n38731), .I0(n2729), 
            .I1(GND_net), .CO(n38732));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n38730), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14627_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5210), 
            .I3(n26334), .O(n28138));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14627_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14628_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4), .I3(n26339), 
            .O(n28139));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14628_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14721_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n23568), .I3(GND_net), .O(n28232));   // verilog/coms.v(127[12] 300[6])
    defparam i14721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14629_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4), .I3(n26334), 
            .O(n28140));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14629_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n38730), .I0(n2730), 
            .I1(GND_net), .CO(n38731));
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n38729), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n38729), .I0(n2731), 
            .I1(VCC_net), .CO(n38730));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n38728), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n38728), .I0(n2732), 
            .I1(GND_net), .CO(n38729));
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n38727), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_10 (.CI(n38098), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n38099));
    SB_LUT4 add_145_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n38097), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n38727), .I0(n2733), 
            .I1(VCC_net), .CO(n38728));
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n38117), .O(n1081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n38727));
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n48634), .I1(n2610), 
            .I2(VCC_net), .I3(n38726), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n38725), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n38725), .I0(n2611), 
            .I1(VCC_net), .CO(n38726));
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n38724), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n38724), .I0(n2612), 
            .I1(VCC_net), .CO(n38725));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n38723), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n38723), .I0(n2613), 
            .I1(VCC_net), .CO(n38724));
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n38722), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n38722), .I0(n2614), 
            .I1(VCC_net), .CO(n38723));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25_adj_5233), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n950));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n38721), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n38721), .I0(n2615), 
            .I1(VCC_net), .CO(n38722));
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n38720), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n38720), .I0(n2616), 
            .I1(VCC_net), .CO(n38721));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n38719), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n38719), .I0(n2617), 
            .I1(VCC_net), .CO(n38720));
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n38718), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n38091), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14998_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n42843), .I3(GND_net), .O(n28509));   // verilog/coms.v(127[12] 300[6])
    defparam i14998_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_184 (.Q(GHC), .C(CLK_c), .E(n27564), .D(GHC_N_403), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n38718), .I0(n2618), 
            .I1(VCC_net), .CO(n38719));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n38717), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHB_182 (.Q(GHB), .C(CLK_c), .E(n27564), .D(GHB_N_389), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n38717), .I0(n2619), 
            .I1(VCC_net), .CO(n38718));
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n2524), .I1(n2523), .I2(n2528), .I3(n2522), 
            .O(n45536));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n38716), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n38716), .I0(n2620), 
            .I1(VCC_net), .CO(n38717));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n38715), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n38715), .I0(n2621), 
            .I1(VCC_net), .CO(n38716));
    SB_LUT4 i14999_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n42843), .I3(GND_net), .O(n28510));   // verilog/coms.v(127[12] 300[6])
    defparam i14999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n2521), .I1(n2525), .I2(n2527), .I3(n2526), 
            .O(n45538));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_CARRY add_145_29 (.CI(n38117), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n38118));
    SB_LUT4 i15000_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n42843), .I3(GND_net), .O(n28511));   // verilog/coms.v(127[12] 300[6])
    defparam i15000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21070_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n34578));
    defparam i21070_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_145_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n38116), .O(n1082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n38714), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n2519), .I1(n2520), .I2(n45538), .I3(n45536), 
            .O(n45544));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n38714), .I0(n2622), 
            .I1(VCC_net), .CO(n38715));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n38713), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n2529), .I1(n34578), .I2(n2530), .I3(n2531), 
            .O(n43900));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n38713), .I0(n2623), 
            .I1(VCC_net), .CO(n38714));
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n38712), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n38712), .I0(n2624), 
            .I1(VCC_net), .CO(n38713));
    SB_LUT4 i15001_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n42843), .I3(GND_net), .O(n28512));   // verilog/coms.v(127[12] 300[6])
    defparam i15001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15002_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n42843), .I3(GND_net), .O(n28513));   // verilog/coms.v(127[12] 300[6])
    defparam i15002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n38711), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n2517), .I1(n43900), .I2(n2518), .I3(n45544), 
            .O(n45550));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n38711), .I0(n2625), 
            .I1(VCC_net), .CO(n38712));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n38710), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n38710), .I0(n2626), 
            .I1(VCC_net), .CO(n38711));
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n38709), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15003_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n42843), .I3(GND_net), .O(n28514));   // verilog/coms.v(127[12] 300[6])
    defparam i15003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15150_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n27595), 
            .I3(GND_net), .O(n28661));   // verilog/coms.v(127[12] 300[6])
    defparam i15150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n45550), 
            .O(n45556));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i15151_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28662));   // verilog/coms.v(127[12] 300[6])
    defparam i15151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33585_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n45556), 
            .O(n2544));
    defparam i33585_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15004_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n42843), .I3(GND_net), .O(n28515));   // verilog/coms.v(127[12] 300[6])
    defparam i15004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n38709), .I0(n2627), 
            .I1(VCC_net), .CO(n38710));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n38708), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n38708), .I0(n2628), 
            .I1(VCC_net), .CO(n38709));
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n38707), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n38707), .I0(n2629), 
            .I1(GND_net), .CO(n38708));
    SB_LUT4 i15005_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n42843), .I3(GND_net), .O(n28516));   // verilog/coms.v(127[12] 300[6])
    defparam i15005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n38706), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n38706), .I0(n2630), 
            .I1(GND_net), .CO(n38707));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n38705), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n38705), .I0(n2631), 
            .I1(VCC_net), .CO(n38706));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n38704), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n38704), .I0(n2632), 
            .I1(GND_net), .CO(n38705));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n38703), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n38703), .I0(n2633), 
            .I1(VCC_net), .CO(n38704));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n38703));
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n48659), .I1(n2511), 
            .I2(VCC_net), .I3(n38702), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n38701), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n38701), .I0(n2512), 
            .I1(VCC_net), .CO(n38702));
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n38700), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n38700), .I0(n2513), 
            .I1(VCC_net), .CO(n38701));
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n38699), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n38699), .I0(n2514), 
            .I1(VCC_net), .CO(n38700));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n38698), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n38698), .I0(n2515), 
            .I1(VCC_net), .CO(n38699));
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n38697), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n38697), .I0(n2516), 
            .I1(VCC_net), .CO(n38698));
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n38696), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n38696), .I0(n2517), 
            .I1(VCC_net), .CO(n38697));
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n38695), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n38695), .I0(n2518), 
            .I1(VCC_net), .CO(n38696));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n38694), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n38694), .I0(n2519), 
            .I1(VCC_net), .CO(n38695));
    SB_LUT4 encoder0_position_31__I_0_i1593_rep_25_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1593_rep_25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n38693), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15018_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n45341), .I3(GND_net), 
            .O(n28529));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15018_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n38693), .I0(n2520), 
            .I1(VCC_net), .CO(n38694));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n38692), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n38692), .I0(n2521), 
            .I1(VCC_net), .CO(n38693));
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n38691), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n38691), .I0(n2522), 
            .I1(VCC_net), .CO(n38692));
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n38690), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_9 (.CI(n38097), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n38098));
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n38690), .I0(n2523), 
            .I1(VCC_net), .CO(n38691));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24_adj_5234), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n949));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28540_3_lut (.I0(n4_adj_5222), .I1(n7647), .I2(n43549), .I3(GND_net), 
            .O(n43556));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_28 (.CI(n38116), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n38117));
    SB_LUT4 i15023_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n27595), 
            .I3(GND_net), .O(n28534));   // verilog/coms.v(127[12] 300[6])
    defparam i15023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n38689), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n38689), .I0(n2524), 
            .I1(VCC_net), .CO(n38690));
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n38688), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n38688), .I0(n2525), 
            .I1(VCC_net), .CO(n38689));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n38687), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n38687), .I0(n2526), 
            .I1(VCC_net), .CO(n38688));
    SB_LUT4 i15025_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n45261), .I3(GND_net), 
            .O(n28536));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n38115), .O(n1083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15026_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n45261), .I3(GND_net), 
            .O(n28537));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n38686), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15027_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n45261), .I3(GND_net), 
            .O(n28538));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15027_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15169_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n27596), .I3(GND_net), .O(n28680));   // verilog/coms.v(127[12] 300[6])
    defparam i15169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15170_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n27596), .I3(GND_net), .O(n28681));   // verilog/coms.v(127[12] 300[6])
    defparam i15170_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n38686), .I0(n2527), 
            .I1(VCC_net), .CO(n38687));
    SB_LUT4 i15028_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n45261), .I3(GND_net), 
            .O(n28539));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n62), .I3(delay_counter[31]), .O(n6_adj_5266));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h00b0;
    SB_LUT4 encoder0_position_31__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32806_3_lut (.I0(n2224), .I1(n2291), .I2(n2247), .I3(GND_net), 
            .O(n2323));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32807_3_lut (.I0(n2323), .I1(n2390), .I2(n2346), .I3(GND_net), 
            .O(n2422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n38685), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n38685), .I0(n2528), 
            .I1(VCC_net), .CO(n38686));
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n38684), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n38684), .I0(n2529), 
            .I1(GND_net), .CO(n38685));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n38683), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_27 (.CI(n38115), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n38116));
    SB_LUT4 i15029_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n45261), .I3(GND_net), 
            .O(n28540));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15029_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n38683), .I0(n2530), 
            .I1(GND_net), .CO(n38684));
    SB_LUT4 encoder0_position_31__I_0_i1584_3_lut (.I0(n46237), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1587_3_lut (.I0(n46235), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15030_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n45261), .I3(GND_net), 
            .O(n28541));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15030_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n38682), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n38682), .I0(n2531), 
            .I1(VCC_net), .CO(n38683));
    SB_LUT4 add_145_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n38114), .O(n1084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n38681), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n38681), .I0(n2532), 
            .I1(GND_net), .CO(n38682));
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n38680), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n38680), .I0(n2533), 
            .I1(VCC_net), .CO(n38681));
    SB_LUT4 i2_3_lut_adj_1697 (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n45261));
    defparam i2_3_lut_adj_1697.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15031_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n45261), .I3(GND_net), 
            .O(n28542));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n46240), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n46236), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28541_3_lut (.I0(encoder0_position[29]), .I1(n43556), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28541_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n38680));
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n48719), .I1(n2412), 
            .I2(VCC_net), .I3(n38679), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n38678), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n38678), .I0(n2413), 
            .I1(VCC_net), .CO(n38679));
    SB_LUT4 i15033_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n27595), 
            .I3(GND_net), .O(n28544));   // verilog/coms.v(127[12] 300[6])
    defparam i15033_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_26 (.CI(n38114), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n38115));
    SB_LUT4 i15034_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n27595), 
            .I3(GND_net), .O(n28545));   // verilog/coms.v(127[12] 300[6])
    defparam i15034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n38677), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n38677), .I0(n2414), 
            .I1(VCC_net), .CO(n38678));
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15036_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n44588), .I3(GND_net), .O(n28547));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15037_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n44588), .I3(GND_net), .O(n28548));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n38676), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n38676), .I0(n2415), 
            .I1(VCC_net), .CO(n38677));
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n38675), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n38675), .I0(n2416), 
            .I1(VCC_net), .CO(n38676));
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n38674), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15038_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n44588), .I3(GND_net), .O(n28549));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15039_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n44588), .I3(GND_net), .O(n28550));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15039_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n38674), .I0(n2417), 
            .I1(VCC_net), .CO(n38675));
    SB_DFFESR GHA_180 (.Q(GHA), .C(CLK_c), .E(n27564), .D(GHA_N_367), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n38673), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n38673), .I0(n2418), 
            .I1(VCC_net), .CO(n38674));
    SB_LUT4 i15040_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n44588), .I3(GND_net), .O(n28551));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2), .I3(n38425), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n38672), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n38672), .I0(n2419), 
            .I1(VCC_net), .CO(n38673));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5203), .I3(n38424), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n38424), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5203), .CO(n38425));
    SB_LUT4 i15041_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n44588), .I3(GND_net), .O(n28552));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n38671), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n38671), .I0(n2420), 
            .I1(VCC_net), .CO(n38672));
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n38670), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5202), .I3(n38423), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n7072), 
            .D(n1097), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n38670), .I0(n2421), 
            .I1(VCC_net), .CO(n38671));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n38669), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n38669), .I0(n2422), 
            .I1(VCC_net), .CO(n38670));
    SB_LUT4 i1_3_lut_adj_1698 (.I0(n5_adj_5182), .I1(n3_adj_5251), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n45760));
    defparam i1_3_lut_adj_1698.LUT_INIT = 16'h8080;
    SB_LUT4 i15042_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n44588), .I3(GND_net), .O(n28553));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14722_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n23568), .I3(GND_net), .O(n28233));   // verilog/coms.v(127[12] 300[6])
    defparam i14722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n38668), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n2425), .I1(n2423), .I2(n2428), .I3(n2427), 
            .O(n45840));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1700 (.I0(n2424), .I1(n2422), .I2(n2426), .I3(GND_net), 
            .O(n45838));
    defparam i1_3_lut_adj_1700.LUT_INIT = 16'hfefe;
    SB_LUT4 i15043_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n44588), .I3(GND_net), .O(n28554));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21076_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n34584));
    defparam i21076_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n7072), 
            .D(n1096), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n2420), .I1(n45838), .I2(n2421), .I3(n45840), 
            .O(n45846));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i14906_3_lut_4_lut (.I0(n1673), .I1(b_prev_adj_5209), .I2(a_new_adj_5349[1]), 
            .I3(direction_N_3907_adj_5211), .O(n28417));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14906_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i15044_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n44588), .I3(GND_net), .O(n28555));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15044_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n38668), .I0(n2423), 
            .I1(VCC_net), .CO(n38669));
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n2429), .I1(n34584), .I2(n2430), .I3(n2431), 
            .O(n43926));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n2418), .I1(n2419), .I2(n43926), .I3(n45846), 
            .O(n45852));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_5178), .I1(n7645), 
            .I2(n45760), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n45852), 
            .O(n45858));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i15045_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n44588), .I3(GND_net), .O(n28556));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33642_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n45858), 
            .O(n2445));
    defparam i33642_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n38667), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28542_3_lut (.I0(n3_adj_5251), .I1(n7646), .I2(n43549), .I3(GND_net), 
            .O(n43558));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15046_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n44588), .I3(GND_net), .O(n28557));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15047_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n44588), .I3(GND_net), .O(n28558));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15048_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n44588), .I3(GND_net), .O(n28559));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15048_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n38667), .I0(n2424), 
            .I1(VCC_net), .CO(n38668));
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5252), .D(commutation_state_7__N_216[0]), .S(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n38666), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n38666), .I0(n2425), 
            .I1(VCC_net), .CO(n38667));
    SB_LUT4 i15049_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n44588), .I3(GND_net), .O(n28560));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28543_3_lut (.I0(encoder0_position[30]), .I1(n43558), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15050_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n44588), .I3(GND_net), .O(n28561));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15051_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n44588), .I3(GND_net), .O(n28562));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15052_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n44588), .I3(GND_net), .O(n28563));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15053_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n44588), .I3(GND_net), .O(n28564));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15054_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n44588), .I3(GND_net), .O(n28565));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15055_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n44588), .I3(GND_net), .O(n28566));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15056_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n44588), .I3(GND_net), .O(n28567));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15057_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n44588), .I3(GND_net), .O(n28568));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n38665), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15058_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n44588), .I3(GND_net), .O(n28569));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1519_rep_30_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_rep_30_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15059_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n44588), .I3(GND_net), .O(n28570));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15060_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n44588), .I3(GND_net), .O(n28571));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15061_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n44588), .I3(GND_net), .O(n28572));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15062_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n44588), .I3(GND_net), .O(n28573));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15062_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n38665), .I0(n2426), 
            .I1(VCC_net), .CO(n38666));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n38664), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n38664), .I0(n2427), 
            .I1(VCC_net), .CO(n38665));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n38663), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n38663), .I0(n2428), 
            .I1(VCC_net), .CO(n38664));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n38423), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5202), .CO(n38424));
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n38662), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n38662), .I0(n2429), 
            .I1(GND_net), .CO(n38663));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5201), .I3(n38422), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n38127), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n38661), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n38661), .I0(n2430), 
            .I1(GND_net), .CO(n38662));
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n38660), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n38422), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5201), .CO(n38423));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5200), .I3(n38421), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15063_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n44588), .I3(GND_net), .O(n28574));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15063_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n38660), .I0(n2431), 
            .I1(VCC_net), .CO(n38661));
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n38659), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n38659), .I0(n2432), 
            .I1(GND_net), .CO(n38660));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n38658), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n38421), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5200), .CO(n38422));
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n38658), .I0(n2433), 
            .I1(VCC_net), .CO(n38659));
    SB_LUT4 add_145_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n38113), .O(n1085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5199), .I3(n38420), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n38658));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n48687), .I1(n2313), 
            .I2(VCC_net), .I3(n38657), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n38656), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n38420), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5199), .CO(n38421));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5198), .I3(n38419), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n38419), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5198), .CO(n38420));
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n38656), .I0(n2314), 
            .I1(VCC_net), .CO(n38657));
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n38655), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5197), .I3(n38418), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n38655), .I0(n2315), 
            .I1(VCC_net), .CO(n38656));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n38418), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5197), .CO(n38419));
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n38654), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n38654), .I0(n2316), 
            .I1(VCC_net), .CO(n38655));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n38653), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n38653), .I0(n2317), 
            .I1(VCC_net), .CO(n38654));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5196), .I3(n38417), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n38652), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_25 (.CI(n38113), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n38114));
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n38652), .I0(n2318), 
            .I1(VCC_net), .CO(n38653));
    SB_LUT4 add_145_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n38096), .O(n1102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n38651), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n38417), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5196), .CO(n38418));
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n38651), .I0(n2319), 
            .I1(VCC_net), .CO(n38652));
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n38650), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n38112), .O(n1086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n38650), .I0(n2320), 
            .I1(VCC_net), .CO(n38651));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5195), .I3(n38416), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n38416), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5195), .CO(n38417));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5194), .I3(n38415), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n38649), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n38415), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5194), .CO(n38416));
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n38649), .I0(n2321), 
            .I1(VCC_net), .CO(n38650));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n38648), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n38648), .I0(n2322), 
            .I1(VCC_net), .CO(n38649));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n38647), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n38647), .I0(n2323), 
            .I1(VCC_net), .CO(n38648));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n46240), 
            .I2(VCC_net), .I3(n38646), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_24 (.CI(n38112), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n38113));
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n38646), .I0(n46240), 
            .I1(VCC_net), .CO(n38647));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n46237), 
            .I2(VCC_net), .I3(n38645), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n38111), .O(n1087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n38645), .I0(n46237), 
            .I1(VCC_net), .CO(n38646));
    SB_CARRY add_145_8 (.CI(n38096), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n38097));
    SB_CARRY add_145_23 (.CI(n38111), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n38112));
    SB_LUT4 add_145_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n38110), .O(n1088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n46236), 
            .I2(VCC_net), .I3(n38644), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5193), .I3(n38414), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n38644), .I0(n46236), 
            .I1(VCC_net), .CO(n38645));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n38643), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n38643), .I0(n2327), 
            .I1(VCC_net), .CO(n38644));
    SB_LUT4 i15064_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n44588), .I3(GND_net), .O(n28575));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_rep_27_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n46236));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1518_rep_27_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23_adj_5235), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n948));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15065_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n44588), .I3(GND_net), .O(n28576));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1520_rep_26_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n46235));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1520_rep_26_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14865_3_lut_4_lut (.I0(n1632), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3907), .O(n28376));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14865_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_31__I_0_i1517_rep_28_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n46237));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1517_rep_28_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GLA_181 (.Q(INLA_c_0), .C(CLK_c), .E(n27564), .D(GLA_N_384), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 add_145_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n38095), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n46235), 
            .I2(VCC_net), .I3(n38642), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n7072), 
            .D(n1095), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n38414), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5193), .CO(n38415));
    SB_LUT4 i15066_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n44588), .I3(GND_net), .O(n28577));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15066_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n7072), 
            .D(n1094), .R(n28015));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n38642), .I0(n46235), 
            .I1(VCC_net), .CO(n38643));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n38641), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n38641), .I0(n2329), 
            .I1(GND_net), .CO(n38642));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n38640), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5192), .I3(n38413), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_22 (.CI(n38110), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n38111));
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n38640), .I0(n2330), 
            .I1(GND_net), .CO(n38641));
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n38639), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n38639), .I0(n2331), 
            .I1(VCC_net), .CO(n38640));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7), .I2(encoder0_position[31]), .I3(GND_net), .O(n731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n4_adj_5222), .I1(n5), .I2(n731), .I3(n6_adj_5229), 
            .O(n5_adj_5182));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'heeea;
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n38638), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1516_rep_31_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n46240));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1516_rep_31_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n38638), .I0(n2332), 
            .I1(GND_net), .CO(n38639));
    SB_DFFESR GLB_183 (.Q(INLB_c_0), .C(CLK_c), .E(n27564), .D(GLB_N_398), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n46240), .I1(n2323), .I2(n46237), .I3(n46235), 
            .O(n45590));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1707 (.I0(n46236), .I1(n2322), .I2(n2327), .I3(GND_net), 
            .O(n45588));
    defparam i1_3_lut_adj_1707.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n38637), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n38637), .I0(n2333), 
            .I1(VCC_net), .CO(n38638));
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n38637));
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n48746), .I1(n2214), 
            .I2(VCC_net), .I3(n38636), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n38635), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n38635), .I0(n2215), 
            .I1(VCC_net), .CO(n38636));
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n38634), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n38413), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5192), .CO(n38414));
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n38634), .I0(n2216), 
            .I1(VCC_net), .CO(n38635));
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n38633), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n38633), .I0(n2217), 
            .I1(VCC_net), .CO(n38634));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n38632), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n38632), .I0(n2218), 
            .I1(VCC_net), .CO(n38633));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n38631), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n38631), .I0(n2219), 
            .I1(VCC_net), .CO(n38632));
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n38630), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n38630), .I0(n2220), 
            .I1(VCC_net), .CO(n38631));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n38629), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n38629), .I0(n2221), 
            .I1(VCC_net), .CO(n38630));
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n38628), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1708 (.I0(n3_adj_5251), .I1(n2_adj_5178), .I2(n5_adj_5182), 
            .I3(GND_net), .O(n43549));
    defparam i1_3_lut_adj_1708.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n38628), .I0(n2222), 
            .I1(VCC_net), .CO(n38629));
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n38627), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n38627), .I0(n2223), 
            .I1(VCC_net), .CO(n38628));
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n38626), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n38626), .I0(n2224), 
            .I1(VCC_net), .CO(n38627));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n38625), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n38625), .I0(n2225), 
            .I1(VCC_net), .CO(n38626));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5191), .I3(n38412), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n38624), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n38624), .I0(n2226), 
            .I1(VCC_net), .CO(n38625));
    SB_LUT4 i28534_rep_56_3_lut (.I0(n7), .I1(n7650), .I2(n43549), .I3(GND_net), 
            .O(n46265));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28534_rep_56_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28589_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n36539), .I3(GND_net), .O(n43608));
    defparam i28589_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n38623), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n38109), .O(n1089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n38623), .I0(n2227), 
            .I1(VCC_net), .CO(n38624));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n38622), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n38622), .I0(n2228), 
            .I1(VCC_net), .CO(n38623));
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n38621), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n38621), .I0(n2229), 
            .I1(GND_net), .CO(n38622));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n38620), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n38412), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5191), .CO(n38413));
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n38620), .I0(n2230), 
            .I1(GND_net), .CO(n38621));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n38619), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5190), .I3(n38411), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n38619), .I0(n2231), 
            .I1(VCC_net), .CO(n38620));
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n38618), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n38411), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5190), .CO(n38412));
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n38618), .I0(n2232), 
            .I1(GND_net), .CO(n38619));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n38617), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n38617), .I0(n2233), 
            .I1(VCC_net), .CO(n38618));
    SB_LUT4 i21149_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n34658));
    defparam i21149_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n38617));
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n2320), .I1(n2321), .I2(n45588), .I3(n45590), 
            .O(n45596));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1710 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n45796));
    defparam i1_2_lut_adj_1710.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n45796), .I1(n2319), .I2(n45596), .I3(n34658), 
            .O(n45600));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n45600), 
            .O(n45606));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n48186), .I1(n2115), 
            .I2(VCC_net), .I3(n38616), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33611_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n45606), 
            .O(n2346));
    defparam i33611_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n38615), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n38615), .I0(n2116), 
            .I1(VCC_net), .CO(n38616));
    SB_CARRY add_145_3 (.CI(n38091), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n38092));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n38614), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5189), .I3(n38410), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n38614), .I0(n2117), 
            .I1(VCC_net), .CO(n38615));
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n38613), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n38613), .I0(n2118), 
            .I1(VCC_net), .CO(n38614));
    SB_LUT4 add_2625_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n38203), 
            .O(n7645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n38612), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n38612), .I0(n2119), 
            .I1(VCC_net), .CO(n38613));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n38611), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n38611), .I0(n2120), 
            .I1(VCC_net), .CO(n38612));
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n38610), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n38410), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5189), .CO(n38411));
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n38610), .I0(n2121), 
            .I1(VCC_net), .CO(n38611));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n38609), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2625_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n38202), 
            .O(n7646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n38609), .I0(n2122), 
            .I1(VCC_net), .CO(n38610));
    SB_CARRY add_2625_6 (.CI(n38202), .I0(n622), .I1(GND_net), .CO(n38203));
    SB_LUT4 add_145_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5188), .I3(n38409), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n38409), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5188), .CO(n38410));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n38608), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5187), .I3(n38408), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n38608), .I0(n2123), 
            .I1(VCC_net), .CO(n38609));
    SB_LUT4 i28535_3_lut (.I0(encoder0_position[26]), .I1(n46265), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2625_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n38201), 
            .O(n7647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n38607), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n38607), .I0(n2124), 
            .I1(VCC_net), .CO(n38608));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n38606), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n38606), .I0(n2125), 
            .I1(VCC_net), .CO(n38607));
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n38605), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_7 (.CI(n38095), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n38096));
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n38605), .I0(n2126), 
            .I1(VCC_net), .CO(n38606));
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n38604), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2625_5 (.CI(n38201), .I0(n623), .I1(VCC_net), .CO(n38202));
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n38604), .I0(n2127), 
            .I1(VCC_net), .CO(n38605));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n38408), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5187), .CO(n38409));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n38603), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n38603), .I0(n2128), 
            .I1(VCC_net), .CO(n38604));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n38602), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5186), .I3(n38407), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n38602), .I0(n2129), 
            .I1(GND_net), .CO(n38603));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n38601), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n38601), .I0(n2130), 
            .I1(GND_net), .CO(n38602));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n38407), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5186), .CO(n38408));
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n38600), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28536_3_lut (.I0(n6_adj_5229), .I1(n7649), .I2(n43549), .I3(GND_net), 
            .O(n43552));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28536_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n38600), .I0(n2131), 
            .I1(VCC_net), .CO(n38601));
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n38599), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n38144), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n38599), .I0(n2132), 
            .I1(GND_net), .CO(n38600));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n38598), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5185), .I3(n38406), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n38598), .I0(n2133), 
            .I1(VCC_net), .CO(n38599));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n38598));
    SB_CARRY add_145_21 (.CI(n38109), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n38110));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n48209), .I1(n2016), 
            .I2(VCC_net), .I3(n38597), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n38596), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n38406), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5185), .CO(n38407));
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n38596), .I0(n2017), 
            .I1(VCC_net), .CO(n38597));
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n38595), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n38091));
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n38595), .I0(n2018), 
            .I1(VCC_net), .CO(n38596));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n38594), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5184), .I3(n38405), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n38594), .I0(n2019), 
            .I1(VCC_net), .CO(n38595));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n38405), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5184), .CO(n38406));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n38593), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n38593), .I0(n2020), 
            .I1(VCC_net), .CO(n38594));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n38592), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28537_3_lut (.I0(encoder0_position[27]), .I1(n43552), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28537_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n38592), .I0(n2021), 
            .I1(VCC_net), .CO(n38593));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5183), .I3(n38404), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n38591), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n38591), .I0(n2022), 
            .I1(VCC_net), .CO(n38592));
    SB_LUT4 add_2625_4_lut (.I0(GND_net), .I1(n405), .I2(GND_net), .I3(n38200), 
            .O(n7648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n38590), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n38590), .I0(n2023), 
            .I1(VCC_net), .CO(n38591));
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n38589), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n38404), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5183), .CO(n38405));
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n38589), .I0(n2024), 
            .I1(VCC_net), .CO(n38590));
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n38588), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n38588), .I0(n2025), 
            .I1(VCC_net), .CO(n38589));
    SB_CARRY add_2625_4 (.CI(n38200), .I0(n405), .I1(GND_net), .CO(n38201));
    SB_LUT4 i28538_3_lut (.I0(n5), .I1(n7648), .I2(n43549), .I3(GND_net), 
            .O(n43554));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n38587), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n38587), .I0(n2026), 
            .I1(VCC_net), .CO(n38588));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5181), .I3(n38403), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n38586), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2625_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n38199), 
            .O(n7649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n38094), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n38586), .I0(n2027), 
            .I1(VCC_net), .CO(n38587));
    SB_CARRY add_2625_3 (.CI(n38199), .I0(n625), .I1(VCC_net), .CO(n38200));
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n38585), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n38585), .I0(n2028), 
            .I1(VCC_net), .CO(n38586));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n38584), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n38584), .I0(n2029), 
            .I1(GND_net), .CO(n38585));
    SB_LUT4 add_2625_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n38583), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n38583), .I0(n2030), 
            .I1(GND_net), .CO(n38584));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n38582), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n38582), .I0(n2031), 
            .I1(VCC_net), .CO(n38583));
    SB_CARRY add_145_6 (.CI(n38094), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n38095));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n38403), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5181), .CO(n38404));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n38581), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n38581), .I0(n2032), 
            .I1(GND_net), .CO(n38582));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n38580), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n38143), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_24 (.CI(n38143), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n38144));
    SB_CARRY add_2625_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n38199));
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n38580), .I0(n2033), 
            .I1(VCC_net), .CO(n38581));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5180), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n38580));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5180), .CO(n38403));
    SB_LUT4 unary_minus_10_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_215), 
            .I3(n38198), .O(pwm_setpoint_23__N_191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n48230), .I1(n1917), 
            .I2(VCC_net), .I3(n38579), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n38578), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n38578), .I0(n1918), 
            .I1(VCC_net), .CO(n38579));
    SB_LUT4 add_224_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n38142), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3), 
            .I3(n38197), .O(pwm_setpoint_23__N_191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n38577), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n38577), .I0(n1919), 
            .I1(VCC_net), .CO(n38578));
    SB_LUT4 add_145_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n38108), .O(n1090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n38576), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n38576), .I0(n1920), 
            .I1(VCC_net), .CO(n38577));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n38575), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n38575), .I0(n1921), 
            .I1(VCC_net), .CO(n38576));
    SB_CARRY unary_minus_10_add_3_24 (.CI(n38197), .I0(GND_net), .I1(n3), 
            .CO(n38198));
    SB_CARRY add_224_23 (.CI(n38142), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n38143));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n38574), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n38574), .I0(n1922), 
            .I1(VCC_net), .CO(n38575));
    SB_LUT4 i28539_3_lut (.I0(encoder0_position[28]), .I1(n43554), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i28539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n38573), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n38573), .I0(n1923), 
            .I1(VCC_net), .CO(n38574));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n38572), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4_adj_5162), 
            .I3(n38196), .O(pwm_setpoint_23__N_191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n38572), .I0(n1924), 
            .I1(VCC_net), .CO(n38573));
    SB_LUT4 add_224_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n38141), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_23 (.CI(n38196), .I0(GND_net), .I1(n4_adj_5162), 
            .CO(n38197));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n38571), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n38571), .I0(n1925), 
            .I1(VCC_net), .CO(n38572));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n38570), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n38570), .I0(n1926), 
            .I1(VCC_net), .CO(n38571));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n38569), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n38569), .I0(n1927), 
            .I1(VCC_net), .CO(n38570));
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n38568), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_20 (.CI(n38108), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n38109));
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n38568), .I0(n1928), 
            .I1(VCC_net), .CO(n38569));
    SB_LUT4 add_145_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n38107), .O(n1091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n38567), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n38567), .I0(n1929), 
            .I1(GND_net), .CO(n38568));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n38566), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n38566), .I0(n1930), 
            .I1(GND_net), .CO(n38567));
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n38565), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_22 (.CI(n38141), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n38142));
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n38565), .I0(n1931), 
            .I1(VCC_net), .CO(n38566));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n38564), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n38564), .I0(n1932), 
            .I1(GND_net), .CO(n38565));
    SB_LUT4 i21145_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n34654));
    defparam i21145_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_224_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n38140), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n38563), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n38563), .I0(n1933), 
            .I1(VCC_net), .CO(n38564));
    SB_CARRY add_224_21 (.CI(n38140), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n38141));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21265_4_lut (.I0(n829), .I1(n828), .I2(n34654), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i21265_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 add_224_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n38139), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n38563));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n48248), .I1(n1818), 
            .I2(VCC_net), .I3(n38562), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n38561), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_20 (.CI(n38139), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n38140));
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n38561), .I0(n1819), 
            .I1(VCC_net), .CO(n38562));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n38560), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5_adj_5163), 
            .I3(n38195), .O(pwm_setpoint_23__N_191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n38560), .I0(n1820), 
            .I1(VCC_net), .CO(n38561));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n38559), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n38559), .I0(n1821), 
            .I1(VCC_net), .CO(n38560));
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n38558), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n38558), .I0(n1822), 
            .I1(VCC_net), .CO(n38559));
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n38557), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n38557), .I0(n1823), 
            .I1(VCC_net), .CO(n38558));
    SB_CARRY add_145_19 (.CI(n38107), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n38108));
    SB_CARRY unary_minus_10_add_3_22 (.CI(n38195), .I0(GND_net), .I1(n5_adj_5163), 
            .CO(n38196));
    SB_LUT4 add_145_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n38106), .O(n1092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n38556), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n38556), .I0(n1824), 
            .I1(VCC_net), .CO(n38557));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n38555), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n38555), .I0(n1825), 
            .I1(VCC_net), .CO(n38556));
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n38554), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n38554), .I0(n1826), 
            .I1(VCC_net), .CO(n38555));
    SB_LUT4 unary_minus_10_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6), 
            .I3(n38194), .O(pwm_setpoint_23__N_191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n38553), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n38553), .I0(n1827), 
            .I1(VCC_net), .CO(n38554));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n38552), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_21 (.CI(n38194), .I0(GND_net), .I1(n6), 
            .CO(n38195));
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n38552), .I0(n1828), 
            .I1(VCC_net), .CO(n38553));
    SB_LUT4 unary_minus_10_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7_adj_5164), 
            .I3(n38193), .O(pwm_setpoint_23__N_191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n38551), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n38138), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n38551), .I0(n1829), 
            .I1(GND_net), .CO(n38552));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n38550), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n38550), .I0(n1830), 
            .I1(GND_net), .CO(n38551));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n38549), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_18 (.CI(n38106), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n38107));
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n38549), .I0(n1831), 
            .I1(VCC_net), .CO(n38550));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n38548), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n38105), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n38548), .I0(n1832), 
            .I1(GND_net), .CO(n38549));
    SB_LUT4 i14667_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n23568), .I3(GND_net), .O(n28178));   // verilog/coms.v(127[12] 300[6])
    defparam i14667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n38547), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n38547), .I0(n1833), 
            .I1(VCC_net), .CO(n38548));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n38547));
    SB_CARRY unary_minus_10_add_3_20 (.CI(n38193), .I0(GND_net), .I1(n7_adj_5164), 
            .CO(n38194));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n48271), .I1(n1719), 
            .I2(VCC_net), .I3(n38546), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n38545), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n38545), .I0(n1720), 
            .I1(VCC_net), .CO(n38546));
    SB_LUT4 i33190_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48271));
    defparam i33190_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14668_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n23568), .I3(GND_net), .O(n28179));   // verilog/coms.v(127[12] 300[6])
    defparam i14668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n38544), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n38544), .I0(n1721), 
            .I1(VCC_net), .CO(n38545));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n38543), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n38543), .I0(n1722), 
            .I1(VCC_net), .CO(n38544));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n38542), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n38542), .I0(n1723), 
            .I1(VCC_net), .CO(n38543));
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n38541), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n38541), .I0(n1724), 
            .I1(VCC_net), .CO(n38542));
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n38540), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n38540), .I0(n1725), 
            .I1(VCC_net), .CO(n38541));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n38539), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n43638));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY add_224_19 (.CI(n38138), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n38139));
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n28542));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n28541));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n28540));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n38539), .I0(n1726), 
            .I1(VCC_net), .CO(n38540));
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n28539));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n28538));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n28537));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n28536));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 unary_minus_10_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8), 
            .I3(n38192), .O(pwm_setpoint_23__N_191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_19 (.CI(n38192), .I0(GND_net), .I1(n8), 
            .CO(n38193));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n38538), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n38538), .I0(n1727), 
            .I1(VCC_net), .CO(n38539));
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n38537), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n38537), .I0(n1728), 
            .I1(VCC_net), .CO(n38538));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5250), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n834));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n38536), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n38536), .I0(n1729), 
            .I1(GND_net), .CO(n38537));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n38535), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n38137), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n38535), .I0(n1730), 
            .I1(GND_net), .CO(n38536));
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n38534), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n38534), .I0(n1731), 
            .I1(VCC_net), .CO(n38535));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n38533), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n38533), .I0(n1732), 
            .I1(GND_net), .CO(n38534));
    SB_DFFESR GLC_185 (.Q(INLC_c_0), .C(CLK_c), .E(n27564), .D(GLC_N_412), 
            .R(n27904));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n38532), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n38532), .I0(n1733), 
            .I1(VCC_net), .CO(n38533));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n38191), .O(pwm_setpoint_23__N_191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n38532));
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_18 (.CI(n38191), .I0(GND_net), .I1(n9), 
            .CO(n38192));
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n48291), .I1(n1620), 
            .I2(VCC_net), .I3(n38531), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n38530), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n38530), .I0(n1621), 
            .I1(VCC_net), .CO(n38531));
    SB_LUT4 unary_minus_10_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10_adj_5165), 
            .I3(n38190), .O(pwm_setpoint_23__N_191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_17 (.CI(n38105), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n38106));
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n38529), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_17 (.CI(n38190), .I0(GND_net), .I1(n10_adj_5165), 
            .CO(n38191));
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n38529), .I0(n1622), 
            .I1(VCC_net), .CO(n38530));
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n38528), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n38528), .I0(n1623), 
            .I1(VCC_net), .CO(n38529));
    SB_LUT4 unary_minus_10_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11), 
            .I3(n38189), .O(pwm_setpoint_23__N_191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n38527), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_18 (.CI(n38137), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n38138));
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n38527), .I0(n1624), 
            .I1(VCC_net), .CO(n38528));
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n38526), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n38136), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n38526), .I0(n1625), 
            .I1(VCC_net), .CO(n38527));
    SB_CARRY add_224_17 (.CI(n38136), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n38137));
    SB_LUT4 add_145_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n38104), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n38525), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n38525), .I0(n1626), 
            .I1(VCC_net), .CO(n38526));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n38524), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_16 (.CI(n38104), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n38105));
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n28362));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY unary_minus_10_add_3_16 (.CI(n38189), .I0(GND_net), .I1(n11), 
            .CO(n38190));
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n38524), .I0(n1627), 
            .I1(VCC_net), .CO(n38525));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n38523), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n38523), .I0(n1628), 
            .I1(VCC_net), .CO(n38524));
    SB_LUT4 add_145_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n38103), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n38522), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n38522), .I0(n1629), 
            .I1(GND_net), .CO(n38523));
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n38521), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_15 (.CI(n38103), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n38104));
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n38521), .I0(n1630), 
            .I1(GND_net), .CO(n38522));
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n38520), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n38520), .I0(n1631), 
            .I1(VCC_net), .CO(n38521));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22_adj_5236), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n947));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF read_189 (.Q(read), .C(CLK_c), .D(n45320));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632_adj_5263), 
            .I2(GND_net), .I3(n38519), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n38519), .I0(n1632_adj_5263), 
            .I1(GND_net), .CO(n38520));
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n38518), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n38188), .O(pwm_setpoint_23__N_191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n38518), .I0(n1633), 
            .I1(VCC_net), .CO(n38519));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n38518));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n48309), .I1(n1521), 
            .I2(VCC_net), .I3(n38517), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_224_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n38135), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n38516), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n38516), .I0(n1522), 
            .I1(VCC_net), .CO(n38517));
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n38515), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n38515), .I0(n1523), 
            .I1(VCC_net), .CO(n38516));
    SB_CARRY add_224_16 (.CI(n38135), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n38136));
    SB_LUT4 add_145_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n38102), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n38514), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_15 (.CI(n38188), .I0(GND_net), .I1(n12), 
            .CO(n38189));
    SB_LUT4 unary_minus_10_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13), 
            .I3(n38187), .O(pwm_setpoint_23__N_191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n38514), .I0(n1524), 
            .I1(VCC_net), .CO(n38515));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n38513), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n38513), .I0(n1525), 
            .I1(VCC_net), .CO(n38514));
    SB_LUT4 add_224_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n38134), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n38512), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n38512), .I0(n1526), 
            .I1(VCC_net), .CO(n38513));
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n38511), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_15 (.CI(n38134), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n38135));
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n38511), .I0(n1527), 
            .I1(VCC_net), .CO(n38512));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n38510), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_14 (.CI(n38102), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n38103));
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n38510), .I0(n1528), 
            .I1(VCC_net), .CO(n38511));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n38509), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n38509), .I0(n1529), 
            .I1(GND_net), .CO(n38510));
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n38508), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n38508), .I0(n1530), 
            .I1(GND_net), .CO(n38509));
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n38507), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n38507), .I0(n1531), 
            .I1(VCC_net), .CO(n38508));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n38506), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n38506), .I0(n1532), 
            .I1(GND_net), .CO(n38507));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n38505), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n38505), .I0(n1533), 
            .I1(VCC_net), .CO(n38506));
    SB_CARRY unary_minus_10_add_3_14 (.CI(n38187), .I0(GND_net), .I1(n13), 
            .CO(n38188));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n38505));
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(GND_net), .I1(n1422), 
            .I2(VCC_net), .I3(n38504), .O(n1489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n38503), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    motorControl control (.GND_net(GND_net), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Ki[1] (Ki[1]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[9] (Ki[9]), .IntegralLimit({IntegralLimit}), 
            .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), 
            .\Ki[3] (Ki[3]), .\Ki[12] (Ki[12]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Kp[2] (Kp[2]), .\Ki[13] (Ki[13]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .duty({duty}), 
            .clk32MHz(clk32MHz), .VCC_net(VCC_net), .setpoint({setpoint}), 
            .motor_state({motor_state}), .PWMLimit({PWMLimit})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(271[16] 283[4])
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    GND i1 (.Y(GND_net));
    SB_LUT4 unary_minus_10_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n38186), .O(pwm_setpoint_23__N_191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n38503), .I0(n1423), 
            .I1(VCC_net), .CO(n38504));
    SB_LUT4 encoder0_position_31__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n38502), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n38502), .I0(n1424), 
            .I1(VCC_net), .CO(n38503));
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n38501), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_13 (.CI(n38186), .I0(GND_net), .I1(n14), 
            .CO(n38187));
    SB_LUT4 add_224_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n38133), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5166), 
            .I3(n38185), .O(pwm_setpoint_23__N_191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n38501), .I0(n1425), 
            .I1(VCC_net), .CO(n38502));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n38500), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n38500), .I0(n1426), 
            .I1(VCC_net), .CO(n38501));
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n38499), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n38499), .I0(n1427), 
            .I1(VCC_net), .CO(n38500));
    SB_CARRY unary_minus_10_add_3_12 (.CI(n38185), .I0(GND_net), .I1(n15_adj_5166), 
            .CO(n38186));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n38498), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33665_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48746));
    defparam i33665_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n2226), .I1(n2224), .I2(n2227), .I3(n2225), 
            .O(n45804));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n38498), .I0(n1428), 
            .I1(VCC_net), .CO(n38499));
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n38497), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21080_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n34588));
    defparam i21080_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n2222), .I1(n45804), .I2(n2223), .I3(n2228), 
            .O(n45808));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n2229), .I1(n34588), .I2(n2230), .I3(n2231), 
            .O(n43911));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n2220), .I1(n43911), .I2(n2221), .I3(n45808), 
            .O(n45814));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n38497), .I0(n1429), 
            .I1(GND_net), .CO(n38498));
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n38496), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n38496), .I0(n1430), 
            .I1(GND_net), .CO(n38497));
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21179_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n34688));
    defparam i21179_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n45814), 
            .O(n45820));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i33668_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n45820), 
            .O(n2247));
    defparam i33668_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i32286_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n47224));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32286_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i32300_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n47188));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32300_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i32299_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n47187));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32299_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1718 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n45668));
    defparam i1_2_lut_adj_1718.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1373_rep_40_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1373_rep_40_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32298_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n47186));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32298_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i32297_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n47185));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32297_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n927), .I1(n45668), .I2(n928), .I3(n34688), 
            .O(n960));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hfefa;
    SB_LUT4 i32296_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n47184));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32296_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i32247_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n47183));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32247_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32216_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n47182));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i32216_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5267), 
            .I2(commutation_state_prev[0]), .I3(dti_N_416), .O(n27540));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21_adj_5237), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n946));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5164));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.b_prev(b_prev), .GND_net(GND_net), 
            .a_new({a_new[1], Open_0}), .direction_N_3907(direction_N_3907), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1668(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .encoder0_position({encoder0_position}), .VCC_net(VCC_net), 
            .n28376(n28376), .n1632(n1632)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(285[57] 292[6])
    SB_LUT4 i28618_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n43638));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i28618_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33105_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48186));
    defparam i33105_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1720 (.I0(n2128), .I1(n2127), .I2(GND_net), .I3(GND_net), 
            .O(n45562));
    defparam i1_2_lut_adj_1720.LUT_INIT = 16'heeee;
    SB_LUT4 i5358_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_367));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i5358_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5249), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n934));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21153_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n34662));
    defparam i21153_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n2122), .I1(n2126), .I2(n45562), .I3(n2125), 
            .O(n45568));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n2129), .I1(n45568), .I2(n34662), .I3(n2130), 
            .O(n45570));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'heccc;
    SB_LUT4 i5360_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_384));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i5360_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n2118), .I1(n2119), .I2(n45570), .I3(n2120), 
            .O(n45576));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n2121), .I1(n2117), .I2(n2123), .I3(n2124), 
            .O(n44948));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_LUT4 i33108_4_lut (.I0(n44948), .I1(n2115), .I2(n2116), .I3(n45576), 
            .O(n2148));
    defparam i33108_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5248), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5163));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33167_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48248));
    defparam i33167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1321_rep_41_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1321_rep_41_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20_adj_5238), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n945));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33128_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48209));
    defparam i33128_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21086_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n34594));
    defparam i21086_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1725 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n45770));
    defparam i1_2_lut_adj_1725.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n2025), .I1(n45770), .I2(n2024), .I3(n2028), 
            .O(n45774));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n2029), .I1(n34594), .I2(n2030), .I3(n2031), 
            .O(n43904));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n45774), 
            .O(n45780));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n2019), .I1(n2020), .I2(n45780), .I3(n43904), 
            .O(n45786));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5298));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33131_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n45786), 
            .O(n2049));
    defparam i33131_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1730 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10), .I3(control_mode[2]), .O(n26211));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam i1_2_lut_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5297));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5296));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33696_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26226), .I3(GND_net), .O(n7072));
    defparam i33696_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19_adj_5239), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n944));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32324_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n47237));
    defparam i32324_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 unary_minus_10_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5162));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33149_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48230));
    defparam i33149_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5180));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1246_rep_44_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_rep_44_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1247_rep_43_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1247_rep_43_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1245_rep_45_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1245_rep_45_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1248_rep_42_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1248_rep_42_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n1928), .I1(n1925), .I2(n1927), .I3(n1926), 
            .O(n45616));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n29908), 
            .I2(n4452), .I3(GND_net), .O(n9_adj_5309));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i21088_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n34596));
    defparam i21088_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1732 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26226), .I3(GND_net), .O(n26227));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut_adj_1732.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n1922), .I1(n1923), .I2(n45616), .I3(n1924), 
            .O(n45622));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n1929), .I1(n34596), .I2(n1930), .I3(n1931), 
            .O(n43868));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n1920), .I1(n43868), .I2(n1921), .I3(n45622), 
            .O(n45628));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 i33153_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n45628), 
            .O(n1950));
    defparam i33153_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1173_rep_46_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1173_rep_46_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5229), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5388[2]), .I1(r_SM_Main_adj_5388[0]), 
            .I2(r_SM_Main_adj_5388[1]), .I3(r_SM_Main_2__N_3613[1]), .O(n48986));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1180_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1178_3_lut (.I0(n1727), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5181));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49_4_lut_4_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n6976), .I3(n47230), .O(n42022));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i49_4_lut_4_lut.LUT_INIT = 16'hf7c4;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5), .I2(encoder0_position[31]), .I3(GND_net), .O(n405));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_5240), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n943));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5183));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21090_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n34598));
    defparam i21090_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5184));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n1829), .I1(n34598), .I2(n1830), .I3(n1831), 
            .O(n43883));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n1822), .I1(n1824), .I2(n1826), .I3(n1828), 
            .O(n45746));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1738 (.I0(n1823), .I1(n1825), .I2(n1827), .I3(GND_net), 
            .O(n45830));
    defparam i1_3_lut_adj_1738.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n1821), .I1(n45830), .I2(n45746), .I3(n43883), 
            .O(n45750));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5185));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5186));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5222), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21102_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n34610));
    defparam i21102_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5187));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33174_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n45750), 
            .O(n1851));
    defparam i33174_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5188));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21108_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n34616));
    defparam i21108_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1740 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n45686));
    defparam i1_3_lut_adj_1740.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5251), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n1029), .I1(n34616), .I2(n1030), .I3(n1031), 
            .O(n43826));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4798_2_lut (.I0(n2_adj_5178), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4798_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5189));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14723_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n23568), .I3(GND_net), .O(n28234));   // verilog/coms.v(127[12] 300[6])
    defparam i14723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5190));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5191));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1117_rep_47_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1117_rep_47_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14577_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n23568), .I3(GND_net), .O(n28088));   // verilog/coms.v(127[12] 300[6])
    defparam i14577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4551_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(107[7:14])
    defparam i4551_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14578_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n23568), .I3(GND_net), .O(n28089));   // verilog/coms.v(127[12] 300[6])
    defparam i14578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632_adj_5263), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_5241), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n942));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5192));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    coms neopxl_color_23__I_0 (.n28234(n28234), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .CLK_c(CLK_c), .n28233(n28233), .n26879(n26879), .n28232(n28232), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n28231(n28231), 
         .n28230(n28230), .GND_net(GND_net), .n28229(n28229), .n28228(n28228), 
         .n28227(n28227), .n28226(n28226), .n28225(n28225), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\FRAME_MATCHER.state ({Open_1, 
         Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
         Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, 
         Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, Open_22, 
         Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, \FRAME_MATCHER.state [3:0]}), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[21][4] (\data_out_frame[21] [4]), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .rx_data_ready(rx_data_ready), 
         .n28224(n28224), .n28223(n28223), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n27595(n27595), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[21][2] (\data_out_frame[21] [2]), .n9(n9_adj_5309), 
         .n3813(n3813), .n4452(n4452), .n23534(n23534), .n29908(n29908), 
         .\FRAME_MATCHER.i_31__N_2626 (\FRAME_MATCHER.i_31__N_2626 ), .\data_in[0] ({\data_in[0] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[2] ({\data_in[2] }), .\data_in[3] ({\data_in[3] }), 
         .n28222(n28222), .n28221(n28221), .n3303(n3303), .n63(n63), 
         .\FRAME_MATCHER.i_31__N_2624 (\FRAME_MATCHER.i_31__N_2624 ), .\FRAME_MATCHER.i_31__N_2622 (\FRAME_MATCHER.i_31__N_2622 ), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .setpoint({setpoint}), 
         .n28220(n28220), .n28219(n28219), .n28218(n28218), .n28217(n28217), 
         .n28216(n28216), .n28215(n28215), .n28214(n28214), .n28213(n28213), 
         .n28212(n28212), .n28211(n28211), .n28210(n28210), .n28209(n28209), 
         .n28208(n28208), .n28207(n28207), .n27596(n27596), .n28206(n28206), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .n28205(n28205), .\data_out_frame[21][1] (\data_out_frame[21] [1]), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .n28204(n28204), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .n28203(n28203), .n28202(n28202), .\data_out_frame[21][0] (\data_out_frame[21] [0]), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_out_frame[21][3] (\data_out_frame[21] [3]), 
         .tx_active(tx_active), .n28200(n28200), .n36539(n36539), .n28199(n28199), 
         .n28198(n28198), .n28197(n28197), .n28196(n28196), .n28195(n28195), 
         .n28194(n28194), .n28193(n28193), .n28192(n28192), .n28191(n28191), 
         .n28190(n28190), .n28189(n28189), .n28188(n28188), .n28187(n28187), 
         .n28186(n28186), .n28185(n28185), .n28184(n28184), .n28183(n28183), 
         .n28182(n28182), .n28181(n28181), .n28180(n28180), .\data_out_frame[27][1] (\data_out_frame[27] [1]), 
         .ID({ID}), .n28179(n28179), .n28178(n28178), .rx_data({rx_data}), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n122(n122), .n5(n5_adj_5274), .n49229(n49229), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .n28177(n28177), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .n28176(n28176), .n28175(n28175), .n28715(n28715), .n28714(n28714), 
         .n28713(n28713), .n28712(n28712), .n28711(n28711), .n28710(n28710), 
         .neopxl_color({neopxl_color}), .n28709(n28709), .n28708(n28708), 
         .n28707(n28707), .n28706(n28706), .n28705(n28705), .n28704(n28704), 
         .n28703(n28703), .n28702(n28702), .n28701(n28701), .n28700(n28700), 
         .n28699(n28699), .n28698(n28698), .n28697(n28697), .n28696(n28696), 
         .n28695(n28695), .n28694(n28694), .n28693(n28693), .n28692(n28692), 
         .n28691(n28691), .n28690(n28690), .n28689(n28689), .n28688(n28688), 
         .n28687(n28687), .n28686(n28686), .n28685(n28685), .n28684(n28684), 
         .n28683(n28683), .n28174(n28174), .n28173(n28173), .n28172(n28172), 
         .n28171(n28171), .n28170(n28170), .n28169(n28169), .n28168(n28168), 
         .n28167(n28167), .n28166(n28166), .n28165(n28165), .n28164(n28164), 
         .n28163(n28163), .n28162(n28162), .n28161(n28161), .n28160(n28160), 
         .n28156(n28156), .n28152(n28152), .n28151(n28151), .n42180(n42180), 
         .n28149(n28149), .PWMLimit({PWMLimit}), .n28148(n28148), .control_mode({control_mode}), 
         .n28146(n28146), .n28145(n28145), .\Ki[0] (Ki[0]), .n28144(n28144), 
         .\Kp[0] (Kp[0]), .n28143(n28143), .DE_c(DE_c), .LED_c(LED_c), 
         .n28682(n28682), .n28681(n28681), .n28680(n28680), .n28662(n28662), 
         .n28661(n28661), .\Kp[1] (Kp[1]), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n28638(n28638), .n28637(n28637), .n28636(n28636), .n28635(n28635), 
         .\Kp[2] (Kp[2]), .n28634(n28634), .n28633(n28633), .n28632(n28632), 
         .n49000(n49000), .n28630(n28630), .n28629(n28629), .n28109(n28109), 
         .IntegralLimit({IntegralLimit}), .n28106(n28106), .n28105(n28105), 
         .n28104(n28104), .n28103(n28103), .n28102(n28102), .n28101(n28101), 
         .n28100(n28100), .n28099(n28099), .n28098(n28098), .n28097(n28097), 
         .n28095(n28095), .n28094(n28094), .n28093(n28093), .n28092(n28092), 
         .n4(n4_adj_5310), .n7(n7_adj_5175), .n28091(n28091), .n27804(n27804), 
         .n28090(n28090), .n28089(n28089), .n28088(n28088), .n28545(n28545), 
         .\Kp[3] (Kp[3]), .n28544(n28544), .\Kp[4] (Kp[4]), .n28534(n28534), 
         .\Kp[5] (Kp[5]), .n28516(n28516), .n28515(n28515), .n28514(n28514), 
         .n28513(n28513), .n28512(n28512), .n28511(n28511), .n28510(n28510), 
         .n28509(n28509), .n28452(n28452), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .n28451(n28451), .n28450(n28450), .n28449(n28449), .n28448(n28448), 
         .n28447(n28447), .n28446(n28446), .n28445(n28445), .n28438(n28438), 
         .n28437(n28437), .n28433(n28433), .n28432(n28432), .n28431(n28431), 
         .n28430(n28430), .n28429(n28429), .n28428(n28428), .n28426(n28426), 
         .n28425(n28425), .n28424(n28424), .n28423(n28423), .n28422(n28422), 
         .n28421(n28421), .n28420(n28420), .n28416(n28416), .\Kp[6] (Kp[6]), 
         .n28415(n28415), .n28414(n28414), .n28413(n28413), .n28412(n28412), 
         .n28411(n28411), .n28410(n28410), .n28409(n28409), .n28408(n28408), 
         .n28407(n28407), .\Kp[7] (Kp[7]), .n28406(n28406), .\Kp[8] (Kp[8]), 
         .n28405(n28405), .\Kp[9] (Kp[9]), .n28404(n28404), .\Kp[10] (Kp[10]), 
         .n28403(n28403), .\Kp[11] (Kp[11]), .n28402(n28402), .\Kp[12] (Kp[12]), 
         .n28401(n28401), .\Kp[13] (Kp[13]), .n28400(n28400), .\Kp[14] (Kp[14]), 
         .n28399(n28399), .\Kp[15] (Kp[15]), .n28398(n28398), .\Ki[1] (Ki[1]), 
         .n28397(n28397), .\Ki[2] (Ki[2]), .n28396(n28396), .\Ki[3] (Ki[3]), 
         .n28395(n28395), .\Ki[4] (Ki[4]), .n28394(n28394), .\Ki[5] (Ki[5]), 
         .n28393(n28393), .\Ki[6] (Ki[6]), .n28392(n28392), .\Ki[7] (Ki[7]), 
         .n28391(n28391), .\Ki[8] (Ki[8]), .n28390(n28390), .\Ki[9] (Ki[9]), 
         .n28389(n28389), .\Ki[10] (Ki[10]), .n28388(n28388), .\Ki[11] (Ki[11]), 
         .n28387(n28387), .\Ki[12] (Ki[12]), .n28386(n28386), .\Ki[13] (Ki[13]), 
         .n28385(n28385), .\Ki[14] (Ki[14]), .n28384(n28384), .\Ki[15] (Ki[15]), 
         .n28383(n28383), .n28382(n28382), .n28381(n28381), .n28380(n28380), 
         .n28379(n28379), .n28378(n28378), .n28377(n28377), .n28373(n28373), 
         .n28361(n28361), .n28360(n28360), .n28359(n28359), .n28358(n28358), 
         .n28357(n28357), .n28356(n28356), .n28355(n28355), .n28354(n28354), 
         .n28353(n28353), .n28352(n28352), .n28351(n28351), .n28350(n28350), 
         .n28349(n28349), .n28348(n28348), .n28347(n28347), .n28346(n28346), 
         .n28345(n28345), .n28344(n28344), .n28343(n28343), .n28342(n28342), 
         .n28341(n28341), .n28340(n28340), .n28339(n28339), .n28338(n28338), 
         .n28337(n28337), .n28336(n28336), .n28335(n28335), .n28329(n28329), 
         .n28328(n28328), .n28327(n28327), .n28326(n28326), .n28325(n28325), 
         .n28324(n28324), .n28323(n28323), .n28322(n28322), .n28321(n28321), 
         .n28320(n28320), .n28319(n28319), .n28318(n28318), .n28317(n28317), 
         .n28316(n28316), .n28315(n28315), .n28314(n28314), .n28313(n28313), 
         .n28312(n28312), .n28311(n28311), .n28310(n28310), .n28309(n28309), 
         .n28308(n28308), .n28307(n28307), .n28306(n28306), .n28305(n28305), 
         .n28304(n28304), .n28303(n28303), .n28302(n28302), .n28301(n28301), 
         .n28300(n28300), .n28299(n28299), .n28298(n28298), .n28297(n28297), 
         .n42822(n42822), .n28296(n28296), .n28295(n28295), .n28294(n28294), 
         .n28293(n28293), .n28292(n28292), .n28291(n28291), .n28290(n28290), 
         .n28289(n28289), .n28288(n28288), .n28287(n28287), .n28286(n28286), 
         .n28285(n28285), .n28284(n28284), .n28283(n28283), .n28282(n28282), 
         .n28281(n28281), .n28280(n28280), .n28279(n28279), .n28278(n28278), 
         .n28277(n28277), .n28276(n28276), .n28275(n28275), .n28274(n28274), 
         .n28273(n28273), .n28272(n28272), .n28271(n28271), .n28270(n28270), 
         .n28269(n28269), .n28268(n28268), .n28267(n28267), .n28266(n28266), 
         .n28262(n28262), .n28261(n28261), .n28260(n28260), .n28258(n28258), 
         .n28257(n28257), .n42836(n42836), .n28256(n28256), .n28255(n28255), 
         .n28254(n28254), .n28253(n28253), .n28252(n28252), .n28251(n28251), 
         .n42843(n42843), .n28250(n28250), .n28249(n28249), .n28248(n28248), 
         .n28247(n28247), .n28246(n28246), .n28245(n28245), .n28243(n28243), 
         .n28242(n28242), .n28241(n28241), .n28240(n28240), .n28239(n28239), 
         .n28087(n28087), .n28238(n28238), .n28237(n28237), .n28236(n28236), 
         .n28235(n28235), .n43608(n43608), .n42830(n42830), .n23568(n23568), 
         .\state[0] (state_adj_5401[0]), .\state[3] (state_adj_5401[3]), 
         .\state[2] (state_adj_5401[2]), .n7233(n7233), .\r_SM_Main_2__N_3613[1] (r_SM_Main_2__N_3613[1]), 
         .r_SM_Main({r_SM_Main_adj_5388}), .n18940(n18940), .\r_Bit_Index[0] (r_Bit_Index_adj_5390[0]), 
         .tx_o(tx_o), .n27763(n27763), .n28054(n28054), .VCC_net(VCC_net), 
         .n48986(n48986), .n28365(n28365), .n28159(n28159), .n4_adj_10(n4_adj_5177), 
         .tx_enable(tx_enable), .\r_Bit_Index[0]_adj_11 (r_Bit_Index[0]), 
         .n27767(n27767), .r_SM_Main_adj_18({r_SM_Main}), .n28056(n28056), 
         .\r_SM_Main_2__N_3542[2] (r_SM_Main_2__N_3542[2]), .r_Rx_Data(r_Rx_Data), 
         .n26339(n26339), .n26334(n26334), .n33899(n33899), .RX_N_10(RX_N_10), 
         .n28368(n28368), .n42422(n42422), .n28142(n28142), .n28141(n28141), 
         .n28140(n28140), .n28139(n28139), .n28138(n28138), .n28128(n28128), 
         .n28127(n28127), .n42722(n42722), .n4_adj_15(n4_adj_5223), .n4_adj_16(n4_adj_5210), 
         .n4_adj_17(n4), .n28372(n28372)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(238[8] 261[4])
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1742 (.I0(n1728), .I1(n1726), .I2(n1727), .I3(GND_net), 
            .O(n45512));
    defparam i1_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i14579_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n23568), .I3(GND_net), .O(n28090));   // verilog/coms.v(127[12] 300[6])
    defparam i14579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5193));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21163_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n34672));
    defparam i21163_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n1723), .I1(n1724), .I2(n45512), .I3(n1725), 
            .O(n45518));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5194));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5195));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1744 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n45738));
    defparam i1_2_lut_adj_1744.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n45738), .I1(n1722), .I2(n45518), .I3(n34672), 
            .O(n45522));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'hfefc;
    SB_LUT4 i33194_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n45522), 
            .O(n1752));
    defparam i33194_4_lut.LUT_INIT = 16'h0001;
    \grp_debouncer(3,1000)  debounce (.reg_B({reg_B}), .CLK_c(CLK_c), .n45341(n45341), 
            .GND_net(GND_net), .data_i({hall1, hall2, hall3}), .VCC_net(VCC_net), 
            .n28107(n28107), .data_o({h1, h2, h3}), .n28529(n28529), 
            .n28419(n28419));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    SB_LUT4 i33306_4_lut (.I0(n1026), .I1(n43826), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i33306_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i20365_1_lut_2_lut (.I0(n23755), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n1964));
    defparam i20365_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1997_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1195), .I3(n26226), .O(n6976));   // verilog/TinyFPGA_B.v(360[5] 384[12])
    defparam i1997_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n27636), 
            .I3(rx_data_ready), .O(n42422));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n27636));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5295));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    EEPROM eeprom (.\state[0] (state_adj_5373[0]), .GND_net(GND_net), .read(read), 
           .\state[1] (state_adj_5373[1]), .\state[3] (state_adj_5401[3]), 
           .\state[0]_adj_6 (state_adj_5401[0]), .CLK_c(CLK_c), .\state[2] (state_adj_5401[2]), 
           .n5614({n5615}), .n28155(n28155), .rw(rw), .n42504(n42504), 
           .data_ready(data_ready), .n122(n122_adj_5176), .n10(n10_adj_5275), 
           .\state_7__N_4103[3] (state_7__N_4103[3]), .n7233(n7233), .\saved_addr[0] (saved_addr[0]), 
           .sda_enable(sda_enable), .VCC_net(VCC_net), .\state_7__N_4087[0] (state_7__N_4087[0]), 
           .scl_enable(scl_enable), .scl(scl), .sda_out(sda_out), .n28135(n28135), 
           .data({data}), .n28134(n28134), .n28133(n28133), .n28132(n28132), 
           .n28131(n28131), .n28130(n28130), .n28129(n28129), .n4(n4_adj_5232), 
           .n4_adj_7(n4_adj_5161), .n33869(n33869), .n28259(n28259), .n28244(n28244), 
           .n26367(n26367), .n26372(n26372)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(387[10] 398[6])
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095_adj_5255), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(1,500000)  quad_counter1 (.b_prev(b_prev_adj_5209), 
            .GND_net(GND_net), .a_new({a_new_adj_5349[1], Open_29}), .direction_N_3907(direction_N_3907_adj_5211), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1668(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .encoder1_position({encoder1_position}), .VCC_net(VCC_net), 
            .n28417(n28417), .n1673(n1673)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(294[57] 301[6])
    SB_LUT4 i5366_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_403));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i5366_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i5368_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_412));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i5368_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1039_rep_48_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1039_rep_48_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5294));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094_adj_5254), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .GND_net(GND_net), 
            .state_7__N_4293(state_7__N_4293), .\data[15] (data_adj_5377[15]), 
            .n44589(n44589), .n9(n9_adj_5230), .CLK_c(CLK_c), .n11(n11_adj_5231), 
            .VCC_net(VCC_net), .n5(n5_adj_5212), .n5_adj_1(n5_adj_5207), 
            .n33894(n33894), .n28153(n28153), .current({current}), .n28623(n28623), 
            .n28622(n28622), .n28621(n28621), .n28620(n28620), .n28619(n28619), 
            .n28618(n28618), .n28617(n28617), .n28616(n28616), .n28615(n28615), 
            .n28614(n28614), .n28613(n28613), .n28612(n28612), .n28125(n28125), 
            .n28124(n28124), .\data[12] (data_adj_5377[12]), .n28123(n28123), 
            .\data[11] (data_adj_5377[11]), .n28122(n28122), .\data[10] (data_adj_5377[10]), 
            .n28121(n28121), .\data[9] (data_adj_5377[9]), .n28120(n28120), 
            .\data[8] (data_adj_5377[8]), .n28119(n28119), .\data[7] (data_adj_5377[7]), 
            .n28118(n28118), .\data[6] (data_adj_5377[6]), .n28117(n28117), 
            .\data[5] (data_adj_5377[5]), .n28116(n28116), .\data[4] (data_adj_5377[4]), 
            .n28115(n28115), .\data[3] (data_adj_5377[3]), .n28114(n28114), 
            .\data[2] (data_adj_5377[2]), .n28113(n28113), .\data[1] (data_adj_5377[1]), 
            .n26390(n26390), .n26377(n26377), .n26385(n26385), .n26380(n26380), 
            .n28427(n28427), .\data[0] (data_adj_5377[0])) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(400[11] 406[4])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5293));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n42722));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5292));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i1_3_lut_4_lut (.I0(n26211), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5291));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21175_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n34684));
    defparam i21175_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1746 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n45636));
    defparam i1_3_lut_adj_1746.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632_adj_5263));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_5242), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n941));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5290));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5289));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .pwm_setpoint({pwm_setpoint}), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (\neo_pixel_transmitter.done , 
            CLK_c, \neo_pixel_transmitter.t0 , GND_net, \state_3__N_528[1] , 
            start, LED_c, \state[1] , n44588, timer, VCC_net, neopxl_color, 
            n28137, n27713, n43584, n41744, n28096, n14, n28577, 
            n28576, n28575, n28574, n28573, n28572, n28571, n28570, 
            n28569, n28568, n28567, n28566, n28565, n28564, n28563, 
            n28562, n28561, n28560, n28559, n28558, n28557, n28556, 
            n28555, n28554, n28553, n28552, n28551, n28550, n28549, 
            n28548, n28547, \neo_pixel_transmitter.done_N_742 , NEOPXL_c, 
            n47171) /* synthesis syn_module_defined=1 */ ;
    output \neo_pixel_transmitter.done ;
    input CLK_c;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    output \state_3__N_528[1] ;
    output start;
    input LED_c;
    output \state[1] ;
    output n44588;
    output [31:0]timer;
    input VCC_net;
    input [23:0]neopxl_color;
    input n28137;
    output n27713;
    output n43584;
    input n41744;
    input n28096;
    output n14;
    input n28577;
    input n28576;
    input n28575;
    input n28574;
    input n28573;
    input n28572;
    input n28571;
    input n28570;
    input n28569;
    input n28568;
    input n28567;
    input n28566;
    input n28565;
    input n28564;
    input n28563;
    input n28562;
    input n28561;
    input n28560;
    input n28559;
    input n28558;
    input n28557;
    input n28556;
    input n28555;
    input n28554;
    input n28553;
    input n28552;
    input n28551;
    input n28550;
    input n28549;
    input n28548;
    input n28547;
    input \neo_pixel_transmitter.done_N_742 ;
    output NEOPXL_c;
    output n47171;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire \neo_pixel_transmitter.done_N_736 , n45343;
    wire [31:0]n1;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    wire [31:0]color_bit_N_722;
    wire [31:0]n282;
    
    wire n27566, n27970, n28, n26, n27, n25, n16_adj_5148, n22_adj_5149, 
        n45253, n20_adj_5150, n24;
    wire [31:0]one_wire_N_679;
    
    wire n4_adj_5151, n39761, n26356, n4_adj_5152, n46094, n46100, 
        n26417, n26235, n1977, n34471, n6921, n47235, n43560, 
        n44621, n44620, n34520, n43780, n91, n43766, n42775, n42715;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n27587, n38333, n46088, n38332, n46086;
    wire [31:0]n133;
    
    wire n38175, n38953, n38952, n38951, n38950, n38949, n38948, 
        n38947, n38946, n38945, n38944, n38943, n38942, n38941, 
        n38940, n38939, n38938, n38937, n38936, n38935, n38934, 
        n38933, n38932, n38931, n38930, n38929, n38928, n38174, 
        n38927, n38926, n38925, n38924, n38923, n46358, n46359, 
        n38173, n38331, n46084, n46365, n46364, n38330, n46082, 
        n38329, n46080, n38172, n38328, n46078, n38327, n46076, 
        n38326, n46074, n38325, n46072, n38171, n38324, n46070, 
        n38323, n46068, n38170, n38322, n46066, n38169, n38168, 
        n38321, n46064, n38320, n46062, n38167, n38166, n38319, 
        n46060, n38165, n38318, n46058, n38164, n38163, n38317, 
        n46056, n48930, n48933, n38316, n46054, n38315, n46052, 
        n38314, n38162, n38313, n48879, n47821, n34432, n40277, 
        n48843, n47897, n48789, n47241;
    wire [3:0]state_3__N_528;
    
    wire n38312, n48840, n46421, n46422, n38161, n38160, n38311, 
        n38159, n46329, n46328, n34542, n38158, n47169, n38310, 
        n38309, n38308, n38307, n38306, n38157, n42814, n38305, 
        n38304, n38303, n38156, n48876, n38155, n43535, n1991, 
        n38154, n38153, n38152, n38151, n38150, n38149, n38148, 
        n38147, n38146, n38145, n48786, n44917, n12_adj_5159, n11_adj_5160, 
        n103;
    
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n45343), .D(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_722[1]));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n27566), .D(n282[1]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n27566), .D(n282[2]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n27566), .D(n282[3]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n27566), .D(n282[4]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n27566), .D(n282[5]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i12_4_lut (.I0(bit_ctr[12]), .I1(bit_ctr[23]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[20]), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n27566), .D(n282[6]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n27566), .D(n282[7]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n27566), .D(n282[8]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n27566), .D(n282[9]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n27566), 
            .D(n282[10]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n27566), 
            .D(n282[11]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n27566), 
            .D(n282[12]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n27566), 
            .D(n282[13]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n27566), 
            .D(n282[14]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n27566), 
            .D(n282[15]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n27566), 
            .D(n282[16]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n27566), 
            .D(n282[17]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n27566), 
            .D(n282[18]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n27566), 
            .D(n282[19]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i10_4_lut (.I0(bit_ctr[25]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n27566), 
            .D(n282[20]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n27566), 
            .D(n282[21]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n27566), 
            .D(n282[22]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n27566), 
            .D(n282[23]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n27566), 
            .D(n282[24]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n27566), 
            .D(n282[25]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n27566), 
            .D(n282[26]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n27566), 
            .D(n282[27]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n27566), 
            .D(n282[28]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n27566), 
            .D(n282[29]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n27566), 
            .D(n282[30]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n27566), 
            .D(n282[31]), .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i11_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[31]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[21]), .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(bit_ctr[22]), .I1(bit_ctr[5]), .I2(bit_ctr[17]), 
            .I3(bit_ctr[14]), .O(n25));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_5148));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1565 (.I0(bit_ctr[9]), .I1(bit_ctr[27]), .I2(bit_ctr[10]), 
            .I3(bit_ctr[15]), .O(n22_adj_5149));
    defparam i9_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n45253));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut (.I0(bit_ctr[26]), .I1(bit_ctr[3]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n20_adj_5150));
    defparam i7_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i11_4_lut_adj_1566 (.I0(n45253), .I1(n22_adj_5149), .I2(n16_adj_5148), 
            .I3(bit_ctr[11]), .O(n24));
    defparam i11_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1567 (.I0(bit_ctr[18]), .I1(n24), .I2(n20_adj_5150), 
            .I3(bit_ctr[8]), .O(\state_3__N_528[1] ));
    defparam i12_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(one_wire_N_679[2]), .I1(n4_adj_5151), .I2(GND_net), 
            .I3(GND_net), .O(n39761));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n26356));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5152));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1570 (.I0(one_wire_N_679[5]), .I1(one_wire_N_679[4]), 
            .I2(GND_net), .I3(GND_net), .O(n46094));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1570.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[7]), .I2(one_wire_N_679[6]), 
            .I3(n46094), .O(n46100));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(one_wire_N_679[10]), .I1(n26417), .I2(one_wire_N_679[9]), 
            .I3(n46100), .O(n26235));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i495_2_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1977));   // verilog/neopixel.v(40[18] 45[12])
    defparam i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4557_4_lut (.I0(n34471), .I1(n1977), .I2(\state[1] ), .I3(n26356), 
            .O(n6921));
    defparam i4557_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i32284_3_lut (.I0(n39761), .I1(n26356), .I2(n26235), .I3(GND_net), 
            .O(n47235));
    defparam i32284_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(\state[1] ), .I1(n26235), .I2(\neo_pixel_transmitter.done ), 
            .I3(n43560), .O(n44621));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'hfafb;
    SB_LUT4 i1_4_lut_adj_1573 (.I0(n44620), .I1(start), .I2(\state[1] ), 
            .I3(n44621), .O(n44588));
    defparam i1_4_lut_adj_1573.LUT_INIT = 16'ha280;
    SB_LUT4 i116_4_lut (.I0(n34520), .I1(n43780), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n91));
    defparam i116_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(n43766), .I1(n4_adj_5152), .I2(n39761), 
            .I3(n42775), .O(n42715));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'h1511;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n26417), .I1(state[0]), .I2(n42715), 
            .I3(n91), .O(n27587));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'h5150;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n46088), .I1(timer[31]), .I2(n1[31]), 
            .I3(n38333), .O(n26417)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n46086), .I1(timer[30]), .I2(n1[30]), 
            .I3(n38332), .O(n46088)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_DFF timer_2189__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n38175), .O(n282[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2189_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n38953), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2189_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n38952), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_32 (.CI(n38952), .I0(GND_net), .I1(timer[30]), 
            .CO(n38953));
    SB_LUT4 timer_2189_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n38951), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_31 (.CI(n38951), .I0(GND_net), .I1(timer[29]), 
            .CO(n38952));
    SB_LUT4 timer_2189_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n38950), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_30 (.CI(n38950), .I0(GND_net), .I1(timer[28]), 
            .CO(n38951));
    SB_LUT4 timer_2189_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n38949), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_29 (.CI(n38949), .I0(GND_net), .I1(timer[27]), 
            .CO(n38950));
    SB_LUT4 timer_2189_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n38948), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_28 (.CI(n38948), .I0(GND_net), .I1(timer[26]), 
            .CO(n38949));
    SB_LUT4 timer_2189_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n38947), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_27 (.CI(n38947), .I0(GND_net), .I1(timer[25]), 
            .CO(n38948));
    SB_LUT4 timer_2189_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n38946), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_26 (.CI(n38946), .I0(GND_net), .I1(timer[24]), 
            .CO(n38947));
    SB_LUT4 timer_2189_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n38945), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_25 (.CI(n38945), .I0(GND_net), .I1(timer[23]), 
            .CO(n38946));
    SB_LUT4 timer_2189_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n38944), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_24 (.CI(n38944), .I0(GND_net), .I1(timer[22]), 
            .CO(n38945));
    SB_LUT4 timer_2189_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n38943), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_23 (.CI(n38943), .I0(GND_net), .I1(timer[21]), 
            .CO(n38944));
    SB_LUT4 timer_2189_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n38942), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_22 (.CI(n38942), .I0(GND_net), .I1(timer[20]), 
            .CO(n38943));
    SB_LUT4 timer_2189_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n38941), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_32 (.CI(n38332), .I0(timer[30]), .I1(n1[30]), 
            .CO(n38333));
    SB_CARRY timer_2189_add_4_21 (.CI(n38941), .I0(GND_net), .I1(timer[19]), 
            .CO(n38942));
    SB_LUT4 timer_2189_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n38940), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_20 (.CI(n38940), .I0(GND_net), .I1(timer[18]), 
            .CO(n38941));
    SB_LUT4 timer_2189_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n38939), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_19 (.CI(n38939), .I0(GND_net), .I1(timer[17]), 
            .CO(n38940));
    SB_LUT4 timer_2189_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n38938), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_18 (.CI(n38938), .I0(GND_net), .I1(timer[16]), 
            .CO(n38939));
    SB_LUT4 timer_2189_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n38937), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_17 (.CI(n38937), .I0(GND_net), .I1(timer[15]), 
            .CO(n38938));
    SB_LUT4 timer_2189_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n38936), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_16 (.CI(n38936), .I0(GND_net), .I1(timer[14]), 
            .CO(n38937));
    SB_LUT4 timer_2189_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n38935), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_15 (.CI(n38935), .I0(GND_net), .I1(timer[13]), 
            .CO(n38936));
    SB_LUT4 timer_2189_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n38934), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_14 (.CI(n38934), .I0(GND_net), .I1(timer[12]), 
            .CO(n38935));
    SB_LUT4 timer_2189_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n38933), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_13 (.CI(n38933), .I0(GND_net), .I1(timer[11]), 
            .CO(n38934));
    SB_LUT4 timer_2189_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n38932), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_12 (.CI(n38932), .I0(GND_net), .I1(timer[10]), 
            .CO(n38933));
    SB_LUT4 timer_2189_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n38931), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_11 (.CI(n38931), .I0(GND_net), .I1(timer[9]), 
            .CO(n38932));
    SB_LUT4 timer_2189_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n38930), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_10 (.CI(n38930), .I0(GND_net), .I1(timer[8]), 
            .CO(n38931));
    SB_LUT4 timer_2189_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n38929), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_9 (.CI(n38929), .I0(GND_net), .I1(timer[7]), 
            .CO(n38930));
    SB_LUT4 timer_2189_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n38928), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n38174), .O(n282[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_8 (.CI(n38928), .I0(GND_net), .I1(timer[6]), 
            .CO(n38929));
    SB_LUT4 timer_2189_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n38927), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_7 (.CI(n38927), .I0(GND_net), .I1(timer[5]), 
            .CO(n38928));
    SB_LUT4 timer_2189_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n38926), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_6 (.CI(n38926), .I0(GND_net), .I1(timer[4]), 
            .CO(n38927));
    SB_LUT4 timer_2189_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n38925), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_5 (.CI(n38925), .I0(GND_net), .I1(timer[3]), 
            .CO(n38926));
    SB_LUT4 timer_2189_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n38924), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_4 (.CI(n38924), .I0(GND_net), .I1(timer[2]), 
            .CO(n38925));
    SB_LUT4 timer_2189_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n38923), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_3 (.CI(n38923), .I0(GND_net), .I1(timer[1]), 
            .CO(n38924));
    SB_LUT4 timer_2189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n38923));
    SB_LUT4 i31277_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46358));
    defparam i31277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31278_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46359));
    defparam i31278_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_32 (.CI(n38174), .I0(bit_ctr[30]), .I1(GND_net), .CO(n38175));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n38173), .O(n282[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_31_lut (.I0(n46084), .I1(timer[29]), .I2(n1[29]), 
            .I3(n38331), .O(n46086)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n38331), .I0(timer[29]), .I1(n1[29]), 
            .CO(n38332));
    SB_LUT4 i31284_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46365));
    defparam i31284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31283_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n46364));
    defparam i31283_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_31 (.CI(n38173), .I0(bit_ctr[29]), .I1(GND_net), .CO(n38174));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n46082), .I1(timer[28]), .I2(n1[28]), 
            .I3(n38330), .O(n46084)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n38330), .I0(timer[28]), .I1(n1[28]), 
            .CO(n38331));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n46080), .I1(timer[27]), .I2(n1[27]), 
            .I3(n38329), .O(n46082)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n38329), .I0(timer[27]), .I1(n1[27]), 
            .CO(n38330));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n38172), .O(n282[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_28_lut (.I0(n46078), .I1(timer[26]), .I2(n1[26]), 
            .I3(n38328), .O(n46080)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_28 (.CI(n38328), .I0(timer[26]), .I1(n1[26]), 
            .CO(n38329));
    SB_LUT4 sub_14_add_2_27_lut (.I0(n46076), .I1(timer[25]), .I2(n1[25]), 
            .I3(n38327), .O(n46078)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n38327), .I0(timer[25]), .I1(n1[25]), 
            .CO(n38328));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n46074), .I1(timer[24]), .I2(n1[24]), 
            .I3(n38326), .O(n46076)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_26 (.CI(n38326), .I0(timer[24]), .I1(n1[24]), 
            .CO(n38327));
    SB_CARRY add_21_30 (.CI(n38172), .I0(bit_ctr[28]), .I1(GND_net), .CO(n38173));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n46072), .I1(timer[23]), .I2(n1[23]), 
            .I3(n38325), .O(n46074)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n38171), .O(n282[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n38171), .I0(bit_ctr[27]), .I1(GND_net), .CO(n38172));
    SB_CARRY sub_14_add_2_25 (.CI(n38325), .I0(timer[23]), .I1(n1[23]), 
            .CO(n38326));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n46070), .I1(timer[22]), .I2(n1[22]), 
            .I3(n38324), .O(n46072)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n38324), .I0(timer[22]), .I1(n1[22]), 
            .CO(n38325));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n46068), .I1(timer[21]), .I2(n1[21]), 
            .I3(n38323), .O(n46070)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n38170), .O(n282[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_23 (.CI(n38323), .I0(timer[21]), .I1(n1[21]), 
            .CO(n38324));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n46066), .I1(timer[20]), .I2(n1[20]), 
            .I3(n38322), .O(n46068)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_28 (.CI(n38170), .I0(bit_ctr[26]), .I1(GND_net), .CO(n38171));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n38169), .O(n282[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n38169), .I0(bit_ctr[25]), .I1(GND_net), .CO(n38170));
    SB_CARRY sub_14_add_2_22 (.CI(n38322), .I0(timer[20]), .I1(n1[20]), 
            .CO(n38323));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n38168), .O(n282[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n46064), .I1(timer[19]), .I2(n1[19]), 
            .I3(n38321), .O(n46066)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n38321), .I0(timer[19]), .I1(n1[19]), 
            .CO(n38322));
    SB_CARRY add_21_26 (.CI(n38168), .I0(bit_ctr[24]), .I1(GND_net), .CO(n38169));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n46062), .I1(timer[18]), .I2(n1[18]), 
            .I3(n38320), .O(n46064)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_20 (.CI(n38320), .I0(timer[18]), .I1(n1[18]), 
            .CO(n38321));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n38167), .O(n282[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_25 (.CI(n38167), .I0(bit_ctr[23]), .I1(GND_net), .CO(n38168));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n38166), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n38166), .I0(bit_ctr[22]), .I1(GND_net), .CO(n38167));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n46060), .I1(timer[17]), .I2(n1[17]), 
            .I3(n38319), .O(n46062)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n38165), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_19 (.CI(n38319), .I0(timer[17]), .I1(n1[17]), 
            .CO(n38320));
    SB_CARRY add_21_23 (.CI(n38165), .I0(bit_ctr[21]), .I1(GND_net), .CO(n38166));
    SB_LUT4 sub_14_add_2_18_lut (.I0(n46058), .I1(timer[16]), .I2(n1[16]), 
            .I3(n38318), .O(n46060)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n38164), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n38164), .I0(bit_ctr[20]), .I1(GND_net), .CO(n38165));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n38163), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n38318), .I0(timer[16]), .I1(n1[16]), 
            .CO(n38319));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n46056), .I1(timer[15]), .I2(n1[15]), 
            .I3(n38317), .O(n46058)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_21 (.CI(n38163), .I0(bit_ctr[19]), .I1(GND_net), .CO(n38164));
    SB_LUT4 n48930_bdd_4_lut (.I0(n48930), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_722[1]), .O(n48933));
    defparam n48930_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY sub_14_add_2_17 (.CI(n38317), .I0(timer[15]), .I1(n1[15]), 
            .CO(n38318));
    SB_LUT4 sub_14_add_2_16_lut (.I0(n46054), .I1(timer[14]), .I2(n1[14]), 
            .I3(n38316), .O(n46056)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n38316), .I0(timer[14]), .I1(n1[14]), 
            .CO(n38317));
    SB_LUT4 sub_14_add_2_15_lut (.I0(n46052), .I1(timer[13]), .I2(n1[13]), 
            .I3(n38315), .O(n46054)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n38315), .I0(timer[13]), .I1(n1[13]), 
            .CO(n38316));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_679[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n38314), .O(n46052)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n38162), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n38314), .I0(timer[12]), .I1(n1[12]), 
            .CO(n38315));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n38313), .O(one_wire_N_679[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n38313), .I0(timer[11]), .I1(n1[11]), 
            .CO(n38314));
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n28137));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i32740_3_lut (.I0(n48879), .I1(n48933), .I2(color_bit_N_722[2]), 
            .I3(GND_net), .O(n47821));
    defparam i32740_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n34432), .I3(GND_net), 
            .O(n40277));
    defparam i1_3_lut.LUT_INIT = 16'h6a6a;
    SB_DFF timer_2189__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i32816_4_lut (.I0(n47821), .I1(n48843), .I2(bit_ctr[3]), .I3(n34432), 
            .O(n47897));   // verilog/neopixel.v(22[26:38])
    defparam i32816_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i32246_3_lut (.I0(n48789), .I1(bit_ctr[3]), .I2(n34432), .I3(GND_net), 
            .O(n47241));
    defparam i32246_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i20366_4_lut (.I0(n47241), .I1(\state_3__N_528[1] ), .I2(n47897), 
            .I3(n40277), .O(state_3__N_528[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i20366_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_21_20 (.CI(n38162), .I0(bit_ctr[18]), .I1(GND_net), .CO(n38163));
    SB_DFFESS state_i0 (.Q(state[0]), .C(CLK_c), .E(n27713), .D(state_3__N_528[0]), 
            .S(n43584));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n38312), .O(one_wire_N_679[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 color_bit_N_722_1__bdd_4_lut (.I0(color_bit_N_722[1]), .I1(n46364), 
            .I2(n46365), .I3(color_bit_N_722[2]), .O(n48840));
    defparam color_bit_N_722_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48840_bdd_4_lut (.I0(n48840), .I1(n46359), .I2(n46358), .I3(color_bit_N_722[2]), 
            .O(n48843));
    defparam n48840_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i31340_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n46421));
    defparam i31340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31341_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n46422));
    defparam i31341_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_12 (.CI(n38312), .I0(timer[10]), .I1(n1[10]), 
            .CO(n38313));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n38161), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n38161), .I0(bit_ctr[17]), .I1(GND_net), .CO(n38162));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n38160), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_18 (.CI(n38160), .I0(bit_ctr[16]), .I1(GND_net), .CO(n38161));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n38311), .O(one_wire_N_679[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n38159), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF start_103 (.Q(start), .C(CLK_c), .D(n41744));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n28096));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i31248_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n46329));
    defparam i31248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31247_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n46328));
    defparam i31247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21013_3_lut (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[10]), 
            .I2(one_wire_N_679[9]), .I3(GND_net), .O(n34520));
    defparam i21013_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i21034_2_lut (.I0(n34520), .I1(n26417), .I2(GND_net), .I3(GND_net), 
            .O(n34542));
    defparam i21034_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28568_4_lut (.I0(n26235), .I1(n39761), .I2(n4_adj_5152), 
            .I3(state[0]), .O(n14));   // verilog/neopixel.v(35[12] 117[6])
    defparam i28568_4_lut.LUT_INIT = 16'hfaee;
    SB_CARRY add_21_17 (.CI(n38159), .I0(bit_ctr[15]), .I1(GND_net), .CO(n38160));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n38158), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1576 (.I0(n14), .I1(n47169), .I2(\state[1] ), 
            .I3(n26356), .O(n43584));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1576.LUT_INIT = 16'h303a;
    SB_CARRY sub_14_add_2_11 (.CI(n38311), .I0(timer[9]), .I1(n1[9]), 
            .CO(n38312));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n38310), .O(one_wire_N_679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n38310), .I0(timer[8]), .I1(n1[8]), 
            .CO(n38311));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n38309), .O(one_wire_N_679[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n38309), .I0(timer[7]), .I1(n1[7]), .CO(n38310));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n38308), .O(one_wire_N_679[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n38308), .I0(timer[6]), .I1(n1[6]), .CO(n38309));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n38307), .O(one_wire_N_679[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n38307), .I0(timer[5]), .I1(n1[5]), .CO(n38308));
    SB_CARRY add_21_16 (.CI(n38158), .I0(bit_ctr[14]), .I1(GND_net), .CO(n38159));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n38306), .O(one_wire_N_679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n38157), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n38306), .I0(timer[4]), .I1(n1[4]), .CO(n38307));
    SB_LUT4 i1_3_lut_2_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n42814));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n38305), .O(one_wire_N_679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n38305), .I0(timer[3]), .I1(n1[3]), .CO(n38306));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n38304), .O(one_wire_N_679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n27566), .D(n282[0]), 
            .R(n27970));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_4 (.CI(n38304), .I0(timer[2]), .I1(n1[2]), .CO(n38305));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_679[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n38303), .O(n4_adj_5151)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_15 (.CI(n38157), .I0(bit_ctr[13]), .I1(GND_net), .CO(n38158));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n38156), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n38303), .I0(timer[1]), .I1(n1[1]), .CO(n38304));
    SB_LUT4 bit_ctr_0__bdd_4_lut_33821_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n48876));   // verilog/neopixel.v(19[6:15])
    defparam bit_ctr_0__bdd_4_lut_33821_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_CARRY add_21_14 (.CI(n38156), .I0(bit_ctr[12]), .I1(GND_net), .CO(n38157));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n38303));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n38155), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n38155), .I0(bit_ctr[11]), .I1(GND_net), .CO(n38156));
    SB_LUT4 i32434_2_lut_4_lut (.I0(n34520), .I1(n26417), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n47169));   // verilog/neopixel.v(35[12] 117[6])
    defparam i32434_2_lut_4_lut.LUT_INIT = 16'hfff1;
    SB_LUT4 i1_2_lut_3_lut (.I0(n14), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n43535));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i509_2_lut_3_lut (.I0(n34520), .I1(n26417), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n1991));   // verilog/neopixel.v(103[9] 111[12])
    defparam i509_2_lut_3_lut.LUT_INIT = 16'hf1f1;
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n38154), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_12 (.CI(n38154), .I0(bit_ctr[10]), .I1(GND_net), .CO(n38155));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n38153), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n48930));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_CARRY add_21_11 (.CI(n38153), .I0(bit_ctr[9]), .I1(GND_net), .CO(n38154));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n38152), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_10 (.CI(n38152), .I0(bit_ctr[8]), .I1(GND_net), .CO(n38153));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n38151), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n38151), .I0(bit_ctr[7]), .I1(GND_net), .CO(n38152));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n38150), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_8 (.CI(n38150), .I0(bit_ctr[6]), .I1(GND_net), .CO(n38151));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n38149), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_7 (.CI(n38149), .I0(bit_ctr[5]), .I1(GND_net), .CO(n38150));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n38148), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n38148), .I0(bit_ctr[4]), .I1(GND_net), .CO(n38149));
    SB_LUT4 i28758_2_lut_3_lut (.I0(n43766), .I1(one_wire_N_679[2]), .I2(n4_adj_5151), 
            .I3(GND_net), .O(n43780));
    defparam i28758_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n38147), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_5 (.CI(n38147), .I0(bit_ctr[3]), .I1(GND_net), .CO(n38148));
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n38146), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n38146), .I0(bit_ctr[2]), .I1(GND_net), .CO(n38147));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n38145), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n38145), .I0(bit_ctr[1]), .I1(GND_net), .CO(n38146));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n282[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n38145));
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[1] ), .I1(state[0]), .I2(n1991), 
            .I3(n43535), .O(n27713));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hdf8a;
    SB_LUT4 i33012_4_lut_4_lut (.I0(\state[1] ), .I1(state[0]), .I2(n6921), 
            .I3(n47235), .O(n27566));
    defparam i33012_4_lut_4_lut.LUT_INIT = 16'h0c1d;
    SB_LUT4 i1_3_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n14), .I3(\state[1] ), .O(n44620));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i23_3_lut_4_lut (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(n4_adj_5151), .I3(state[0]), .O(n43560));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'ha0ee;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n28577));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n28576));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n28575));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n28574));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n28573));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n28572));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n28571));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n28570));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n28569));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n28568));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n28567));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n28566));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n28565));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n28564));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n28563));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n28562));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n28561));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n28560));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n28559));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n28558));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n28557));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n28556));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n28555));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n28554));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n28553));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n28552));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n28551));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n28550));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n28549));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n28548));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n28547));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 color_bit_N_722_1__bdd_4_lut_33748 (.I0(color_bit_N_722[1]), .I1(n46328), 
            .I2(n46329), .I3(color_bit_N_722[2]), .O(n48786));
    defparam color_bit_N_722_1__bdd_4_lut_33748.LUT_INIT = 16'he4aa;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n48786_bdd_4_lut (.I0(n48786), .I1(n46422), .I2(n46421), .I3(color_bit_N_722[2]), 
            .O(n48789));
    defparam n48786_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i20928_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n34432));
    defparam i20928_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1577 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_722[2]));
    defparam i1_2_lut_3_lut_adj_1577.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1_2_lut_adj_1578 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n42775));
    defparam i1_2_lut_adj_1578.LUT_INIT = 16'h2222;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n27587), .D(\neo_pixel_transmitter.done_N_742 ), 
            .R(n44917));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 n48876_bdd_4_lut_4_lut (.I0(color_bit_N_722[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n48876), .O(n48879));   // verilog/neopixel.v(19[6:15])
    defparam n48876_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[5]), .I2(one_wire_N_679[6]), 
            .I3(one_wire_N_679[9]), .O(n12_adj_5159));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(one_wire_N_679[7]), .I1(one_wire_N_679[4]), .I2(one_wire_N_679[10]), 
            .I3(GND_net), .O(n11_adj_5160));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n34542), .I3(\state[1] ), .O(n44917));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n11_adj_5160), .I2(start), 
            .I3(n12_adj_5159), .O(n43766));
    defparam i2_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32289_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n34542), .I3(start), .O(n47171));
    defparam i32289_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(one_wire_N_679[2]), .I1(n42814), .I2(one_wire_N_679[3]), 
            .I3(n4_adj_5151), .O(n103));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'h45cd;
    SB_LUT4 i33000_3_lut (.I0(n43766), .I1(n103), .I2(n26417), .I3(GND_net), 
            .O(n45343));
    defparam i33000_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 mux_1255_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1255_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i2_2_lut_3_lut (.I0(n26235), .I1(one_wire_N_679[2]), .I2(one_wire_N_679[3]), 
            .I3(GND_net), .O(n34471));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1580 (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_528[1] ), .O(n27970));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut_adj_1580.LUT_INIT = 16'h8000;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Ki[4] , \Ki[5] , \Ki[1] , \Ki[6] , 
            \Ki[7] , \Ki[8] , \Kp[14] , \Kp[15] , \Ki[9] , IntegralLimit, 
            \Ki[10] , \Ki[11] , \Ki[0] , \Ki[2] , \Ki[3] , \Ki[12] , 
            \Kp[1] , \Kp[0] , \Kp[2] , \Ki[13] , \Kp[3] , \Kp[4] , 
            \Ki[14] , \Ki[15] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , 
            \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , duty, 
            clk32MHz, VCC_net, setpoint, motor_state, PWMLimit) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[1] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Ki[9] ;
    input [23:0]IntegralLimit;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[12] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Ki[13] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    output [23:0]duty;
    input clk32MHz;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    input [23:0]PWMLimit;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n13, n10, n12, n35, n30;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3672 ;
    
    wire n299, n13_adj_4726, n39161;
    wire [5:0]n18513;
    
    wire n195, n39162, n372, n33, n31, n29, n47462, n47458, 
        n47454, n48005, n18, n38034, n4, n44653;
    wire [6:0]n18416;
    
    wire n53, n122, n47918, n47607, n48053, n37, n48054, n39, 
        n48040, n7, n6, n21, n47919, n23, n47920, n445, n518, 
        n591;
    wire [23:0]n1;
    
    wire n1044, n1117, n664, n320, n43, n25, n47468, n47445;
    wire [12:0]n16869;
    wire [11:0]n17233;
    
    wire n980, n39160;
    wire [23:0]n1_adj_5146;
    
    wire n24, n8, n45, n47442, n47805, n393, n737, n47605, n38370, 
        n38371, n41, n48023, n47448, n907, n39159, n47959, n27, 
        n38369, n47613, n810, n119, n50, n192, n48015, n4_adj_4729;
    wire [23:0]duty_23__N_3772;
    wire [47:0]n106;
    wire [47:0]n155;
    
    wire n38257, n38258, n834, n39158, n38368, n761, n39157, n466, 
        n47925, n265, n883, n539, n338, n688, n39156, n47926, 
        n49304, n47739, n47493, n125, n49328, n56, n198;
    wire [16:0]n15136;
    wire [15:0]n15713;
    
    wire n895, n39469, n30_adj_4732, n10_adj_4733, n47491, n48003, 
        n47597, n48051, n48052, n48042, n49295, n48047, n47484, 
        n47595, n47803, n49291, n47482, n47957, n47603;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3723 ;
    
    wire \PID_CONTROLLER.integral_23__N_3722 , n48013, n341, n381, \PID_CONTROLLER.integral_23__N_3720 , 
        n414, n113, n44, n956, n411, n271, n344, n615, n39155, 
        n39321;
    wire [19:0]n12529;
    
    wire n39322;
    wire [20:0]n11605;
    
    wire n39320, n542, n39154, n39176, n831, n39177, n39470, n469, 
        n39153, n396, n39152, n822, n39468;
    wire [13:0]n16449;
    
    wire n758, n39175, n749, n39467, n676, n39466, n38367, n603, 
        n39465, n323, n39151, n530, n39464, n685, n39174, n612, 
        n250, n39150, n177, n39149, n35_adj_4736, n104;
    wire [10:0]n17545;
    
    wire n910, n39148, n38366, n837, n39147, n764, n39146, n691, 
        n39145, n618, n39144, n545, n39143, n1029, n487, n560, 
        n186, n39319, n457, n39463, n384, n39462, n311, n39461, 
        n104_adj_4737, n238, n39460, n165, n39459, n23_adj_4738, 
        n92, n35_adj_4740, n39318;
    wire [7:0]n18209;
    wire [6:0]n18353;
    
    wire n630, n39458, n39317, n454, n527, n177_adj_4741, n98, 
        n29_adj_4744, n101, n32, n174, n1111, n247;
    wire [23:0]n4236;
    
    wire n320_adj_4745, n393_adj_4746, n165_adj_4747, n110, n417, 
        n6_adj_4749;
    wire [3:0]n18633;
    wire [4:0]n18584;
    
    wire n600, n41_adj_4750, n183, n472, n39142, n204, n557, n39457, 
        n399, n39141, n238_adj_4752;
    wire [1:0]n18681;
    
    wire n256, n311_adj_4754, n250_adj_4755, n259, n673, n384_adj_4756, 
        n332, n326, n39140, n1102, n39316, n484, n39456, n171, 
        n329, n405, n131, n244, n323_adj_4757, n396_adj_4758, n62, 
        n466_adj_4760, n746, n86, n478, n469_adj_4761, n17_adj_4762, 
        n317, n159, n551, n539_adj_4763, n253, n39139, n232, n624, 
        n4_adj_4764;
    wire [2:0]n18664;
    
    wire n490, n390, n697, n12_adj_4765, n463, n542_adj_4766, n8_adj_4767, 
        n11_adj_4768, n6_adj_4769, n37861, n18_adj_4770, n13_adj_4771, 
        n4_adj_4772, n44771, n305, n770, n612_adj_4773, n378, n83, 
        n14_adj_4774, n685_adj_4775, n451, n524, n597, n156, n229, 
        n180, n39138, n536, n107, n38, n19_adj_4777, n38365, n39137, 
        n39136, n758_adj_4778, n38256, n39315, n39173, n402, n670, 
        n341_adj_4780, n39135, n302, n39134, n39455, n39314, n609, 
        n39133, n682, n375, n448, n755, n828, n521, n594, n901, 
        n17_adj_4781, n38364, n39454, n39172, n819, n615_adj_4782, 
        n39313, n39453, n39171, n39452, n39312, n39311, n39170, 
        n457_adj_4783, n15_adj_4784, n38363, n39169, n39310;
    wire [14:0]n16224;
    
    wire n39451, n39450, n39449, n667, n39309, n39308, n39307, 
        n39306, n475, n39305, n974, n688_adj_4785, n740, n1047, 
        n548, n1120, n892, n113_adj_4786, n831_adj_4787, n813, n44_adj_4788, 
        n886, n971, n39448, n95, n26_adj_4789, n965, n168, n761_adj_4790, 
        n834_adj_4791, n530_adj_4792, n186_adj_4793, n247_adj_4794, 
        n39168, n226, n39304, n174_adj_4795, n39167, n898, n39447, 
        n259_adj_4796, n603_adj_4797, n621, n332_adj_4798, n405_adj_4799, 
        n38362, n38255;
    wire [23:0]duty_23__N_3648;
    
    wire n825, n39446, n153, n39303, n676_adj_4801, n32_adj_4802, 
        n101_adj_4803, n11_adj_4804, n80, n694, n38254, n560_adj_4805, 
        n39166, n487_adj_4806, n39165, n478_adj_4807, n752, n39445, 
        n749_adj_4808, n551_adj_4809, n822_adj_4810, n767, n11_adj_4811, 
        n38361, n907_adj_4812, n9_adj_4813, n38360, n679, n39444, 
        n624_adj_4816, n1038, n743;
    wire [18:0]n13369;
    
    wire n39302, n980_adj_4817, n606, n39443;
    wire [9:0]n17809;
    
    wire n840, n39101, n767_adj_4818, n39100, n39301, n414_adj_4819, 
        n39164, n895_adj_4820, n533, n39442, n840_adj_4821, n39300, 
        n39299, n38359, n694_adj_4822, n39099, n460, n39441, n38253, 
        n621_adj_4823, n39098, n387, n39440, n548_adj_4824, n39097, 
        n475_adj_4825, n39096, n402_adj_4826, n39095, n329_adj_4827, 
        n39094, n256_adj_4828, n39093, n697_adj_4829, n770_adj_4830, 
        n968, n107_adj_4831, n183_adj_4832, n39092, n38_adj_4833, 
        n1041, n1114, n180_adj_4834, n253_adj_4835, n326_adj_4836, 
        n399_adj_4837, n5_adj_4838, n38358, n3_adj_4840, n38357, n41_adj_4842, 
        n110_adj_4843, n116, n47, n39298, n314, n39439, n1105, 
        n39297, n189_adj_4845, n1032, n39296, n472_adj_4846, n262, 
        n959, n39295, n241, n39438, n545_adj_4847, n335, n618_adj_4848, 
        n408, n481, n554, n691_adj_4849, n627, n764_adj_4851, n700, 
        n38252, n38356, n38355, n38354, n38251, n38250, n39437, 
        n39294, n39293, n38353;
    wire [23:0]n257;
    
    wire n256_adj_4853;
    wire [23:0]duty_23__N_3747;
    
    wire duty_23__N_3771, n38352;
    wire [13:0]n16673;
    
    wire n39436, n38351, n38350, n39435, n39292, n38349, n39434, 
        n38348, n38347, n38346, n38345, n39291, n38249, n39433, 
        n39290, n38344, n968_adj_4859, n816, n39289, n889, n38343, 
        n39432, n38248, n38342, n904, n38341, n39431, n39288, 
        n38247, n39287, n39430, n39429, n39286, n39163, n38340, 
        n38339, n1041_adj_4862, n1114_adj_4863, n904_adj_4864, n38338, 
        n39428, n39285, n39284, n89, n20_adj_4866, n38337, n38246, 
        n77, n8_adj_4869, n38336;
    wire [9:0]n17929;
    wire [8:0]n18128;
    
    wire n39283, n39427, n39282, n38245, n39426, n162, n39281, 
        n38335, n38334, n38244, n39280, n39425, n150_adj_4874, n977, 
        n39279, n235, n38243, n39424, n39278, n837_adj_4876, n89_adj_4877, 
        n20_adj_4878, n910_adj_4879, n1050, n39423, n962, n98_adj_4881, 
        n38242, n39277, n29_adj_4883, n39276, n171_adj_4885, n223, 
        n308;
    wire [23:0]n1_adj_5147;
    
    wire n39275;
    wire [5:0]n18465;
    
    wire n39422, n39421, n39420;
    wire [17:0]n14129;
    
    wire n39274, n39273, n39419, n39272, n39271, n268_adj_4889, 
        n39418, n195_adj_4890, n39417, n53_adj_4891, n122_adj_4892, 
        n1108, n39270;
    wire [12:0]n17064;
    
    wire n1050_adj_4893, n39416, n977_adj_4894, n39415, n1035, n39269, 
        n39268, n39414, n39267, n39266, n244_adj_4895, n296, n39265, 
        n39413, n39264, n39412, n39263, n39262, n39261, n39411, 
        n39260, n39410, n381_adj_4897, n47440, n369, n454_adj_4901, 
        n6_adj_4902, n39259, n527_adj_4903, n39258, n39409, n600_adj_4904, 
        n673_adj_4905, n47406, n6_adj_4906, n746_adj_4907, n819_adj_4908, 
        n39257, n39408, n892_adj_4909, n965_adj_4910, n1038_adj_4911;
    wire [16:0]n14813;
    
    wire n39256, n1111_adj_4912, n317_adj_4913, n116_adj_4914, n47_adj_4915, 
        n189_adj_4916, n39407, n39255, n39254, n39406, n262_adj_4917, 
        n335_adj_4918, n408_adj_4919, n481_adj_4920, n39405, n39253, 
        n39404, n554_adj_4921, n627_adj_4922;
    wire [11:0]n17401;
    
    wire n39403, n39252, n39402, n39401, n39400, n39251, n39250, 
        n39399, n39398, n39249, n39397, n39396, n39248, n39395, 
        n39394, n39247, n162_adj_4923, n125_adj_4924, n56_adj_4925, 
        n198_adj_4926, n39393, n39246, n39392, n235_adj_4927, n39245, 
        n271_adj_4928, n39244, n39243, n490_adj_4929, n39391, n344_adj_4930;
    wire [4:0]n18549;
    
    wire n417_adj_4931, n39390, n308_adj_4932, n39242, n268_adj_4933, 
        n39389, n39388, n39241, n39387, n39240;
    wire [10:0]n17688;
    
    wire n39386, n39385, n442, n4_adj_4935;
    wire [3:0]n18609;
    
    wire n6_adj_4936;
    wire [7:0]n18289;
    
    wire n39239, n39384, n39238, n39383, n39237, n39236, n39235, 
        n39382, n39234, n39381, n39233, n39380, n39232, n39379, 
        n39378, n8_adj_4937, n37836;
    wire [1:0]n18673;
    
    wire n39377;
    wire [15:0]n15425;
    
    wire n39231, n39230;
    wire [2:0]n18649;
    
    wire n37877, n4_adj_4938, n39376, n39229, n39228, n47408, n47418, 
        n47310, n39227;
    wire [8:0]n18029;
    
    wire n38434, n47340, n38433, n39375, n39226, n38432, n39374, 
        n39225, n38431, n37918, n39224, n38430, n39373, n39223, 
        n38429, n38428, n39372, n39222, n38427, n38426, n39221, 
        n700_adj_4939, n86_adj_4940, n12_adj_4941, n17_adj_4942, n8_adj_4943, 
        n11_adj_4944, n6_adj_4945, n159_adj_4946, n39371, n232_adj_4947, 
        n39370, n305_adj_4948, n378_adj_4949, n39220, n451_adj_4950, 
        n524_adj_4951, n597_adj_4952, n670_adj_4953, n39369, n743_adj_4954, 
        n816_adj_4955, n889_adj_4956, n39368, n39219, n39218, n39367, 
        n39217, n39366;
    wire [0:0]n10081;
    wire [21:0]n10588;
    
    wire n39365, n39216, n38287, n38286, n23_adj_4957, n92_adj_4958;
    wire [14:0]n15969;
    
    wire n39215, n38285, n1117_adj_4959, n39214, n39364, n1044_adj_4960, 
        n39213, n962_adj_4961, n1035_adj_4962, n38284, n1108_adj_4963, 
        n38283, n971_adj_4964, n39212, n83_adj_4965, n14_adj_4966, 
        n38282, n156_adj_4967, n39363, n515, n39362, n898_adj_4969, 
        n39211, n229_adj_4970, n302_adj_4971, n39361, n375_adj_4973, 
        n390_adj_4974, n825_adj_4975, n39210, n39360, n752_adj_4976, 
        n39209, n588, n679_adj_4977, n39208, n39359, n448_adj_4979, 
        n39358, n38281, n606_adj_4980, n39207, n521_adj_4981, n661, 
        n1096, n39357, n533_adj_4982, n39206, n38280, n594_adj_4983;
    wire [0:0]n10612;
    wire [21:0]n11119;
    
    wire n39599, n39598, n39597, n39596, n39595, n39594, n39593, 
        n39592, n1023, n39356, n460_adj_4984, n39205, n1096_adj_4985, 
        n39591, n1023_adj_4986, n39590, n950, n39589, n877, n39588, 
        n387_adj_4988, n39204, n667_adj_4989, n38279, n804, n39587, 
        n731, n39586, n740_adj_4990, n38278, n658, n39585, n585, 
        n39584, n950_adj_4991, n39355, n877_adj_4992, n39354, n314_adj_4993, 
        n39203, n512, n39583, n439, n39582, n804_adj_4994, n39353, 
        n241_adj_4995, n39202, n366, n39581, n293, n39580, n220, 
        n39579, n147_adj_4996, n39578, n5_adj_4997, n74, n38277;
    wire [20:0]n12088;
    
    wire n39577, n39576, n39575, n38276, n39574, n813_adj_4998, 
        n38275, n39573, n39572, n39571, n731_adj_4999, n39352, n168_adj_5000, 
        n39201, n886_adj_5001, n959_adj_5002, n1099, n39570, n1026, 
        n39569, n953, n39568, n658_adj_5003, n39351, n26_adj_5004, 
        n95_adj_5005, n880, n39567, n38274, n807, n39566, n734, 
        n39565, n661_adj_5006, n39564, n588_adj_5007, n39563, n585_adj_5008, 
        n39350, n630_adj_5009, n39200, n515_adj_5010, n39562, n512_adj_5011, 
        n39349, n557_adj_5012, n39199, n442_adj_5013, n39561, n369_adj_5014, 
        n39560, n38402, n38401, n296_adj_5017, n39559, n223_adj_5018, 
        n39558, n150_adj_5019, n39557, n8_adj_5020, n77_adj_5021;
    wire [19:0]n12969;
    
    wire n39556, n484_adj_5022, n39198, n39555, n39554, n39553, 
        n39552, n38400, n39551, n439_adj_5024, n39348, n411_adj_5025, 
        n39197, n38273, n366_adj_5026, n39347, n293_adj_5027, n39346, 
        n220_adj_5028, n39345, n38399, n338_adj_5030, n39196, n147_adj_5031, 
        n39344, n1102_adj_5032, n39550, n1029_adj_5033, n39549, n956_adj_5034, 
        n39548, n265_adj_5035, n39195, n883_adj_5036, n39547, n38272, 
        n810_adj_5037, n39546, n737_adj_5038, n39545, n664_adj_5039, 
        n39544, n591_adj_5040, n39543, n38398, n518_adj_5042, n39542, 
        n192_adj_5043, n39194, n38397, n5_adj_5045, n74_adj_5046, 
        n445_adj_5047, n39541, n50_adj_5048, n119_adj_5049, n39343, 
        n39342, n38271, n1120_adj_5050, n39193, n38396, n39341, 
        n1047_adj_5052, n39192, n38395, n38270, n39340, n372_adj_5054, 
        n39540, n974_adj_5055, n39191, n38394, n38393, n299_adj_5058, 
        n39539, n1032_adj_5059, n38392, n39339, n39338, n901_adj_5061, 
        n39190, n39337, n828_adj_5062, n39189, n1099_adj_5063, n39336, 
        n38391, n38390, n755_adj_5066, n39188, n38389, n38269, n682_adj_5068, 
        n39187, n38268, n1026_adj_5069, n39335, n609_adj_5070, n39186, 
        n38388, n226_adj_5072, n39538, n38267, n953_adj_5073, n39334, 
        n153_adj_5074, n39537, n536_adj_5075, n39185, n11_adj_5076, 
        n80_adj_5077;
    wire [18:0]n13768;
    
    wire n39536, n39535, n38266, n880_adj_5078, n39333, n39534, 
        n39533, n807_adj_5079, n39332, n734_adj_5080, n39331, n463_adj_5081, 
        n39184, n39532, n1105_adj_5083, n39531, n38387, n39530, 
        n39529, n39528, n39527, n39526, n39525, n38386, n39524, 
        n39330, n39523, n39522, n39329, n39183, n39521, n38385, 
        n39520, n39519, n39328, n38265, n39518;
    wire [17:0]n14489;
    
    wire n39517, n39516, n39515, n39514, n39513, n39512, n39511, 
        n39510, n39509, n39508, n39507, n39506, n39505, n39504, 
        n39503, n39502, n39501, n39500, n39499, n39327, n38384, 
        n39498, n39497, n39496, n39495, n39494, n39493, n39492, 
        n39182, n39491, n39490, n39489, n39488, n39487, n39486, 
        n39485, n39484, n39483, n39482, n39481, n39480, n39479, 
        n39326, n38383, n38382, n38264, n38381, n39478, n38263, 
        n38380, n38262, n39325, n39181, n38261, n38260, n38379, 
        n38378, n39477, n38377, n39324, n39180, n38376, n38375, 
        n39179, n38374, n39476, n39178, n39323, n38373, n39475, 
        n39474, n39473, n39472, n39471, n38259, n38372, n4_adj_5084, 
        n38050, n41_adj_5085, n39_adj_5086, n45_adj_5087, n37_adj_5088, 
        n29_adj_5089, n31_adj_5090, n43_adj_5091, n35_adj_5092, n23_adj_5093, 
        n25_adj_5094, n33_adj_5095, n11_adj_5096, n13_adj_5097, n15_adj_5098, 
        n27_adj_5099, n9_adj_5100, n17_adj_5101, n19_adj_5102, n21_adj_5103, 
        n37968, n47394, n47387, n12_adj_5104, n10_adj_5105, n30_adj_5106, 
        n47650, n47644, n47971, n47813, n48011, n16_adj_5107, n47827, 
        n47828, n8_adj_5108, n24_adj_5109, n47312, n47809, n47625, 
        n4_adj_5110, n47823, n47824, n47349, n48029, n47627, n48067, 
        n48068, n48058, n47315, n47965, n40, n47967, n39_adj_5111, 
        n41_adj_5112, n45_adj_5113, n37_adj_5114, n43_adj_5115, n23_adj_5116, 
        n25_adj_5117, n29_adj_5118, n31_adj_5119, n35_adj_5120, n11_adj_5121, 
        n13_adj_5122, n27_adj_5123, n15_adj_5124, n33_adj_5125, n9_adj_5126, 
        n17_adj_5127, n19_adj_5128, n21_adj_5129, n47430, n47424, 
        n12_adj_5130, n10_adj_5131, n30_adj_5132, n47689, n47685, 
        n47981, n47837, n48019, n16_adj_5133, n47911, n47912, n8_adj_5134, 
        n24_adj_5135, n47410, n47807, n47615, n4_adj_5136, n47909, 
        n47910, n47420, n47973, n47617, n48055, n48056, n48036, 
        n47412, n47961, n47623, n48017, n17_adj_5137, n9_adj_5138, 
        n11_adj_5139, n47513, n47511, n49340, n47875, n47749, n49322, 
        n47747, n47745, n49316, n16_adj_5140, n47478, n47721, n47717, 
        n47991, n47853, n47751, n49309, n12_adj_5141, n47939, n47499, 
        n49307, n47869, n49333, n47995, n49298, n16_adj_5142, n47480, 
        n24_adj_5143, n6_adj_5144, n47927, n47928, n4_adj_5145, n47917;
    
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [22]), .O(n13_adj_4726));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_5267_3 (.CI(n39161), .I0(n18513[0]), .I1(n195), .CO(n39162));
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32377_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n47462), 
            .O(n47458));
    defparam i32377_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32924_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n47454), 
            .O(n48005));   // verilog/motorControl.v(31[38:63])
    defparam i32924_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4726), .I1(n18), .I2(n38034), .I3(n4), 
            .O(n44653));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5267_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n18416[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32526_3_lut (.I0(n47918), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n47607));   // verilog/motorControl.v(31[38:63])
    defparam i32526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32972_4_lut (.I0(n47607), .I1(n48005), .I2(n35), .I3(n47458), 
            .O(n48053));   // verilog/motorControl.v(31[38:63])
    defparam i32972_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32973_3_lut (.I0(n48053), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n48054));   // verilog/motorControl.v(31[38:63])
    defparam i32973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32959_3_lut (.I0(n48054), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n48040));   // verilog/motorControl.v(31[38:63])
    defparam i32959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7), .I3(GND_net), 
            .O(n6));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32838_3_lut (.I0(n6), .I1(\PID_CONTROLLER.integral [10]), .I2(n21), 
            .I3(GND_net), .O(n47919));   // verilog/motorControl.v(31[38:63])
    defparam i32838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32839_3_lut (.I0(n47919), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23), .I3(GND_net), .O(n47920));   // verilog/motorControl.v(31[38:63])
    defparam i32839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32364_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n47468), 
            .O(n47445));
    defparam i32364_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5267_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n39161));
    SB_LUT4 add_5140_14_lut (.I0(GND_net), .I1(n17233[11]), .I2(n980), 
            .I3(n39160), .O(n16869[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32724_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n47442), 
            .O(n47805));   // verilog/motorControl.v(31[38:63])
    defparam i32724_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32524_3_lut (.I0(n47920), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25), .I3(GND_net), .O(n47605));   // verilog/motorControl.v(31[38:63])
    defparam i32524_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n38370), .I0(GND_net), .I1(n1_adj_5146[14]), 
            .CO(n38371));
    SB_LUT4 i32367_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n48023), 
            .O(n47448));
    defparam i32367_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5140_13_lut (.I0(GND_net), .I1(n17233[10]), .I2(n907), 
            .I3(n39159), .O(n16869[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32878_4_lut (.I0(n47605), .I1(n47805), .I2(n45), .I3(n47445), 
            .O(n47959));   // verilog/motorControl.v(31[38:63])
    defparam i32878_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_5146[13]), .I3(n38369), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32532_3_lut (.I0(n48040), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n47613));   // verilog/motorControl.v(31[38:63])
    defparam i32532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n38369), .I0(GND_net), .I1(n1_adj_5146[13]), 
            .CO(n38370));
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5140_13 (.CI(n39159), .I0(n17233[10]), .I1(n907), .CO(n39160));
    SB_LUT4 i32934_4_lut (.I0(n47613), .I1(n47959), .I2(n45), .I3(n47448), 
            .O(n48015));   // verilog/motorControl.v(31[38:63])
    defparam i32934_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4729));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n38257), .O(duty_23__N_3772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n38257), .I0(n106[16]), .I1(n155[16]), .CO(n38258));
    SB_LUT4 add_5140_12_lut (.I0(GND_net), .I1(n17233[9]), .I2(n834), 
            .I3(n39158), .O(n16869[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_12 (.CI(n39158), .I0(n17233[9]), .I1(n834), .CO(n39159));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_5146[12]), .I3(n38368), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5140_11_lut (.I0(GND_net), .I1(n17233[8]), .I2(n761), 
            .I3(n39157), .O(n16869[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32844_3_lut (.I0(n4_adj_4729), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n47925));   // verilog/motorControl.v(31[10:34])
    defparam i32844_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5140_11 (.CI(n39157), .I0(n17233[8]), .I1(n761), .CO(n39158));
    SB_LUT4 add_5140_10_lut (.I0(GND_net), .I1(n17233[7]), .I2(n688), 
            .I3(n39156), .O(n16869[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32845_3_lut (.I0(n47925), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n47926));   // verilog/motorControl.v(31[10:34])
    defparam i32845_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32412_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n49304), 
            .I2(IntegralLimit[16]), .I3(n47739), .O(n47493));
    defparam i32412_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_364_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n49328));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_364_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5037_13_lut (.I0(GND_net), .I1(n15713[10]), .I2(n895), 
            .I3(n39469), .O(n15136[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32922_4_lut (.I0(n30_adj_4732), .I1(n10_adj_4733), .I2(n49328), 
            .I3(n47491), .O(n48003));   // verilog/motorControl.v(31[10:34])
    defparam i32922_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5140_10 (.CI(n39156), .I0(n17233[7]), .I1(n688), .CO(n39157));
    SB_LUT4 i32516_3_lut (.I0(n47926), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n47597));   // verilog/motorControl.v(31[10:34])
    defparam i32516_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32970_4_lut (.I0(n47597), .I1(n48003), .I2(n49328), .I3(n47493), 
            .O(n48051));   // verilog/motorControl.v(31[10:34])
    defparam i32970_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32971_3_lut (.I0(n48051), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n48052));   // verilog/motorControl.v(31[10:34])
    defparam i32971_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32961_3_lut (.I0(n48052), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n48042));   // verilog/motorControl.v(31[10:34])
    defparam i32961_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32403_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n49295), 
            .I2(IntegralLimit[21]), .I3(n48047), .O(n47484));
    defparam i32403_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i32876_4_lut (.I0(n47595), .I1(n47803), .I2(n49291), .I3(n47482), 
            .O(n47957));   // verilog/motorControl.v(31[10:34])
    defparam i32876_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32522_3_lut (.I0(n48042), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n47603));   // verilog/motorControl.v(31[10:34])
    defparam i32522_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32935_3_lut (.I0(n48015), .I1(\PID_CONTROLLER.integral_23__N_3723 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3722 ));   // verilog/motorControl.v(31[38:63])
    defparam i32935_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32932_4_lut (.I0(n47603), .I1(n47957), .I2(n49291), .I3(n47484), 
            .O(n48013));   // verilog/motorControl.v(31[10:34])
    defparam i32932_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_850_4_lut  (.I0(n48013), .I1(\PID_CONTROLLER.integral_23__N_3722 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3720 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_850_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5140_9_lut (.I0(GND_net), .I1(n17233[6]), .I2(n615), .I3(n39155), 
            .O(n16869[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_9 (.CI(n39155), .I0(n17233[6]), .I1(n615), .CO(n39156));
    SB_CARRY add_4868_21 (.CI(n39321), .I0(n12529[18]), .I1(GND_net), 
            .CO(n39322));
    SB_LUT4 add_4868_20_lut (.I0(GND_net), .I1(n12529[17]), .I2(GND_net), 
            .I3(n39320), .O(n11605[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_8_lut (.I0(GND_net), .I1(n17233[5]), .I2(n542), .I3(n39154), 
            .O(n16869[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_8 (.CI(n39154), .I0(n17233[5]), .I1(n542), .CO(n39155));
    SB_CARRY add_5113_12 (.CI(n39176), .I0(n16869[9]), .I1(n831), .CO(n39177));
    SB_CARRY add_5037_13 (.CI(n39469), .I0(n15713[10]), .I1(n895), .CO(n39470));
    SB_LUT4 add_5140_7_lut (.I0(GND_net), .I1(n17233[4]), .I2(n469), .I3(n39153), 
            .O(n16869[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_7 (.CI(n39153), .I0(n17233[4]), .I1(n469), .CO(n39154));
    SB_LUT4 add_5140_6_lut (.I0(GND_net), .I1(n17233[3]), .I2(n396), .I3(n39152), 
            .O(n16869[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_6 (.CI(n39152), .I0(n17233[3]), .I1(n396), .CO(n39153));
    SB_LUT4 add_5037_12_lut (.I0(GND_net), .I1(n15713[9]), .I2(n822), 
            .I3(n39468), .O(n15136[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n38368), .I0(GND_net), .I1(n1_adj_5146[12]), 
            .CO(n38369));
    SB_LUT4 add_5113_11_lut (.I0(GND_net), .I1(n16869[8]), .I2(n758), 
            .I3(n39175), .O(n16449[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_12 (.CI(n39468), .I0(n15713[9]), .I1(n822), .CO(n39469));
    SB_LUT4 add_5037_11_lut (.I0(GND_net), .I1(n15713[8]), .I2(n749), 
            .I3(n39467), .O(n15136[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_11 (.CI(n39467), .I0(n15713[8]), .I1(n749), .CO(n39468));
    SB_LUT4 add_5037_10_lut (.I0(GND_net), .I1(n15713[7]), .I2(n676), 
            .I3(n39466), .O(n15136[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_10 (.CI(n39466), .I0(n15713[7]), .I1(n676), .CO(n39467));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_5146[11]), .I3(n38367), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5113_11 (.CI(n39175), .I0(n16869[8]), .I1(n758), .CO(n39176));
    SB_LUT4 add_5037_9_lut (.I0(GND_net), .I1(n15713[6]), .I2(n603), .I3(n39465), 
            .O(n15136[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5140_5_lut (.I0(GND_net), .I1(n17233[2]), .I2(n323), .I3(n39151), 
            .O(n16869[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_9 (.CI(n39465), .I0(n15713[6]), .I1(n603), .CO(n39466));
    SB_LUT4 add_5037_8_lut (.I0(GND_net), .I1(n15713[5]), .I2(n530), .I3(n39464), 
            .O(n15136[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_8 (.CI(n39464), .I0(n15713[5]), .I1(n530), .CO(n39465));
    SB_LUT4 add_5113_10_lut (.I0(GND_net), .I1(n16869[7]), .I2(n685), 
            .I3(n39174), .O(n16449[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_20 (.CI(n39320), .I0(n12529[17]), .I1(GND_net), 
            .CO(n39321));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n38367), .I0(GND_net), .I1(n1_adj_5146[11]), 
            .CO(n38368));
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5140_5 (.CI(n39151), .I0(n17233[2]), .I1(n323), .CO(n39152));
    SB_LUT4 add_5140_4_lut (.I0(GND_net), .I1(n17233[1]), .I2(n250), .I3(n39150), 
            .O(n16869[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_4 (.CI(n39150), .I0(n17233[1]), .I1(n250), .CO(n39151));
    SB_LUT4 add_5140_3_lut (.I0(GND_net), .I1(n17233[0]), .I2(n177), .I3(n39149), 
            .O(n16869[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_3 (.CI(n39149), .I0(n17233[0]), .I1(n177), .CO(n39150));
    SB_LUT4 add_5140_2_lut (.I0(GND_net), .I1(n35_adj_4736), .I2(n104), 
            .I3(GND_net), .O(n16869[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5140_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5140_2 (.CI(GND_net), .I0(n35_adj_4736), .I1(n104), .CO(n39149));
    SB_LUT4 add_5165_13_lut (.I0(GND_net), .I1(n17545[10]), .I2(n910), 
            .I3(n39148), .O(n17233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_5146[10]), .I3(n38366), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5165_12_lut (.I0(GND_net), .I1(n17545[9]), .I2(n837), 
            .I3(n39147), .O(n17233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_12 (.CI(n39147), .I0(n17545[9]), .I1(n837), .CO(n39148));
    SB_LUT4 add_5165_11_lut (.I0(GND_net), .I1(n17545[8]), .I2(n764), 
            .I3(n39146), .O(n17233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_11 (.CI(n39146), .I0(n17545[8]), .I1(n764), .CO(n39147));
    SB_LUT4 add_5165_10_lut (.I0(GND_net), .I1(n17545[7]), .I2(n691), 
            .I3(n39145), .O(n17233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_10 (.CI(n39145), .I0(n17545[7]), .I1(n691), .CO(n39146));
    SB_LUT4 add_5165_9_lut (.I0(GND_net), .I1(n17545[6]), .I2(n618), .I3(n39144), 
            .O(n17233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_9 (.CI(n39144), .I0(n17545[6]), .I1(n618), .CO(n39145));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n38366), .I0(GND_net), .I1(n1_adj_5146[10]), 
            .CO(n38367));
    SB_LUT4 add_5165_8_lut (.I0(GND_net), .I1(n17545[5]), .I2(n545), .I3(n39143), 
            .O(n17233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4868_19_lut (.I0(GND_net), .I1(n12529[16]), .I2(GND_net), 
            .I3(n39319), .O(n11605[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_7_lut (.I0(GND_net), .I1(n15713[4]), .I2(n457), .I3(n39463), 
            .O(n15136[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_7 (.CI(n39463), .I0(n15713[4]), .I1(n457), .CO(n39464));
    SB_LUT4 add_5037_6_lut (.I0(GND_net), .I1(n15713[3]), .I2(n384), .I3(n39462), 
            .O(n15136[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_19 (.CI(n39319), .I0(n12529[16]), .I1(GND_net), 
            .CO(n39320));
    SB_CARRY add_5037_6 (.CI(n39462), .I0(n15713[3]), .I1(n384), .CO(n39463));
    SB_LUT4 add_5037_5_lut (.I0(GND_net), .I1(n15713[2]), .I2(n311), .I3(n39461), 
            .O(n15136[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5037_5 (.CI(n39461), .I0(n15713[2]), .I1(n311), .CO(n39462));
    SB_LUT4 add_5037_4_lut (.I0(GND_net), .I1(n15713[1]), .I2(n238), .I3(n39460), 
            .O(n15136[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_4 (.CI(n39460), .I0(n15713[1]), .I1(n238), .CO(n39461));
    SB_LUT4 add_5037_3_lut (.I0(GND_net), .I1(n15713[0]), .I2(n165), .I3(n39459), 
            .O(n15136[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_3 (.CI(n39459), .I0(n15713[0]), .I1(n165), .CO(n39460));
    SB_CARRY add_5113_10 (.CI(n39174), .I0(n16869[7]), .I1(n685), .CO(n39175));
    SB_LUT4 add_5037_2_lut (.I0(GND_net), .I1(n23_adj_4738), .I2(n92), 
            .I3(GND_net), .O(n15136[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5037_2 (.CI(GND_net), .I0(n23_adj_4738), .I1(n92), .CO(n39459));
    SB_LUT4 add_4868_18_lut (.I0(GND_net), .I1(n12529[15]), .I2(GND_net), 
            .I3(n39318), .O(n11605[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_9_lut (.I0(GND_net), .I1(n18353[6]), .I2(n630), .I3(n39458), 
            .O(n18209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_18 (.CI(n39318), .I0(n12529[15]), .I1(GND_net), 
            .CO(n39319));
    SB_LUT4 add_4868_17_lut (.I0(GND_net), .I1(n12529[14]), .I2(GND_net), 
            .I3(n39317), .O(n11605[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4741));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4744));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20568_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20568_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4745));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4747));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4749), .I1(\Kp[4] ), .I2(n18633[2]), 
            .I3(n1[18]), .O(n18584[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4750));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5165_8 (.CI(n39143), .I0(n17545[5]), .I1(n545), .CO(n39144));
    SB_LUT4 add_5165_7_lut (.I0(GND_net), .I1(n17545[4]), .I2(n472), .I3(n39142), 
            .O(n17233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5245_8_lut (.I0(GND_net), .I1(n18353[5]), .I2(n557), .I3(n39457), 
            .O(n18209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_7 (.CI(n39142), .I0(n17545[4]), .I1(n472), .CO(n39143));
    SB_LUT4 add_5165_6_lut (.I0(GND_net), .I1(n17545[3]), .I2(n399), .I3(n39141), 
            .O(n17233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_6 (.CI(n39141), .I0(n17545[3]), .I1(n399), .CO(n39142));
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5245_8 (.CI(n39457), .I0(n18353[5]), .I1(n557), .CO(n39458));
    SB_LUT4 i24374_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n18681[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24374_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4754));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4756));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5165_5_lut (.I0(GND_net), .I1(n17545[2]), .I2(n326), .I3(n39140), 
            .O(n17233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_5 (.CI(n39140), .I0(n17545[2]), .I1(n326), .CO(n39141));
    SB_CARRY add_4868_17 (.CI(n39317), .I0(n12529[14]), .I1(GND_net), 
            .CO(n39318));
    SB_LUT4 add_4868_16_lut (.I0(GND_net), .I1(n12529[13]), .I2(n1102), 
            .I3(n39316), .O(n11605[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_7_lut (.I0(GND_net), .I1(n18353[4]), .I2(n484), .I3(n39456), 
            .O(n18209[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4868_16 (.CI(n39316), .I0(n12529[13]), .I1(n1102), .CO(n39317));
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(n1[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4757));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4760));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4762));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4763));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5165_4_lut (.I0(GND_net), .I1(n17545[1]), .I2(n253), .I3(n39139), 
            .O(n17233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1549 (.I0(n4_adj_4764), .I1(\Kp[3] ), .I2(n18664[1]), 
            .I3(n1[19]), .O(n18633[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1549.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1550 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4765));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1550.LUT_INIT = 16'h9c50;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4766));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24578_4_lut (.I0(n18633[2]), .I1(\Kp[4] ), .I2(n6_adj_4749), 
            .I3(n1[18]), .O(n8_adj_4767));   // verilog/motorControl.v(34[16:22])
    defparam i24578_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), .I3(n1[21]), 
            .O(n11_adj_4768));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i24524_4_lut (.I0(n18664[1]), .I1(\Kp[3] ), .I2(n4_adj_4764), 
            .I3(n1[19]), .O(n6_adj_4769));   // verilog/motorControl.v(34[16:22])
    defparam i24524_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i24376_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n37861));   // verilog/motorControl.v(34[16:22])
    defparam i24376_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4769), .I1(n11_adj_4768), .I2(n8_adj_4767), 
            .I3(n12_adj_4765), .O(n18_adj_4770));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1551 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), 
            .I3(n1[22]), .O(n13_adj_4771));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1551.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1552 (.I0(n13_adj_4771), .I1(n18_adj_4770), .I2(n37861), 
            .I3(n4_adj_4772), .O(n44771));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1552.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4773));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4774));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4775));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5165_4 (.CI(n39139), .I0(n17545[1]), .I1(n253), .CO(n39140));
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5165_3_lut (.I0(GND_net), .I1(n17545[0]), .I2(n180), .I3(n39138), 
            .O(n17233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_3 (.CI(n39138), .I0(n17545[0]), .I1(n180), .CO(n39139));
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5165_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n17233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_5146[9]), .I3(n38365), .O(n19_adj_4777)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5165_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n39138));
    SB_LUT4 add_5279_7_lut (.I0(GND_net), .I1(n44771), .I2(n490), .I3(n39137), 
            .O(n18513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5279_6_lut (.I0(GND_net), .I1(n18584[3]), .I2(n417), .I3(n39136), 
            .O(n18513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_7 (.CI(n39456), .I0(n18353[4]), .I1(n484), .CO(n39457));
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4778));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n38256), .O(duty_23__N_3772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4868_15_lut (.I0(GND_net), .I1(n12529[12]), .I2(n1029), 
            .I3(n39315), .O(n11605[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5113_9_lut (.I0(GND_net), .I1(n16869[6]), .I2(n612), .I3(n39173), 
            .O(n16449[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4780));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5279_6 (.CI(n39136), .I0(n18584[3]), .I1(n417), .CO(n39137));
    SB_LUT4 add_5279_5_lut (.I0(GND_net), .I1(n18584[2]), .I2(n344), .I3(n39135), 
            .O(n18513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5279_5 (.CI(n39135), .I0(n18584[2]), .I1(n344), .CO(n39136));
    SB_LUT4 add_5279_4_lut (.I0(GND_net), .I1(n18584[1]), .I2(n271), .I3(n39134), 
            .O(n18513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5279_4 (.CI(n39134), .I0(n18584[1]), .I1(n271), .CO(n39135));
    SB_LUT4 add_5245_6_lut (.I0(GND_net), .I1(n18353[3]), .I2(n411), .I3(n39455), 
            .O(n18209[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_15 (.CI(n39315), .I0(n12529[12]), .I1(n1029), .CO(n39316));
    SB_LUT4 add_4868_14_lut (.I0(GND_net), .I1(n12529[11]), .I2(n956), 
            .I3(n39314), .O(n11605[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5279_3_lut (.I0(GND_net), .I1(n18584[0]), .I2(n198), .I3(n39133), 
            .O(n18513[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n38365), .I0(GND_net), .I1(n1_adj_5146[9]), 
            .CO(n38366));
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5245_6 (.CI(n39455), .I0(n18353[3]), .I1(n411), .CO(n39456));
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5279_3 (.CI(n39133), .I0(n18584[0]), .I1(n198), .CO(n39134));
    SB_LUT4 add_5279_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n18513[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5279_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4868_14 (.CI(n39314), .I0(n12529[11]), .I1(n956), .CO(n39315));
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5113_9 (.CI(n39173), .I0(n16869[6]), .I1(n612), .CO(n39174));
    SB_CARRY add_5279_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n39133));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_5146[8]), .I3(n38364), .O(n17_adj_4781)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5245_5_lut (.I0(GND_net), .I1(n18353[2]), .I2(n338), .I3(n39454), 
            .O(n18209[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_5 (.CI(n39454), .I0(n18353[2]), .I1(n338), .CO(n39455));
    SB_LUT4 add_5113_8_lut (.I0(GND_net), .I1(n16869[5]), .I2(n539), .I3(n39172), 
            .O(n16449[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4782));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4868_13_lut (.I0(GND_net), .I1(n12529[10]), .I2(n883), 
            .I3(n39313), .O(n11605[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_4_lut (.I0(GND_net), .I1(n18353[1]), .I2(n265), .I3(n39453), 
            .O(n18209[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_4 (.CI(n39453), .I0(n18353[1]), .I1(n265), .CO(n39454));
    SB_CARRY add_5113_8 (.CI(n39172), .I0(n16869[5]), .I1(n539), .CO(n39173));
    SB_LUT4 add_5113_7_lut (.I0(GND_net), .I1(n16869[4]), .I2(n466), .I3(n39171), 
            .O(n16449[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5245_3_lut (.I0(GND_net), .I1(n18353[0]), .I2(n192), .I3(n39452), 
            .O(n18209[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_3 (.CI(n39452), .I0(n18353[0]), .I1(n192), .CO(n39453));
    SB_LUT4 add_5245_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n18209[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5245_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_13 (.CI(n39313), .I0(n12529[10]), .I1(n883), .CO(n39314));
    SB_LUT4 add_4868_12_lut (.I0(GND_net), .I1(n12529[9]), .I2(n810), 
            .I3(n39312), .O(n11605[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_12 (.CI(n39312), .I0(n12529[9]), .I1(n810), .CO(n39313));
    SB_CARRY add_5113_7 (.CI(n39171), .I0(n16869[4]), .I1(n466), .CO(n39172));
    SB_LUT4 add_4868_11_lut (.I0(GND_net), .I1(n12529[8]), .I2(n737), 
            .I3(n39311), .O(n11605[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5113_6_lut (.I0(GND_net), .I1(n16869[3]), .I2(n393), .I3(n39170), 
            .O(n16449[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5113_6 (.CI(n39170), .I0(n16869[3]), .I1(n393), .CO(n39171));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n38364), .I0(GND_net), .I1(n1_adj_5146[8]), 
            .CO(n38365));
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4783));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_5146[7]), .I3(n38363), .O(n15_adj_4784)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5113_5_lut (.I0(GND_net), .I1(n16869[2]), .I2(n320), .I3(n39169), 
            .O(n16449[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5245_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n39452));
    SB_CARRY add_4868_11 (.CI(n39311), .I0(n12529[8]), .I1(n737), .CO(n39312));
    SB_LUT4 add_4868_10_lut (.I0(GND_net), .I1(n12529[7]), .I2(n664), 
            .I3(n39310), .O(n11605[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_17_lut (.I0(GND_net), .I1(n16224[14]), .I2(GND_net), 
            .I3(n39451), .O(n15713[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_16_lut (.I0(GND_net), .I1(n16224[13]), .I2(n1117), 
            .I3(n39450), .O(n15713[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_16 (.CI(n39450), .I0(n16224[13]), .I1(n1117), .CO(n39451));
    SB_LUT4 add_5069_15_lut (.I0(GND_net), .I1(n16224[12]), .I2(n1044), 
            .I3(n39449), .O(n15713[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4868_10 (.CI(n39310), .I0(n12529[7]), .I1(n664), .CO(n39311));
    SB_LUT4 add_4868_9_lut (.I0(GND_net), .I1(n12529[6]), .I2(n591), .I3(n39309), 
            .O(n11605[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_9 (.CI(n39309), .I0(n12529[6]), .I1(n591), .CO(n39310));
    SB_LUT4 add_4868_8_lut (.I0(GND_net), .I1(n12529[5]), .I2(n518), .I3(n39308), 
            .O(n11605[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_8 (.CI(n39308), .I0(n12529[5]), .I1(n518), .CO(n39309));
    SB_LUT4 add_4868_7_lut (.I0(GND_net), .I1(n12529[4]), .I2(n445), .I3(n39307), 
            .O(n11605[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_7 (.CI(n39307), .I0(n12529[4]), .I1(n445), .CO(n39308));
    SB_CARRY add_5069_15 (.CI(n39449), .I0(n16224[12]), .I1(n1044), .CO(n39450));
    SB_LUT4 add_4868_6_lut (.I0(GND_net), .I1(n12529[3]), .I2(n372), .I3(n39306), 
            .O(n11605[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_6 (.CI(n39306), .I0(n12529[3]), .I1(n372), .CO(n39307));
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4868_5_lut (.I0(GND_net), .I1(n12529[2]), .I2(n299), .I3(n39305), 
            .O(n11605[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4785));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4786));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4787));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4788));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5069_14_lut (.I0(GND_net), .I1(n16224[11]), .I2(n971), 
            .I3(n39448), .O(n15713[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4789));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_17 (.CI(n38256), .I0(n106[15]), .I1(n155[15]), .CO(n38257));
    SB_CARRY add_5113_5 (.CI(n39169), .I0(n16869[2]), .I1(n320), .CO(n39170));
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4790));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4791));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4792));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4793));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4868_5 (.CI(n39305), .I0(n12529[2]), .I1(n299), .CO(n39306));
    SB_LUT4 add_5113_4_lut (.I0(GND_net), .I1(n16869[1]), .I2(n247_adj_4794), 
            .I3(n39168), .O(n16449[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_14 (.CI(n39448), .I0(n16224[11]), .I1(n971), .CO(n39449));
    SB_LUT4 add_4868_4_lut (.I0(GND_net), .I1(n12529[1]), .I2(n226), .I3(n39304), 
            .O(n11605[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5113_4 (.CI(n39168), .I0(n16869[1]), .I1(n247_adj_4794), 
            .CO(n39169));
    SB_LUT4 add_5113_3_lut (.I0(GND_net), .I1(n16869[0]), .I2(n174_adj_4795), 
            .I3(n39167), .O(n16449[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5113_3 (.CI(n39167), .I0(n16869[0]), .I1(n174_adj_4795), 
            .CO(n39168));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n38363), .I0(GND_net), .I1(n1_adj_5146[7]), 
            .CO(n38364));
    SB_LUT4 add_5069_13_lut (.I0(GND_net), .I1(n16224[10]), .I2(n898), 
            .I3(n39447), .O(n15713[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4796));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4797));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4798));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4799));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_5146[6]), .I3(n38362), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n38255), .O(duty_23__N_3772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_13 (.CI(n39447), .I0(n16224[10]), .I1(n898), .CO(n39448));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3648[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5069_12_lut (.I0(GND_net), .I1(n16224[9]), .I2(n825), 
            .I3(n39446), .O(n15713[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_4868_4 (.CI(n39304), .I0(n12529[1]), .I1(n226), .CO(n39305));
    SB_CARRY add_5069_12 (.CI(n39446), .I0(n16224[9]), .I1(n825), .CO(n39447));
    SB_LUT4 add_4868_3_lut (.I0(GND_net), .I1(n12529[0]), .I2(n153), .I3(n39303), 
            .O(n11605[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4868_3 (.CI(n39303), .I0(n12529[0]), .I1(n153), .CO(n39304));
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4801));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5113_2_lut (.I0(GND_net), .I1(n32_adj_4802), .I2(n101_adj_4803), 
            .I3(GND_net), .O(n16449[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4868_2_lut (.I0(GND_net), .I1(n11_adj_4804), .I2(n80), 
            .I3(GND_net), .O(n11605[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n38362), .I0(GND_net), .I1(n1_adj_5146[6]), 
            .CO(n38363));
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5113_2 (.CI(GND_net), .I0(n32_adj_4802), .I1(n101_adj_4803), 
            .CO(n39167));
    SB_CARRY add_12_16 (.CI(n38255), .I0(n106[14]), .I1(n155[14]), .CO(n38256));
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n38254), .O(duty_23__N_3772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_8_lut (.I0(GND_net), .I1(n18513[5]), .I2(n560_adj_4805), 
            .I3(n39166), .O(n18416[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_7_lut (.I0(GND_net), .I1(n18513[4]), .I2(n487_adj_4806), 
            .I3(n39165), .O(n18416[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5069_11_lut (.I0(GND_net), .I1(n16224[8]), .I2(n752), 
            .I3(n39445), .O(n15713[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4808));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_15 (.CI(n38254), .I0(n106[13]), .I1(n155[13]), .CO(n38255));
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4809));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_5146[5]), .I3(n38361), .O(n11_adj_4811)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5069_11 (.CI(n39445), .I0(n16224[8]), .I1(n752), .CO(n39446));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n38361), .I0(GND_net), .I1(n1_adj_5146[5]), 
            .CO(n38362));
    SB_CARRY add_4868_2 (.CI(GND_net), .I0(n11_adj_4804), .I1(n80), .CO(n39303));
    SB_CARRY add_5267_7 (.CI(n39165), .I0(n18513[4]), .I1(n487_adj_4806), 
            .CO(n39166));
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4812));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_5146[4]), .I3(n38360), .O(n9_adj_4813)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5069_10_lut (.I0(GND_net), .I1(n16224[7]), .I2(n679), 
            .I3(n39444), .O(n15713[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5069_10 (.CI(n39444), .I0(n16224[7]), .I1(n679), .CO(n39445));
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_21_lut (.I0(GND_net), .I1(n13369[18]), .I2(GND_net), 
            .I3(n39302), .O(n12529[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4817));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5069_9_lut (.I0(GND_net), .I1(n16224[6]), .I2(n606), .I3(n39443), 
            .O(n15713[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5188_12_lut (.I0(GND_net), .I1(n17809[9]), .I2(n840), 
            .I3(n39101), .O(n17545[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5188_11_lut (.I0(GND_net), .I1(n17809[8]), .I2(n767_adj_4818), 
            .I3(n39100), .O(n17545[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_9 (.CI(n39443), .I0(n16224[6]), .I1(n606), .CO(n39444));
    SB_LUT4 add_4909_20_lut (.I0(GND_net), .I1(n13369[17]), .I2(GND_net), 
            .I3(n39301), .O(n12529[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_6_lut (.I0(GND_net), .I1(n18513[3]), .I2(n414_adj_4819), 
            .I3(n39164), .O(n18416[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4820));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4909_20 (.CI(n39301), .I0(n13369[17]), .I1(GND_net), 
            .CO(n39302));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n38360), .I0(GND_net), .I1(n1_adj_5146[4]), 
            .CO(n38361));
    SB_LUT4 add_5069_8_lut (.I0(GND_net), .I1(n16224[5]), .I2(n533), .I3(n39442), 
            .O(n15713[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4821));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5188_11 (.CI(n39100), .I0(n17809[8]), .I1(n767_adj_4818), 
            .CO(n39101));
    SB_LUT4 add_4909_19_lut (.I0(GND_net), .I1(n13369[16]), .I2(GND_net), 
            .I3(n39300), .O(n12529[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_19 (.CI(n39300), .I0(n13369[16]), .I1(GND_net), 
            .CO(n39301));
    SB_LUT4 add_4909_18_lut (.I0(GND_net), .I1(n13369[15]), .I2(GND_net), 
            .I3(n39299), .O(n12529[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_5146[3]), .I3(n38359), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5188_10_lut (.I0(GND_net), .I1(n17809[7]), .I2(n694_adj_4822), 
            .I3(n39099), .O(n17545[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_8 (.CI(n39442), .I0(n16224[5]), .I1(n533), .CO(n39443));
    SB_LUT4 add_5069_7_lut (.I0(GND_net), .I1(n16224[4]), .I2(n460), .I3(n39441), 
            .O(n15713[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n38253), .O(duty_23__N_3772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_7 (.CI(n39441), .I0(n16224[4]), .I1(n460), .CO(n39442));
    SB_CARRY add_5267_6 (.CI(n39164), .I0(n18513[3]), .I1(n414_adj_4819), 
            .CO(n39165));
    SB_LUT4 add_5267_3_lut (.I0(GND_net), .I1(n18513[0]), .I2(n195), .I3(n39161), 
            .O(n18416[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_10 (.CI(n39099), .I0(n17809[7]), .I1(n694_adj_4822), 
            .CO(n39100));
    SB_LUT4 add_5188_9_lut (.I0(GND_net), .I1(n17809[6]), .I2(n621_adj_4823), 
            .I3(n39098), .O(n17545[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_9 (.CI(n39098), .I0(n17809[6]), .I1(n621_adj_4823), 
            .CO(n39099));
    SB_LUT4 add_5069_6_lut (.I0(GND_net), .I1(n16224[3]), .I2(n387), .I3(n39440), 
            .O(n15713[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5188_8_lut (.I0(GND_net), .I1(n17809[5]), .I2(n548_adj_4824), 
            .I3(n39097), .O(n17545[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_8 (.CI(n39097), .I0(n17809[5]), .I1(n548_adj_4824), 
            .CO(n39098));
    SB_LUT4 add_5188_7_lut (.I0(GND_net), .I1(n17809[4]), .I2(n475_adj_4825), 
            .I3(n39096), .O(n17545[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_7 (.CI(n39096), .I0(n17809[4]), .I1(n475_adj_4825), 
            .CO(n39097));
    SB_LUT4 add_5188_6_lut (.I0(GND_net), .I1(n17809[3]), .I2(n402_adj_4826), 
            .I3(n39095), .O(n17545[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_6 (.CI(n39095), .I0(n17809[3]), .I1(n402_adj_4826), 
            .CO(n39096));
    SB_LUT4 add_5188_5_lut (.I0(GND_net), .I1(n17809[2]), .I2(n329_adj_4827), 
            .I3(n39094), .O(n17545[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_5 (.CI(n39094), .I0(n17809[2]), .I1(n329_adj_4827), 
            .CO(n39095));
    SB_LUT4 add_5188_4_lut (.I0(GND_net), .I1(n17809[1]), .I2(n256_adj_4828), 
            .I3(n39093), .O(n17545[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4829));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4909_18 (.CI(n39299), .I0(n13369[15]), .I1(GND_net), 
            .CO(n39300));
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4830));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5188_4 (.CI(n39093), .I0(n17809[1]), .I1(n256_adj_4828), 
            .CO(n39094));
    SB_CARRY add_5069_6 (.CI(n39440), .I0(n16224[3]), .I1(n387), .CO(n39441));
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5188_3_lut (.I0(GND_net), .I1(n17809[0]), .I2(n183_adj_4832), 
            .I3(n39092), .O(n17545[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4833));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4835));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5188_3 (.CI(n39092), .I0(n17809[0]), .I1(n183_adj_4832), 
            .CO(n39093));
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4836));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n38359), .I0(GND_net), .I1(n1_adj_5146[3]), 
            .CO(n38360));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_5146[2]), .I3(n38358), .O(n5_adj_4838)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n38358), .I0(GND_net), .I1(n1_adj_5146[2]), 
            .CO(n38359));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_5146[1]), .I3(n38357), .O(n3_adj_4840)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5188_2_lut (.I0(GND_net), .I1(n41_adj_4842), .I2(n110_adj_4843), 
            .I3(GND_net), .O(n17545[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5188_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5188_2 (.CI(GND_net), .I0(n41_adj_4842), .I1(n110_adj_4843), 
            .CO(n39092));
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_17_lut (.I0(GND_net), .I1(n13369[14]), .I2(GND_net), 
            .I3(n39298), .O(n12529[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_5_lut (.I0(GND_net), .I1(n16224[2]), .I2(n314), .I3(n39439), 
            .O(n15713[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_17 (.CI(n39298), .I0(n13369[14]), .I1(GND_net), 
            .CO(n39299));
    SB_LUT4 add_4909_16_lut (.I0(GND_net), .I1(n13369[13]), .I2(n1105), 
            .I3(n39297), .O(n12529[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_16 (.CI(n39297), .I0(n13369[13]), .I1(n1105), .CO(n39298));
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4845));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_15_lut (.I0(GND_net), .I1(n13369[12]), .I2(n1032), 
            .I3(n39296), .O(n12529[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5069_5 (.CI(n39439), .I0(n16224[2]), .I1(n314), .CO(n39440));
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4846));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4909_15 (.CI(n39296), .I0(n13369[12]), .I1(n1032), .CO(n39297));
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_14_lut (.I0(GND_net), .I1(n13369[11]), .I2(n959), 
            .I3(n39295), .O(n12529[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_4_lut (.I0(GND_net), .I1(n16224[1]), .I2(n241), .I3(n39438), 
            .O(n15713[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n38357), .I0(GND_net), .I1(n1_adj_5146[1]), 
            .CO(n38358));
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4847));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4909_14 (.CI(n39295), .I0(n13369[11]), .I1(n959), .CO(n39296));
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4848));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4849));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5146[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3723 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4851));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5146[0]), 
            .CO(n38357));
    SB_CARRY add_12_14 (.CI(n38253), .I0(n106[12]), .I1(n155[12]), .CO(n38254));
    SB_CARRY add_5069_4 (.CI(n39438), .I0(n16224[1]), .I1(n241), .CO(n39439));
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n38252), .O(duty_23__N_3772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n38356), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n38252), .I0(n106[11]), .I1(n155[11]), .CO(n38253));
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n38355), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n38355), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n38356));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n38354), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n38251), .O(duty_23__N_3772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n38251), .I0(n106[10]), .I1(n155[10]), .CO(n38252));
    SB_CARRY sub_3_add_2_23 (.CI(n38354), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n38355));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n38250), 
            .O(duty_23__N_3772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5069_3_lut (.I0(GND_net), .I1(n16224[0]), .I2(n168), .I3(n39437), 
            .O(n15713[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_3 (.CI(n39437), .I0(n16224[0]), .I1(n168), .CO(n39438));
    SB_LUT4 add_5069_2_lut (.I0(GND_net), .I1(n26_adj_4789), .I2(n95), 
            .I3(GND_net), .O(n15713[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5069_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5069_2 (.CI(GND_net), .I0(n26_adj_4789), .I1(n95), .CO(n39437));
    SB_LUT4 add_4909_13_lut (.I0(GND_net), .I1(n13369[10]), .I2(n886), 
            .I3(n39294), .O(n12529[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_13 (.CI(n39294), .I0(n13369[10]), .I1(n886), .CO(n39295));
    SB_LUT4 add_4909_12_lut (.I0(GND_net), .I1(n13369[9]), .I2(n813), 
            .I3(n39293), .O(n12529[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n38353), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3772[1]), .I1(n257[1]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3747[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3772[2]), .I1(n257[2]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3747[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3747[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3747[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3747[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3747[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3747[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3747[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3747[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3747[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3747[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3747[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3747[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4843));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4842));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3747[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3747[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3747[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4832));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3747[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3747[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_22 (.CI(n38353), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n38354));
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n38352), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n38352), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n38353));
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3747[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5099_16_lut (.I0(GND_net), .I1(n16673[13]), .I2(n1120), 
            .I3(n39436), .O(n16224[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3747[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n38351), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3747[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4909_12 (.CI(n39293), .I0(n13369[9]), .I1(n813), .CO(n39294));
    SB_CARRY sub_3_add_2_20 (.CI(n38351), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n38352));
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3747[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3772[23]), .I1(n257[23]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3747[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n38350), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_15_lut (.I0(GND_net), .I1(n16673[12]), .I2(n1047), 
            .I3(n39435), .O(n16224[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_15 (.CI(n39435), .I0(n16673[12]), .I1(n1047), .CO(n39436));
    SB_LUT4 add_4909_11_lut (.I0(GND_net), .I1(n13369[8]), .I2(n740), 
            .I3(n39292), .O(n12529[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n38350), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n38351));
    SB_CARRY add_4909_11 (.CI(n39292), .I0(n13369[8]), .I1(n740), .CO(n39293));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n38349), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_18 (.CI(n38349), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n38350));
    SB_LUT4 add_5099_14_lut (.I0(GND_net), .I1(n16673[11]), .I2(n974), 
            .I3(n39434), .O(n16224[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n38348), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n38348), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n38349));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n38347), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n38347), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n38348));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n38346), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n38250), .I0(n106[9]), .I1(n155[9]), .CO(n38251));
    SB_CARRY sub_3_add_2_15 (.CI(n38346), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n38347));
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n38345), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4909_10_lut (.I0(GND_net), .I1(n13369[7]), .I2(n667), 
            .I3(n39291), .O(n12529[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_10 (.CI(n39291), .I0(n13369[7]), .I1(n667), .CO(n39292));
    SB_CARRY add_5099_14 (.CI(n39434), .I0(n16673[11]), .I1(n974), .CO(n39435));
    SB_CARRY sub_3_add_2_14 (.CI(n38345), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n38346));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n38249), 
            .O(duty_23__N_3772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_13_lut (.I0(GND_net), .I1(n16673[10]), .I2(n901), 
            .I3(n39433), .O(n16224[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4909_9_lut (.I0(GND_net), .I1(n13369[6]), .I2(n594), .I3(n39290), 
            .O(n12529[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n38249), .I0(n106[8]), .I1(n155[8]), .CO(n38250));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n38344), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_9 (.CI(n39290), .I0(n13369[6]), .I1(n594), .CO(n39291));
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4859));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_13 (.CI(n38344), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n38345));
    SB_LUT4 add_4909_8_lut (.I0(GND_net), .I1(n13369[5]), .I2(n521), .I3(n39289), 
            .O(n12529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n38343), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_13 (.CI(n39433), .I0(n16673[10]), .I1(n901), .CO(n39434));
    SB_CARRY sub_3_add_2_12 (.CI(n38343), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n38344));
    SB_LUT4 add_5099_12_lut (.I0(GND_net), .I1(n16673[9]), .I2(n828), 
            .I3(n39432), .O(n16224[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_8 (.CI(n39289), .I0(n13369[5]), .I1(n521), .CO(n39290));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n38248), 
            .O(duty_23__N_3772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n38342), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_9 (.CI(n38248), .I0(n106[7]), .I1(n155[7]), .CO(n38249));
    SB_CARRY sub_3_add_2_11 (.CI(n38342), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n38343));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n38341), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5099_12 (.CI(n39432), .I0(n16673[9]), .I1(n828), .CO(n39433));
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4827));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5099_11_lut (.I0(GND_net), .I1(n16673[8]), .I2(n755), 
            .I3(n39431), .O(n16224[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_11 (.CI(n39431), .I0(n16673[8]), .I1(n755), .CO(n39432));
    SB_LUT4 add_4909_7_lut (.I0(GND_net), .I1(n13369[4]), .I2(n448), .I3(n39288), 
            .O(n12529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_7 (.CI(n39288), .I0(n13369[4]), .I1(n448), .CO(n39289));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n38247), 
            .O(duty_23__N_3772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4909_6_lut (.I0(GND_net), .I1(n13369[3]), .I2(n375), .I3(n39287), 
            .O(n12529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n38341), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n38342));
    SB_LUT4 add_5099_10_lut (.I0(GND_net), .I1(n16673[7]), .I2(n682), 
            .I3(n39430), .O(n16224[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4909_6 (.CI(n39287), .I0(n13369[3]), .I1(n375), .CO(n39288));
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4826));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4824));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5099_10 (.CI(n39430), .I0(n16673[7]), .I1(n682), .CO(n39431));
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5099_9_lut (.I0(GND_net), .I1(n16673[6]), .I2(n609), .I3(n39429), 
            .O(n16224[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4823));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_5_lut (.I0(GND_net), .I1(n13369[2]), .I2(n302), .I3(n39286), 
            .O(n12529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_5_lut (.I0(GND_net), .I1(n18513[2]), .I2(n341_adj_4780), 
            .I3(n39163), .O(n18416[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n38340), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n38340), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n38341));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n38339), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n38339), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n38340));
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4862));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4863));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4864));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5099_9 (.CI(n39429), .I0(n16673[6]), .I1(n609), .CO(n39430));
    SB_CARRY add_4909_5 (.CI(n39286), .I0(n13369[2]), .I1(n302), .CO(n39287));
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n38338), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_7 (.CI(n38338), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n38339));
    SB_LUT4 add_5099_8_lut (.I0(GND_net), .I1(n16673[5]), .I2(n536), .I3(n39428), 
            .O(n16224[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4909_4_lut (.I0(GND_net), .I1(n13369[1]), .I2(n229), .I3(n39285), 
            .O(n12529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_4 (.CI(n39285), .I0(n13369[1]), .I1(n229), .CO(n39286));
    SB_LUT4 add_4909_3_lut (.I0(GND_net), .I1(n13369[0]), .I2(n156), .I3(n39284), 
            .O(n12529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4909_3 (.CI(n39284), .I0(n13369[0]), .I1(n156), .CO(n39285));
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_8 (.CI(n38247), .I0(n106[6]), .I1(n155[6]), .CO(n38248));
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4866));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n38337), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n38246), 
            .O(duty_23__N_3772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n38337), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n38338));
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4909_2_lut (.I0(GND_net), .I1(n14_adj_4774), .I2(n83), 
            .I3(GND_net), .O(n12529[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4909_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n38246), .I0(n106[5]), .I1(n155[5]), .CO(n38247));
    SB_CARRY add_5099_8 (.CI(n39428), .I0(n16673[5]), .I1(n536), .CO(n39429));
    SB_CARRY add_4909_2 (.CI(GND_net), .I0(n14_adj_4774), .I1(n83), .CO(n39284));
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4818));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4869));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n38336), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5219_11_lut (.I0(GND_net), .I1(n18128[8]), .I2(n770), 
            .I3(n39283), .O(n17929[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_7_lut (.I0(GND_net), .I1(n16673[4]), .I2(n463), .I3(n39427), 
            .O(n16224[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_7 (.CI(n39427), .I0(n16673[4]), .I1(n463), .CO(n39428));
    SB_LUT4 add_5219_10_lut (.I0(GND_net), .I1(n18128[7]), .I2(n697), 
            .I3(n39282), .O(n17929[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n38336), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n38337));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n38245), 
            .O(duty_23__N_3772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_6_lut (.I0(GND_net), .I1(n16673[3]), .I2(n390), .I3(n39426), 
            .O(n16224[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_10 (.CI(n39282), .I0(n18128[7]), .I1(n697), .CO(n39283));
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5219_9_lut (.I0(GND_net), .I1(n18128[6]), .I2(n624), .I3(n39281), 
            .O(n17929[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n38335), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n38245), .I0(n106[4]), .I1(n155[4]), .CO(n38246));
    SB_CARRY sub_3_add_2_4 (.CI(n38335), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n38336));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n38334), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n38244), 
            .O(duty_23__N_3772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5099_6 (.CI(n39426), .I0(n16673[3]), .I1(n390), .CO(n39427));
    SB_CARRY add_5219_9 (.CI(n39281), .I0(n18128[6]), .I1(n624), .CO(n39282));
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5219_8_lut (.I0(GND_net), .I1(n18128[5]), .I2(n551), .I3(n39280), 
            .O(n17929[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_5_lut (.I0(GND_net), .I1(n16673[2]), .I2(n317), .I3(n39425), 
            .O(n16224[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4874));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_5 (.CI(n38244), .I0(n106[3]), .I1(n155[3]), .CO(n38245));
    SB_CARRY add_5219_8 (.CI(n39280), .I0(n18128[5]), .I1(n551), .CO(n39281));
    SB_CARRY sub_3_add_2_3 (.CI(n38334), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n38335));
    SB_CARRY add_5099_5 (.CI(n39425), .I0(n16673[2]), .I1(n317), .CO(n39426));
    SB_LUT4 add_5219_7_lut (.I0(GND_net), .I1(n18128[4]), .I2(n478), .I3(n39279), 
            .O(n17929[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n38243), 
            .O(duty_23__N_3772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5099_4_lut (.I0(GND_net), .I1(n16673[1]), .I2(n244), .I3(n39424), 
            .O(n16224[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_7 (.CI(n39279), .I0(n18128[4]), .I1(n478), .CO(n39280));
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_4 (.CI(n38243), .I0(n106[2]), .I1(n155[2]), .CO(n38244));
    SB_CARRY add_5099_4 (.CI(n39424), .I0(n16673[1]), .I1(n244), .CO(n39425));
    SB_LUT4 add_5219_6_lut (.I0(GND_net), .I1(n18128[3]), .I2(n405), .I3(n39278), 
            .O(n17929[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4876));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4878));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4879));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5219_6 (.CI(n39278), .I0(n18128[3]), .I1(n405), .CO(n39279));
    SB_LUT4 add_5099_3_lut (.I0(GND_net), .I1(n16673[0]), .I2(n171), .I3(n39423), 
            .O(n16224[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n38334));
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4881));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n38242), 
            .O(duty_23__N_3772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5219_5_lut (.I0(GND_net), .I1(n18128[2]), .I2(n332), .I3(n39277), 
            .O(n17929[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_3 (.CI(n38242), .I0(n106[1]), .I1(n155[1]), .CO(n38243));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5219_5 (.CI(n39277), .I0(n18128[2]), .I1(n332), .CO(n39278));
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n38242));
    SB_LUT4 add_5219_4_lut (.I0(GND_net), .I1(n18128[1]), .I2(n259), .I3(n39276), 
            .O(n17929[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5099_3 (.CI(n39423), .I0(n16673[0]), .I1(n171), .CO(n39424));
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4885));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5099_2_lut (.I0(GND_net), .I1(n29_adj_4744), .I2(n98), 
            .I3(GND_net), .O(n16224[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5099_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_4 (.CI(n39276), .I0(n18128[1]), .I1(n259), .CO(n39277));
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4806));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4805));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5099_2 (.CI(GND_net), .I0(n29_adj_4744), .I1(n98), .CO(n39423));
    SB_LUT4 add_5219_3_lut (.I0(GND_net), .I1(n18128[0]), .I2(n186), .I3(n39275), 
            .O(n17929[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_3 (.CI(n39275), .I0(n18128[0]), .I1(n186), .CO(n39276));
    SB_LUT4 add_5260_8_lut (.I0(GND_net), .I1(n18465[5]), .I2(n560), .I3(n39422), 
            .O(n18353[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5260_7_lut (.I0(GND_net), .I1(n18465[4]), .I2(n487), .I3(n39421), 
            .O(n18353[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_7 (.CI(n39421), .I0(n18465[4]), .I1(n487), .CO(n39422));
    SB_LUT4 add_5219_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n17929[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5260_6_lut (.I0(GND_net), .I1(n18465[3]), .I2(n414), .I3(n39420), 
            .O(n18353[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n39275));
    SB_CARRY add_5260_6 (.CI(n39420), .I0(n18465[3]), .I1(n414), .CO(n39421));
    SB_LUT4 add_4948_20_lut (.I0(GND_net), .I1(n14129[17]), .I2(GND_net), 
            .I3(n39274), .O(n13369[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4948_19_lut (.I0(GND_net), .I1(n14129[16]), .I2(GND_net), 
            .I3(n39273), .O(n13369[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_19 (.CI(n39273), .I0(n14129[16]), .I1(GND_net), 
            .CO(n39274));
    SB_LUT4 add_5260_5_lut (.I0(GND_net), .I1(n18465[2]), .I2(n341), .I3(n39419), 
            .O(n18353[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_5 (.CI(n39419), .I0(n18465[2]), .I1(n341), .CO(n39420));
    SB_LUT4 add_4948_18_lut (.I0(GND_net), .I1(n14129[15]), .I2(GND_net), 
            .I3(n39272), .O(n13369[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_18 (.CI(n39272), .I0(n14129[15]), .I1(GND_net), 
            .CO(n39273));
    SB_LUT4 add_4948_17_lut (.I0(GND_net), .I1(n14129[14]), .I2(GND_net), 
            .I3(n39271), .O(n13369[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5260_4_lut (.I0(GND_net), .I1(n18465[1]), .I2(n268_adj_4889), 
            .I3(n39418), .O(n18353[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_4 (.CI(n39418), .I0(n18465[1]), .I1(n268_adj_4889), 
            .CO(n39419));
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4803));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5260_3_lut (.I0(GND_net), .I1(n18465[0]), .I2(n195_adj_4890), 
            .I3(n39417), .O(n18353[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4802));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5260_3 (.CI(n39417), .I0(n18465[0]), .I1(n195_adj_4890), 
            .CO(n39418));
    SB_LUT4 add_5260_2_lut (.I0(GND_net), .I1(n53_adj_4891), .I2(n122_adj_4892), 
            .I3(GND_net), .O(n18353[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5260_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_17 (.CI(n39271), .I0(n14129[14]), .I1(GND_net), 
            .CO(n39272));
    SB_LUT4 add_4948_16_lut (.I0(GND_net), .I1(n14129[13]), .I2(n1108), 
            .I3(n39270), .O(n13369[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5260_2 (.CI(GND_net), .I0(n53_adj_4891), .I1(n122_adj_4892), 
            .CO(n39417));
    SB_LUT4 add_5127_15_lut (.I0(GND_net), .I1(n17064[12]), .I2(n1050_adj_4893), 
            .I3(n39416), .O(n16673[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_16 (.CI(n39270), .I0(n14129[13]), .I1(n1108), .CO(n39271));
    SB_LUT4 add_5127_14_lut (.I0(GND_net), .I1(n17064[11]), .I2(n977_adj_4894), 
            .I3(n39415), .O(n16673[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4948_15_lut (.I0(GND_net), .I1(n14129[12]), .I2(n1035), 
            .I3(n39269), .O(n13369[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_15 (.CI(n39269), .I0(n14129[12]), .I1(n1035), .CO(n39270));
    SB_CARRY add_5127_14 (.CI(n39415), .I0(n17064[11]), .I1(n977_adj_4894), 
            .CO(n39416));
    SB_LUT4 add_4948_14_lut (.I0(GND_net), .I1(n14129[11]), .I2(n962), 
            .I3(n39268), .O(n13369[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_13_lut (.I0(GND_net), .I1(n17064[10]), .I2(n904), 
            .I3(n39414), .O(n16673[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_14 (.CI(n39268), .I0(n14129[11]), .I1(n962), .CO(n39269));
    SB_LUT4 add_4948_13_lut (.I0(GND_net), .I1(n14129[10]), .I2(n889), 
            .I3(n39267), .O(n13369[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_13 (.CI(n39267), .I0(n14129[10]), .I1(n889), .CO(n39268));
    SB_LUT4 add_4948_12_lut (.I0(GND_net), .I1(n14129[9]), .I2(n816), 
            .I3(n39266), .O(n13369[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_12 (.CI(n39266), .I0(n14129[9]), .I1(n816), .CO(n39267));
    SB_CARRY add_5127_13 (.CI(n39414), .I0(n17064[10]), .I1(n904), .CO(n39415));
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4738));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4736));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4948_11_lut (.I0(GND_net), .I1(n14129[8]), .I2(n743), 
            .I3(n39265), .O(n13369[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_12_lut (.I0(GND_net), .I1(n17064[9]), .I2(n831_adj_4787), 
            .I3(n39413), .O(n16673[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_11 (.CI(n39265), .I0(n14129[8]), .I1(n743), .CO(n39266));
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4948_10_lut (.I0(GND_net), .I1(n14129[7]), .I2(n670), 
            .I3(n39264), .O(n13369[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_10 (.CI(n39264), .I0(n14129[7]), .I1(n670), .CO(n39265));
    SB_CARRY add_5127_12 (.CI(n39413), .I0(n17064[9]), .I1(n831_adj_4787), 
            .CO(n39414));
    SB_LUT4 add_5127_11_lut (.I0(GND_net), .I1(n17064[8]), .I2(n758_adj_4778), 
            .I3(n39412), .O(n16673[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4948_9_lut (.I0(GND_net), .I1(n14129[6]), .I2(n597), .I3(n39263), 
            .O(n13369[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_9 (.CI(n39263), .I0(n14129[6]), .I1(n597), .CO(n39264));
    SB_CARRY add_5127_11 (.CI(n39412), .I0(n17064[8]), .I1(n758_adj_4778), 
            .CO(n39413));
    SB_LUT4 add_4948_8_lut (.I0(GND_net), .I1(n14129[5]), .I2(n524), .I3(n39262), 
            .O(n13369[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_8 (.CI(n39262), .I0(n14129[5]), .I1(n524), .CO(n39263));
    SB_LUT4 add_4948_7_lut (.I0(GND_net), .I1(n14129[4]), .I2(n451), .I3(n39261), 
            .O(n13369[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_10_lut (.I0(GND_net), .I1(n17064[7]), .I2(n685_adj_4775), 
            .I3(n39411), .O(n16673[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_7 (.CI(n39261), .I0(n14129[4]), .I1(n451), .CO(n39262));
    SB_CARRY add_5127_10 (.CI(n39411), .I0(n17064[7]), .I1(n685_adj_4775), 
            .CO(n39412));
    SB_LUT4 add_4948_6_lut (.I0(GND_net), .I1(n14129[3]), .I2(n378), .I3(n39260), 
            .O(n13369[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_6 (.CI(n39260), .I0(n14129[3]), .I1(n378), .CO(n39261));
    SB_LUT4 add_5127_9_lut (.I0(GND_net), .I1(n17064[6]), .I2(n612_adj_4773), 
            .I3(n39410), .O(n16673[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4897));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32359_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(PWMLimit[2]), .O(n47440));   // verilog/motorControl.v(36[10:25])
    defparam i32359_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4901));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(GND_net), .O(n6_adj_4902));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_4948_5_lut (.I0(GND_net), .I1(n14129[2]), .I2(n305), .I3(n39259), 
            .O(n13369[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_5 (.CI(n39259), .I0(n14129[2]), .I1(n305), .CO(n39260));
    SB_CARRY add_5127_9 (.CI(n39410), .I0(n17064[6]), .I1(n612_adj_4773), 
            .CO(n39411));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4903));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4948_4_lut (.I0(GND_net), .I1(n14129[1]), .I2(n232), .I3(n39258), 
            .O(n13369[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4948_4 (.CI(n39258), .I0(n14129[1]), .I1(n232), .CO(n39259));
    SB_LUT4 add_5127_8_lut (.I0(GND_net), .I1(n17064[5]), .I2(n539_adj_4763), 
            .I3(n39409), .O(n16673[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4905));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32325_3_lut_4_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3772[2]), .O(n47406));   // verilog/motorControl.v(38[19:35])
    defparam i32325_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4906));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4908));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4948_3_lut (.I0(GND_net), .I1(n14129[0]), .I2(n159), .I3(n39257), 
            .O(n13369[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_8 (.CI(n39409), .I0(n17064[5]), .I1(n539_adj_4763), 
            .CO(n39410));
    SB_CARRY add_4948_3 (.CI(n39257), .I0(n14129[0]), .I1(n159), .CO(n39258));
    SB_LUT4 add_4948_2_lut (.I0(GND_net), .I1(n17_adj_4762), .I2(n86), 
            .I3(GND_net), .O(n13369[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4948_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_7_lut (.I0(GND_net), .I1(n17064[4]), .I2(n466_adj_4760), 
            .I3(n39408), .O(n16673[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4909));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4911));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4948_2 (.CI(GND_net), .I0(n17_adj_4762), .I1(n86), .CO(n39257));
    SB_LUT4 add_4985_19_lut (.I0(GND_net), .I1(n14813[16]), .I2(GND_net), 
            .I3(n39256), .O(n14129[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4912));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4913));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4914));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4915));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4916));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5127_7 (.CI(n39408), .I0(n17064[4]), .I1(n466_adj_4760), 
            .CO(n39409));
    SB_LUT4 add_5127_6_lut (.I0(GND_net), .I1(n17064[3]), .I2(n393_adj_4746), 
            .I3(n39407), .O(n16673[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_6 (.CI(n39407), .I0(n17064[3]), .I1(n393_adj_4746), 
            .CO(n39408));
    SB_LUT4 add_4985_18_lut (.I0(GND_net), .I1(n14813[15]), .I2(GND_net), 
            .I3(n39255), .O(n14129[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_18 (.CI(n39255), .I0(n14813[15]), .I1(GND_net), 
            .CO(n39256));
    SB_LUT4 add_4985_17_lut (.I0(GND_net), .I1(n14813[14]), .I2(GND_net), 
            .I3(n39254), .O(n14129[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_5_lut (.I0(GND_net), .I1(n17064[2]), .I2(n320_adj_4745), 
            .I3(n39406), .O(n16673[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4917));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4918));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4919));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4920));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5127_5 (.CI(n39406), .I0(n17064[2]), .I1(n320_adj_4745), 
            .CO(n39407));
    SB_CARRY add_4985_17 (.CI(n39254), .I0(n14813[14]), .I1(GND_net), 
            .CO(n39255));
    SB_LUT4 add_5127_4_lut (.I0(GND_net), .I1(n17064[1]), .I2(n247), .I3(n39405), 
            .O(n16673[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_4 (.CI(n39405), .I0(n17064[1]), .I1(n247), .CO(n39406));
    SB_LUT4 add_4985_16_lut (.I0(GND_net), .I1(n14813[13]), .I2(n1111), 
            .I3(n39253), .O(n14129[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_3_lut (.I0(GND_net), .I1(n17064[0]), .I2(n174), .I3(n39404), 
            .O(n16673[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_16 (.CI(n39253), .I0(n14813[13]), .I1(n1111), .CO(n39254));
    SB_CARRY add_5127_3 (.CI(n39404), .I0(n17064[0]), .I1(n174), .CO(n39405));
    SB_LUT4 add_5127_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n16673[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4921));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4922));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5127_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n39404));
    SB_LUT4 add_5153_14_lut (.I0(GND_net), .I1(n17401[11]), .I2(n980_adj_4817), 
            .I3(n39403), .O(n17064[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_15_lut (.I0(GND_net), .I1(n14813[12]), .I2(n1038), 
            .I3(n39252), .O(n14129[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_13_lut (.I0(GND_net), .I1(n17401[10]), .I2(n907_adj_4812), 
            .I3(n39402), .O(n17064[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_13 (.CI(n39402), .I0(n17401[10]), .I1(n907_adj_4812), 
            .CO(n39403));
    SB_CARRY add_4985_15 (.CI(n39252), .I0(n14813[12]), .I1(n1038), .CO(n39253));
    SB_LUT4 add_5153_12_lut (.I0(GND_net), .I1(n17401[9]), .I2(n834_adj_4791), 
            .I3(n39401), .O(n17064[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_12 (.CI(n39401), .I0(n17401[9]), .I1(n834_adj_4791), 
            .CO(n39402));
    SB_LUT4 add_5153_11_lut (.I0(GND_net), .I1(n17401[8]), .I2(n761_adj_4790), 
            .I3(n39400), .O(n17064[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_14_lut (.I0(GND_net), .I1(n14813[11]), .I2(n965), 
            .I3(n39251), .O(n14129[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_14 (.CI(n39251), .I0(n14813[11]), .I1(n965), .CO(n39252));
    SB_CARRY add_5153_11 (.CI(n39400), .I0(n17401[8]), .I1(n761_adj_4790), 
            .CO(n39401));
    SB_LUT4 add_4985_13_lut (.I0(GND_net), .I1(n14813[10]), .I2(n892), 
            .I3(n39250), .O(n14129[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_10_lut (.I0(GND_net), .I1(n17401[7]), .I2(n688_adj_4785), 
            .I3(n39399), .O(n17064[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_13 (.CI(n39250), .I0(n14813[10]), .I1(n892), .CO(n39251));
    SB_CARRY add_5153_10 (.CI(n39399), .I0(n17401[7]), .I1(n688_adj_4785), 
            .CO(n39400));
    SB_LUT4 add_5153_9_lut (.I0(GND_net), .I1(n17401[6]), .I2(n615_adj_4782), 
            .I3(n39398), .O(n17064[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_12_lut (.I0(GND_net), .I1(n14813[9]), .I2(n819), 
            .I3(n39249), .O(n14129[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_9 (.CI(n39398), .I0(n17401[6]), .I1(n615_adj_4782), 
            .CO(n39399));
    SB_CARRY add_4985_12 (.CI(n39249), .I0(n14813[9]), .I1(n819), .CO(n39250));
    SB_LUT4 add_5153_8_lut (.I0(GND_net), .I1(n17401[5]), .I2(n542_adj_4766), 
            .I3(n39397), .O(n17064[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_8 (.CI(n39397), .I0(n17401[5]), .I1(n542_adj_4766), 
            .CO(n39398));
    SB_LUT4 add_5153_7_lut (.I0(GND_net), .I1(n17401[4]), .I2(n469_adj_4761), 
            .I3(n39396), .O(n17064[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_7 (.CI(n39396), .I0(n17401[4]), .I1(n469_adj_4761), 
            .CO(n39397));
    SB_LUT4 add_4985_11_lut (.I0(GND_net), .I1(n14813[8]), .I2(n746), 
            .I3(n39248), .O(n14129[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20332_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20332_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5153_6_lut (.I0(GND_net), .I1(n17401[3]), .I2(n396_adj_4758), 
            .I3(n39395), .O(n17064[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_6 (.CI(n39395), .I0(n17401[3]), .I1(n396_adj_4758), 
            .CO(n39396));
    SB_LUT4 add_5153_5_lut (.I0(GND_net), .I1(n17401[2]), .I2(n323_adj_4757), 
            .I3(n39394), .O(n17064[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_5 (.CI(n39394), .I0(n17401[2]), .I1(n323_adj_4757), 
            .CO(n39395));
    SB_CARRY add_4985_11 (.CI(n39248), .I0(n14813[8]), .I1(n746), .CO(n39249));
    SB_LUT4 add_4985_10_lut (.I0(GND_net), .I1(n14813[7]), .I2(n673), 
            .I3(n39247), .O(n14129[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4923));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4924));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4925));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4926));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4985_10 (.CI(n39247), .I0(n14813[7]), .I1(n673), .CO(n39248));
    SB_LUT4 add_5153_4_lut (.I0(GND_net), .I1(n17401[1]), .I2(n250_adj_4755), 
            .I3(n39393), .O(n17064[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_9_lut (.I0(GND_net), .I1(n14813[6]), .I2(n600), .I3(n39246), 
            .O(n14129[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_9 (.CI(n39246), .I0(n14813[6]), .I1(n600), .CO(n39247));
    SB_CARRY add_5153_4 (.CI(n39393), .I0(n17401[1]), .I1(n250_adj_4755), 
            .CO(n39394));
    SB_LUT4 add_5153_3_lut (.I0(GND_net), .I1(n17401[0]), .I2(n177_adj_4741), 
            .I3(n39392), .O(n17064[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4927));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5153_3 (.CI(n39392), .I0(n17401[0]), .I1(n177_adj_4741), 
            .CO(n39393));
    SB_LUT4 add_4985_8_lut (.I0(GND_net), .I1(n14813[5]), .I2(n527), .I3(n39245), 
            .O(n14129[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_8 (.CI(n39245), .I0(n14813[5]), .I1(n527), .CO(n39246));
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4928));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4985_7_lut (.I0(GND_net), .I1(n14813[4]), .I2(n454), .I3(n39244), 
            .O(n14129[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_2_lut (.I0(GND_net), .I1(n35_adj_4740), .I2(n104_adj_4737), 
            .I3(GND_net), .O(n17064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_7 (.CI(n39244), .I0(n14813[4]), .I1(n454), .CO(n39245));
    SB_CARRY add_5153_2 (.CI(GND_net), .I0(n35_adj_4740), .I1(n104_adj_4737), 
            .CO(n39392));
    SB_LUT4 add_4985_6_lut (.I0(GND_net), .I1(n14813[3]), .I2(n381), .I3(n39243), 
            .O(n14129[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5273_7_lut (.I0(GND_net), .I1(n44653), .I2(n490_adj_4929), 
            .I3(n39391), .O(n18465[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4930));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5273_6_lut (.I0(GND_net), .I1(n18549[3]), .I2(n417_adj_4931), 
            .I3(n39390), .O(n18465[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_6 (.CI(n39243), .I0(n14813[3]), .I1(n381), .CO(n39244));
    SB_CARRY add_5273_6 (.CI(n39390), .I0(n18549[3]), .I1(n417_adj_4931), 
            .CO(n39391));
    SB_CARRY add_5267_5 (.CI(n39163), .I0(n18513[2]), .I1(n341_adj_4780), 
            .CO(n39164));
    SB_LUT4 add_4985_5_lut (.I0(GND_net), .I1(n14813[2]), .I2(n308_adj_4932), 
            .I3(n39242), .O(n14129[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5267_4_lut (.I0(GND_net), .I1(n18513[1]), .I2(n268_adj_4933), 
            .I3(n39162), .O(n18416[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5267_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_5 (.CI(n39242), .I0(n14813[2]), .I1(n308_adj_4932), 
            .CO(n39243));
    SB_LUT4 add_5273_5_lut (.I0(GND_net), .I1(n18549[2]), .I2(n344_adj_4930), 
            .I3(n39389), .O(n18465[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_5 (.CI(n39389), .I0(n18549[2]), .I1(n344_adj_4930), 
            .CO(n39390));
    SB_CARRY add_5267_4 (.CI(n39162), .I0(n18513[1]), .I1(n268_adj_4933), 
            .CO(n39163));
    SB_LUT4 add_5273_4_lut (.I0(GND_net), .I1(n18549[1]), .I2(n271_adj_4928), 
            .I3(n39388), .O(n18465[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_4 (.CI(n39388), .I0(n18549[1]), .I1(n271_adj_4928), 
            .CO(n39389));
    SB_LUT4 add_4985_4_lut (.I0(GND_net), .I1(n14813[1]), .I2(n235_adj_4927), 
            .I3(n39241), .O(n14129[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5273_3_lut (.I0(GND_net), .I1(n18549[0]), .I2(n198_adj_4926), 
            .I3(n39387), .O(n18465[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_4 (.CI(n39241), .I0(n14813[1]), .I1(n235_adj_4927), 
            .CO(n39242));
    SB_CARRY add_5273_3 (.CI(n39387), .I0(n18549[0]), .I1(n198_adj_4926), 
            .CO(n39388));
    SB_LUT4 add_5273_2_lut (.I0(GND_net), .I1(n56_adj_4925), .I2(n125_adj_4924), 
            .I3(GND_net), .O(n18465[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5273_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_3_lut (.I0(GND_net), .I1(n14813[0]), .I2(n162_adj_4923), 
            .I3(n39240), .O(n14129[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5273_2 (.CI(GND_net), .I0(n56_adj_4925), .I1(n125_adj_4924), 
            .CO(n39387));
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4933));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4932));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4985_3 (.CI(n39240), .I0(n14813[0]), .I1(n162_adj_4923), 
            .CO(n39241));
    SB_LUT4 add_5177_13_lut (.I0(GND_net), .I1(n17688[10]), .I2(n910_adj_4879), 
            .I3(n39386), .O(n17401[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4985_2_lut (.I0(GND_net), .I1(n20_adj_4878), .I2(n89_adj_4877), 
            .I3(GND_net), .O(n14129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4985_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4985_2 (.CI(GND_net), .I0(n20_adj_4878), .I1(n89_adj_4877), 
            .CO(n39240));
    SB_LUT4 add_5177_12_lut (.I0(GND_net), .I1(n17688[9]), .I2(n837_adj_4876), 
            .I3(n39385), .O(n17401[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24448_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n4_adj_4935), .I3(n18609[1]), .O(n6_adj_4936));   // verilog/motorControl.v(34[25:36])
    defparam i24448_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3648[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3648[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3648[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3648[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3648[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3648[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3648[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3648[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3648[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3648[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3648[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3648[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3648[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3648[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3648[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3648[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3648[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3648[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3648[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3648[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3648[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3648[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3648[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n18609[1]), .I3(n4_adj_4935), .O(n18549[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 add_5237_10_lut (.I0(GND_net), .I1(n18289[7]), .I2(n700), 
            .I3(n39239), .O(n18128[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5177_12 (.CI(n39385), .I0(n17688[9]), .I1(n837_adj_4876), 
            .CO(n39386));
    SB_LUT4 add_5177_11_lut (.I0(GND_net), .I1(n17688[8]), .I2(n764_adj_4851), 
            .I3(n39384), .O(n17401[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5237_9_lut (.I0(GND_net), .I1(n18289[6]), .I2(n627), .I3(n39238), 
            .O(n18128[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_9 (.CI(n39238), .I0(n18289[6]), .I1(n627), .CO(n39239));
    SB_CARRY add_5177_11 (.CI(n39384), .I0(n17688[8]), .I1(n764_adj_4851), 
            .CO(n39385));
    SB_LUT4 add_5177_10_lut (.I0(GND_net), .I1(n17688[7]), .I2(n691_adj_4849), 
            .I3(n39383), .O(n17401[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5237_8_lut (.I0(GND_net), .I1(n18289[5]), .I2(n554), .I3(n39237), 
            .O(n18128[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_8 (.CI(n39237), .I0(n18289[5]), .I1(n554), .CO(n39238));
    SB_LUT4 add_5237_7_lut (.I0(GND_net), .I1(n18289[4]), .I2(n481), .I3(n39236), 
            .O(n18128[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_7 (.CI(n39236), .I0(n18289[4]), .I1(n481), .CO(n39237));
    SB_LUT4 add_5237_6_lut (.I0(GND_net), .I1(n18289[3]), .I2(n408), .I3(n39235), 
            .O(n18128[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5177_10 (.CI(n39383), .I0(n17688[7]), .I1(n691_adj_4849), 
            .CO(n39384));
    SB_LUT4 add_5177_9_lut (.I0(GND_net), .I1(n17688[6]), .I2(n618_adj_4848), 
            .I3(n39382), .O(n17401[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5177_9 (.CI(n39382), .I0(n17688[6]), .I1(n618_adj_4848), 
            .CO(n39383));
    SB_CARRY add_5237_6 (.CI(n39235), .I0(n18289[3]), .I1(n408), .CO(n39236));
    SB_LUT4 add_5237_5_lut (.I0(GND_net), .I1(n18289[2]), .I2(n335), .I3(n39234), 
            .O(n18128[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5177_8_lut (.I0(GND_net), .I1(n17688[5]), .I2(n545_adj_4847), 
            .I3(n39381), .O(n17401[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_5 (.CI(n39234), .I0(n18289[2]), .I1(n335), .CO(n39235));
    SB_CARRY add_5177_8 (.CI(n39381), .I0(n17688[5]), .I1(n545_adj_4847), 
            .CO(n39382));
    SB_LUT4 add_5237_4_lut (.I0(GND_net), .I1(n18289[1]), .I2(n262), .I3(n39233), 
            .O(n18128[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_4 (.CI(n39233), .I0(n18289[1]), .I1(n262), .CO(n39234));
    SB_LUT4 add_5177_7_lut (.I0(GND_net), .I1(n17688[4]), .I2(n472_adj_4846), 
            .I3(n39380), .O(n17401[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5177_7 (.CI(n39380), .I0(n17688[4]), .I1(n472_adj_4846), 
            .CO(n39381));
    SB_LUT4 add_5237_3_lut (.I0(GND_net), .I1(n18289[0]), .I2(n189_adj_4845), 
            .I3(n39232), .O(n18128[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_3 (.CI(n39232), .I0(n18289[0]), .I1(n189_adj_4845), 
            .CO(n39233));
    SB_LUT4 add_5237_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18128[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5177_6_lut (.I0(GND_net), .I1(n17688[3]), .I2(n399_adj_4837), 
            .I3(n39379), .O(n17401[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n39232));
    SB_CARRY add_5177_6 (.CI(n39379), .I0(n17688[3]), .I1(n399_adj_4837), 
            .CO(n39380));
    SB_LUT4 add_5177_5_lut (.I0(GND_net), .I1(n17688[2]), .I2(n326_adj_4836), 
            .I3(n39378), .O(n17401[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5177_5 (.CI(n39378), .I0(n17688[2]), .I1(n326_adj_4836), 
            .CO(n39379));
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4937));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i24364_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n37836), .I3(n18673[0]), .O(n4));   // verilog/motorControl.v(34[25:36])
    defparam i24364_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_5177_4_lut (.I0(GND_net), .I1(n17688[1]), .I2(n253_adj_4835), 
            .I3(n39377), .O(n17401[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_18_lut (.I0(GND_net), .I1(n15425[15]), .I2(GND_net), 
            .I3(n39231), .O(n14813[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_17_lut (.I0(GND_net), .I1(n15425[14]), .I2(GND_net), 
            .I3(n39230), .O(n14813[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1553 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n18673[0]), .I3(n37836), .O(n18649[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1553.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1554 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(n18649[0]), .I3(n37877), .O(n18609[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1554.LUT_INIT = 16'h8778;
    SB_LUT4 i24402_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(n37877), .I3(n18649[0]), .O(n4_adj_4938));   // verilog/motorControl.v(34[25:36])
    defparam i24402_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_5177_4 (.CI(n39377), .I0(n17688[1]), .I1(n253_adj_4835), 
            .CO(n39378));
    SB_CARRY add_5020_17 (.CI(n39230), .I0(n15425[14]), .I1(GND_net), 
            .CO(n39231));
    SB_LUT4 add_5177_3_lut (.I0(GND_net), .I1(n17688[0]), .I2(n180_adj_4834), 
            .I3(n39376), .O(n17401[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_16_lut (.I0(GND_net), .I1(n15425[13]), .I2(n1114), 
            .I3(n39229), .O(n14813[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24351_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n18649[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24351_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24353_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n37836));   // verilog/motorControl.v(34[25:36])
    defparam i24353_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_5177_3 (.CI(n39376), .I0(n17688[0]), .I1(n180_adj_4834), 
            .CO(n39377));
    SB_CARRY add_5020_16 (.CI(n39229), .I0(n15425[13]), .I1(n1114), .CO(n39230));
    SB_LUT4 add_5020_15_lut (.I0(GND_net), .I1(n15425[12]), .I2(n1041), 
            .I3(n39228), .O(n14813[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32327_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3772[9]), .O(n47408));
    defparam i32327_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5177_2_lut (.I0(GND_net), .I1(n38_adj_4833), .I2(n107_adj_4831), 
            .I3(GND_net), .O(n17401[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5177_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32337_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3772[7]), .O(n47418));
    defparam i32337_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5020_15 (.CI(n39228), .I0(n15425[12]), .I1(n1041), .CO(n39229));
    SB_CARRY add_5177_2 (.CI(GND_net), .I0(n38_adj_4833), .I1(n107_adj_4831), 
            .CO(n39376));
    SB_LUT4 i32229_2_lut_4_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(duty_23__N_3772[9]), .I3(n257[9]), .O(n47310));
    defparam i32229_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5020_14_lut (.I0(GND_net), .I1(n15425[11]), .I2(n968), 
            .I3(n39227), .O(n14813[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5209_11_lut (.I0(GND_net), .I1(n18029[8]), .I2(n770_adj_4830), 
            .I3(n38434), .O(n17809[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32259_2_lut_4_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(duty_23__N_3772[7]), .I3(n257[7]), .O(n47340));
    defparam i32259_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5209_10_lut (.I0(GND_net), .I1(n18029[7]), .I2(n697_adj_4829), 
            .I3(n38433), .O(n17809[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5199_12_lut (.I0(GND_net), .I1(n17929[9]), .I2(n840_adj_4821), 
            .I3(n39375), .O(n17688[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_14 (.CI(n39227), .I0(n15425[11]), .I1(n968), .CO(n39228));
    SB_LUT4 add_5020_13_lut (.I0(GND_net), .I1(n15425[10]), .I2(n895_adj_4820), 
            .I3(n39226), .O(n14813[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24389_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), .I3(\Ki[1] ), 
            .O(n18609[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24389_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24391_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), .I3(\Ki[1] ), 
            .O(n37877));   // verilog/motorControl.v(34[25:36])
    defparam i24391_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_5209_10 (.CI(n38433), .I0(n18029[7]), .I1(n697_adj_4829), 
            .CO(n38434));
    SB_LUT4 add_5209_9_lut (.I0(GND_net), .I1(n18029[6]), .I2(n624_adj_4816), 
            .I3(n38432), .O(n17809[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_9 (.CI(n38432), .I0(n18029[6]), .I1(n624_adj_4816), 
            .CO(n38433));
    SB_LUT4 add_5199_11_lut (.I0(GND_net), .I1(n17929[8]), .I2(n767), 
            .I3(n39374), .O(n17688[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_13 (.CI(n39226), .I0(n15425[10]), .I1(n895_adj_4820), 
            .CO(n39227));
    SB_LUT4 add_5020_12_lut (.I0(GND_net), .I1(n15425[9]), .I2(n822_adj_4810), 
            .I3(n39225), .O(n14813[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5209_8_lut (.I0(GND_net), .I1(n18029[5]), .I2(n551_adj_4809), 
            .I3(n38431), .O(n17809[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1555 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n18609[0]), .I3(n37918), .O(n18549[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1555.LUT_INIT = 16'h8778;
    SB_CARRY add_5209_8 (.CI(n38431), .I0(n18029[5]), .I1(n551_adj_4809), 
            .CO(n38432));
    SB_LUT4 i24440_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n37918), .I3(n18609[0]), .O(n4_adj_4935));   // verilog/motorControl.v(34[25:36])
    defparam i24440_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i24427_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n18549[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24427_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i24429_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n37918));   // verilog/motorControl.v(34[25:36])
    defparam i24429_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_5199_11 (.CI(n39374), .I0(n17929[8]), .I1(n767), .CO(n39375));
    SB_CARRY add_5020_12 (.CI(n39225), .I0(n15425[9]), .I1(n822_adj_4810), 
            .CO(n39226));
    SB_LUT4 add_5020_11_lut (.I0(GND_net), .I1(n15425[8]), .I2(n749_adj_4808), 
            .I3(n39224), .O(n14813[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5209_7_lut (.I0(GND_net), .I1(n18029[4]), .I2(n478_adj_4807), 
            .I3(n38430), .O(n17809[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_7 (.CI(n38430), .I0(n18029[4]), .I1(n478_adj_4807), 
            .CO(n38431));
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4931));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1556 (.I0(n6_adj_4936), .I1(\Ki[4] ), .I2(n18609[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n18549[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1556.LUT_INIT = 16'h965a;
    SB_LUT4 add_5199_10_lut (.I0(GND_net), .I1(n17929[7]), .I2(n694), 
            .I3(n39373), .O(n17688[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_11 (.CI(n39224), .I0(n15425[8]), .I1(n749_adj_4808), 
            .CO(n39225));
    SB_CARRY add_5199_10 (.CI(n39373), .I0(n17929[7]), .I1(n694), .CO(n39374));
    SB_LUT4 add_5020_10_lut (.I0(GND_net), .I1(n15425[7]), .I2(n676_adj_4801), 
            .I3(n39223), .O(n14813[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5209_6_lut (.I0(GND_net), .I1(n18029[3]), .I2(n405_adj_4799), 
            .I3(n38429), .O(n17809[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_6 (.CI(n38429), .I0(n18029[3]), .I1(n405_adj_4799), 
            .CO(n38430));
    SB_CARRY add_5020_10 (.CI(n39223), .I0(n15425[7]), .I1(n676_adj_4801), 
            .CO(n39224));
    SB_LUT4 add_5209_5_lut (.I0(GND_net), .I1(n18029[2]), .I2(n332_adj_4798), 
            .I3(n38428), .O(n17809[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5199_9_lut (.I0(GND_net), .I1(n17929[6]), .I2(n621), .I3(n39372), 
            .O(n17688[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_9_lut (.I0(GND_net), .I1(n15425[6]), .I2(n603_adj_4797), 
            .I3(n39222), .O(n14813[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_5 (.CI(n38428), .I0(n18029[2]), .I1(n332_adj_4798), 
            .CO(n38429));
    SB_LUT4 add_5209_4_lut (.I0(GND_net), .I1(n18029[1]), .I2(n259_adj_4796), 
            .I3(n38427), .O(n17809[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24534_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n18673[0]));   // verilog/motorControl.v(34[25:36])
    defparam i24534_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_5199_9 (.CI(n39372), .I0(n17929[6]), .I1(n621), .CO(n39373));
    SB_CARRY add_5020_9 (.CI(n39222), .I0(n15425[6]), .I1(n603_adj_4797), 
            .CO(n39223));
    SB_CARRY add_5209_4 (.CI(n38427), .I0(n18029[1]), .I1(n259_adj_4796), 
            .CO(n38428));
    SB_LUT4 add_5209_3_lut (.I0(GND_net), .I1(n18029[0]), .I2(n186_adj_4793), 
            .I3(n38426), .O(n17809[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_8_lut (.I0(GND_net), .I1(n15425[5]), .I2(n530_adj_4792), 
            .I3(n39221), .O(n14813[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4939));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5209_3 (.CI(n38426), .I0(n18029[0]), .I1(n186_adj_4793), 
            .CO(n38427));
    SB_LUT4 i2_4_lut_adj_1557 (.I0(n4_adj_4938), .I1(\Ki[3] ), .I2(n18649[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n18609[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1557.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4940));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4929));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5209_2_lut (.I0(GND_net), .I1(n44_adj_4788), .I2(n113_adj_4786), 
            .I3(GND_net), .O(n17809[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1558 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [20]), .O(n12_adj_4941));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1558.LUT_INIT = 16'h9c50;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4942));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5209_2 (.CI(GND_net), .I0(n44_adj_4788), .I1(n113_adj_4786), 
            .CO(n38426));
    SB_LUT4 i24456_4_lut (.I0(n18609[2]), .I1(\Ki[4] ), .I2(n6_adj_4936), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n8_adj_4943));   // verilog/motorControl.v(34[25:36])
    defparam i24456_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1559 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n11_adj_4944));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1559.LUT_INIT = 16'h6ca0;
    SB_LUT4 i24410_4_lut (.I0(n18649[1]), .I1(\Ki[3] ), .I2(n4_adj_4938), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n6_adj_4945));   // verilog/motorControl.v(34[25:36])
    defparam i24410_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4946));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5199_8_lut (.I0(GND_net), .I1(n17929[5]), .I2(n548), .I3(n39371), 
            .O(n17688[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5199_8 (.CI(n39371), .I0(n17929[5]), .I1(n548), .CO(n39372));
    SB_CARRY add_5020_8 (.CI(n39221), .I0(n15425[5]), .I1(n530_adj_4792), 
            .CO(n39222));
    SB_LUT4 i24536_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n38034));   // verilog/motorControl.v(34[25:36])
    defparam i24536_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4947));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5199_7_lut (.I0(GND_net), .I1(n17929[4]), .I2(n475), .I3(n39370), 
            .O(n17688[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4948));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5199_7 (.CI(n39370), .I0(n17929[4]), .I1(n475), .CO(n39371));
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4949));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5020_7_lut (.I0(GND_net), .I1(n15425[4]), .I2(n457_adj_4783), 
            .I3(n39220), .O(n14813[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4951));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4952));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5199_6_lut (.I0(GND_net), .I1(n17929[3]), .I2(n402), .I3(n39369), 
            .O(n17688[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4954));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4955));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5199_6 (.CI(n39369), .I0(n17929[3]), .I1(n402), .CO(n39370));
    SB_CARRY add_5020_7 (.CI(n39220), .I0(n15425[4]), .I1(n457_adj_4783), 
            .CO(n39221));
    SB_LUT4 add_5199_5_lut (.I0(GND_net), .I1(n17929[2]), .I2(n329), .I3(n39368), 
            .O(n17688[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5020_6_lut (.I0(GND_net), .I1(n15425[3]), .I2(n384_adj_4756), 
            .I3(n39219), .O(n14813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_6 (.CI(n39219), .I0(n15425[3]), .I1(n384_adj_4756), 
            .CO(n39220));
    SB_CARRY add_5199_5 (.CI(n39368), .I0(n17929[2]), .I1(n329), .CO(n39369));
    SB_LUT4 add_5020_5_lut (.I0(GND_net), .I1(n15425[2]), .I2(n311_adj_4754), 
            .I3(n39218), .O(n14813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5199_4_lut (.I0(GND_net), .I1(n17929[1]), .I2(n256), .I3(n39367), 
            .O(n17688[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_5 (.CI(n39218), .I0(n15425[2]), .I1(n311_adj_4754), 
            .CO(n39219));
    SB_LUT4 add_5020_4_lut (.I0(GND_net), .I1(n15425[1]), .I2(n238_adj_4752), 
            .I3(n39217), .O(n14813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5199_4 (.CI(n39367), .I0(n17929[1]), .I1(n256), .CO(n39368));
    SB_LUT4 add_5199_3_lut (.I0(GND_net), .I1(n17929[0]), .I2(n183), .I3(n39366), 
            .O(n17688[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_4 (.CI(n39217), .I0(n15425[1]), .I1(n238_adj_4752), 
            .CO(n39218));
    SB_CARRY add_5199_3 (.CI(n39366), .I0(n17929[0]), .I1(n183), .CO(n39367));
    SB_LUT4 add_5199_2_lut (.I0(GND_net), .I1(n41_adj_4750), .I2(n110), 
            .I3(GND_net), .O(n17688[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5199_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5199_2 (.CI(GND_net), .I0(n41_adj_4750), .I1(n110), .CO(n39366));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I1(n10588[21]), .I2(GND_net), .I3(n39365), .O(n10081[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5020_3_lut (.I0(GND_net), .I1(n15425[0]), .I2(n165_adj_4747), 
            .I3(n39216), .O(n14813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4236[23]), .I3(n38287), .O(\PID_CONTROLLER.integral_23__N_3672 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4236[22]), .I3(n38286), .O(\PID_CONTROLLER.integral_23__N_3672 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_3 (.CI(n39216), .I0(n15425[0]), .I1(n165_adj_4747), 
            .CO(n39217));
    SB_LUT4 add_5020_2_lut (.I0(GND_net), .I1(n23_adj_4957), .I2(n92_adj_4958), 
            .I3(GND_net), .O(n14813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5020_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5020_2 (.CI(GND_net), .I0(n23_adj_4957), .I1(n92_adj_4958), 
            .CO(n39216));
    SB_CARRY add_958_24 (.CI(n38286), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4236[22]), .CO(n38287));
    SB_LUT4 add_5053_17_lut (.I0(GND_net), .I1(n15969[14]), .I2(GND_net), 
            .I3(n39215), .O(n15425[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4236[21]), .I3(n38285), .O(\PID_CONTROLLER.integral_23__N_3672 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_16_lut (.I0(GND_net), .I1(n15969[13]), .I2(n1117_adj_4959), 
            .I3(n39214), .O(n15425[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_16 (.CI(n39214), .I0(n15969[13]), .I1(n1117_adj_4959), 
            .CO(n39215));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10588[20]), .I2(GND_net), 
            .I3(n39364), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_15_lut (.I0(GND_net), .I1(n15969[12]), .I2(n1044_adj_4960), 
            .I3(n39213), .O(n15425[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4961));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_23 (.CI(n39364), .I0(n10588[20]), .I1(GND_net), 
            .CO(n39365));
    SB_CARRY add_958_23 (.CI(n38285), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4236[21]), .CO(n38286));
    SB_LUT4 add_958_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4236[20]), .I3(n38284), .O(\PID_CONTROLLER.integral_23__N_3672 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4963));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5053_15 (.CI(n39213), .I0(n15969[12]), .I1(n1044_adj_4960), 
            .CO(n39214));
    SB_CARRY add_958_22 (.CI(n38284), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4236[20]), .CO(n38285));
    SB_LUT4 add_958_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4236[19]), .I3(n38283), .O(\PID_CONTROLLER.integral_23__N_3672 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_14_lut (.I0(GND_net), .I1(n15969[11]), .I2(n971_adj_4964), 
            .I3(n39212), .O(n15425[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4966));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_21 (.CI(n38283), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4236[19]), .CO(n38284));
    SB_LUT4 add_958_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4236[18]), .I3(n38282), .O(\PID_CONTROLLER.integral_23__N_3672 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_14 (.CI(n39212), .I0(n15969[11]), .I1(n971_adj_4964), 
            .CO(n39213));
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4967));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10588[19]), .I2(GND_net), 
            .I3(n39363), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n39363), .I0(n10588[19]), .I1(GND_net), 
            .CO(n39364));
    SB_LUT4 i20590_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10588[18]), .I2(GND_net), 
            .I3(n39362), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_13_lut (.I0(GND_net), .I1(n15969[10]), .I2(n898_adj_4969), 
            .I3(n39211), .O(n15425[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_20 (.CI(n38282), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4236[18]), .CO(n38283));
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4970));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_21 (.CI(n39362), .I0(n10588[18]), .I1(GND_net), 
            .CO(n39363));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10588[17]), .I2(GND_net), 
            .I3(n39361), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4973));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_20 (.CI(n39361), .I0(n10588[17]), .I1(GND_net), 
            .CO(n39362));
    SB_CARRY add_5053_13 (.CI(n39211), .I0(n15969[10]), .I1(n898_adj_4969), 
            .CO(n39212));
    SB_LUT4 add_5053_12_lut (.I0(GND_net), .I1(n15969[9]), .I2(n825_adj_4975), 
            .I3(n39210), .O(n15425[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_12 (.CI(n39210), .I0(n15969[9]), .I1(n825_adj_4975), 
            .CO(n39211));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10588[16]), .I2(GND_net), 
            .I3(n39360), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_11_lut (.I0(GND_net), .I1(n15969[8]), .I2(n752_adj_4976), 
            .I3(n39209), .O(n15425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_11 (.CI(n39209), .I0(n15969[8]), .I1(n752_adj_4976), 
            .CO(n39210));
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_19 (.CI(n39360), .I0(n10588[16]), .I1(GND_net), 
            .CO(n39361));
    SB_LUT4 add_5053_10_lut (.I0(GND_net), .I1(n15969[7]), .I2(n679_adj_4977), 
            .I3(n39208), .O(n15425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10588[15]), .I2(GND_net), 
            .I3(n39359), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n39359), .I0(n10588[15]), .I1(GND_net), 
            .CO(n39360));
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4979));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5053_10 (.CI(n39208), .I0(n15969[7]), .I1(n679_adj_4977), 
            .CO(n39209));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10588[14]), .I2(GND_net), 
            .I3(n39358), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n39358), .I0(n10588[14]), .I1(GND_net), 
            .CO(n39359));
    SB_LUT4 add_958_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4236[17]), .I3(n38281), .O(\PID_CONTROLLER.integral_23__N_3672 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_19 (.CI(n38281), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4236[17]), .CO(n38282));
    SB_LUT4 add_5053_9_lut (.I0(GND_net), .I1(n15969[6]), .I2(n606_adj_4980), 
            .I3(n39207), .O(n15425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4981));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10588[13]), .I2(n1096), 
            .I3(n39357), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_9 (.CI(n39207), .I0(n15969[6]), .I1(n606_adj_4980), 
            .CO(n39208));
    SB_LUT4 add_5053_8_lut (.I0(GND_net), .I1(n15969[5]), .I2(n533_adj_4982), 
            .I3(n39206), .O(n15425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4236[16]), .I3(n38280), .O(\PID_CONTROLLER.integral_23__N_3672 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4983));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5053_8 (.CI(n39206), .I0(n15969[5]), .I1(n533_adj_4982), 
            .CO(n39207));
    SB_CARRY mult_11_add_1225_16 (.CI(n39357), .I0(n10588[13]), .I1(n1096), 
            .CO(n39358));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n11119[21]), .I2(GND_net), 
            .I3(n39599), .O(n10612[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n11119[20]), .I2(GND_net), 
            .I3(n39598), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n39598), .I0(n11119[20]), .I1(GND_net), 
            .CO(n39599));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n11119[19]), .I2(GND_net), 
            .I3(n39597), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n39597), .I0(n11119[19]), .I1(GND_net), 
            .CO(n39598));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n11119[18]), .I2(GND_net), 
            .I3(n39596), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n39596), .I0(n11119[18]), .I1(GND_net), 
            .CO(n39597));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n11119[17]), .I2(GND_net), 
            .I3(n39595), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n39595), .I0(n11119[17]), .I1(GND_net), 
            .CO(n39596));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n11119[16]), .I2(GND_net), 
            .I3(n39594), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n39594), .I0(n11119[16]), .I1(GND_net), 
            .CO(n39595));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n11119[15]), .I2(GND_net), 
            .I3(n39593), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n39593), .I0(n11119[15]), .I1(GND_net), 
            .CO(n39594));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n11119[14]), .I2(GND_net), 
            .I3(n39592), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10588[12]), .I2(n1023), 
            .I3(n39356), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_7_lut (.I0(GND_net), .I1(n15969[4]), .I2(n460_adj_4984), 
            .I3(n39205), .O(n15425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n39592), .I0(n11119[14]), .I1(GND_net), 
            .CO(n39593));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n11119[13]), .I2(n1096_adj_4985), 
            .I3(n39591), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_18 (.CI(n38280), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4236[16]), .CO(n38281));
    SB_CARRY mult_10_add_1225_16 (.CI(n39591), .I0(n11119[13]), .I1(n1096_adj_4985), 
            .CO(n39592));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n11119[12]), .I2(n1023_adj_4986), 
            .I3(n39590), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n39590), .I0(n11119[12]), .I1(n1023_adj_4986), 
            .CO(n39591));
    SB_CARRY mult_11_add_1225_15 (.CI(n39356), .I0(n10588[12]), .I1(n1023), 
            .CO(n39357));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n11119[11]), .I2(n950), 
            .I3(n39589), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_7 (.CI(n39205), .I0(n15969[4]), .I1(n460_adj_4984), 
            .CO(n39206));
    SB_CARRY mult_10_add_1225_14 (.CI(n39589), .I0(n11119[11]), .I1(n950), 
            .CO(n39590));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n11119[10]), .I2(n877), 
            .I3(n39588), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n39588), .I0(n11119[10]), .I1(n877), 
            .CO(n39589));
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5053_6_lut (.I0(GND_net), .I1(n15969[3]), .I2(n387_adj_4988), 
            .I3(n39204), .O(n15425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4989));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_958_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4236[15]), .I3(n38279), .O(\PID_CONTROLLER.integral_23__N_3672 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n11119[9]), .I2(n804), 
            .I3(n39587), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n39587), .I0(n11119[9]), .I1(n804), 
            .CO(n39588));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n11119[8]), .I2(n731), 
            .I3(n39586), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4990));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_17 (.CI(n38279), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4236[15]), .CO(n38280));
    SB_CARRY mult_10_add_1225_11 (.CI(n39586), .I0(n11119[8]), .I1(n731), 
            .CO(n39587));
    SB_LUT4 add_958_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4236[14]), .I3(n38278), .O(\PID_CONTROLLER.integral_23__N_3672 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n11119[7]), .I2(n658), 
            .I3(n39585), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n39585), .I0(n11119[7]), .I1(n658), 
            .CO(n39586));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n11119[6]), .I2(n585), 
            .I3(n39584), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10588[11]), .I2(n950_adj_4991), 
            .I3(n39355), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_6 (.CI(n39204), .I0(n15969[3]), .I1(n387_adj_4988), 
            .CO(n39205));
    SB_CARRY mult_11_add_1225_14 (.CI(n39355), .I0(n10588[11]), .I1(n950_adj_4991), 
            .CO(n39356));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10588[10]), .I2(n877_adj_4992), 
            .I3(n39354), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_5_lut (.I0(GND_net), .I1(n15969[2]), .I2(n314_adj_4993), 
            .I3(n39203), .O(n15425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n39354), .I0(n10588[10]), .I1(n877_adj_4992), 
            .CO(n39355));
    SB_CARRY mult_10_add_1225_9 (.CI(n39584), .I0(n11119[6]), .I1(n585), 
            .CO(n39585));
    SB_CARRY add_958_16 (.CI(n38278), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4236[14]), .CO(n38279));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n11119[5]), .I2(n512), 
            .I3(n39583), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5053_5 (.CI(n39203), .I0(n15969[2]), .I1(n314_adj_4993), 
            .CO(n39204));
    SB_CARRY mult_10_add_1225_8 (.CI(n39583), .I0(n11119[5]), .I1(n512), 
            .CO(n39584));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n11119[4]), .I2(n439), 
            .I3(n39582), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10588[9]), .I2(n804_adj_4994), 
            .I3(n39353), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n39582), .I0(n11119[4]), .I1(n439), 
            .CO(n39583));
    SB_LUT4 add_5053_4_lut (.I0(GND_net), .I1(n15969[1]), .I2(n241_adj_4995), 
            .I3(n39202), .O(n15425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n11119[3]), .I2(n366), 
            .I3(n39581), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n39581), .I0(n11119[3]), .I1(n366), 
            .CO(n39582));
    SB_CARRY add_5053_4 (.CI(n39202), .I0(n15969[1]), .I1(n241_adj_4995), 
            .CO(n39203));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n11119[2]), .I2(n293), 
            .I3(n39580), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n39580), .I0(n11119[2]), .I1(n293), 
            .CO(n39581));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n11119[1]), .I2(n220), 
            .I3(n39579), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n39579), .I0(n11119[1]), .I1(n220), 
            .CO(n39580));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n11119[0]), .I2(n147_adj_4996), 
            .I3(n39578), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n39578), .I0(n11119[0]), .I1(n147_adj_4996), 
            .CO(n39579));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4997), .I2(n74), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4236[13]), .I3(n38277), .O(\PID_CONTROLLER.integral_23__N_3672 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4997), .I1(n74), 
            .CO(n39578));
    SB_LUT4 add_4846_23_lut (.I0(GND_net), .I1(n12088[20]), .I2(GND_net), 
            .I3(n39577), .O(n11119[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_15 (.CI(n38277), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4236[13]), .CO(n38278));
    SB_LUT4 add_4846_22_lut (.I0(GND_net), .I1(n12088[19]), .I2(GND_net), 
            .I3(n39576), .O(n11119[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_22 (.CI(n39576), .I0(n12088[19]), .I1(GND_net), 
            .CO(n39577));
    SB_LUT4 add_4846_21_lut (.I0(GND_net), .I1(n12088[18]), .I2(GND_net), 
            .I3(n39575), .O(n11119[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4236[12]), .I3(n38276), .O(\PID_CONTROLLER.integral_23__N_3672 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_21 (.CI(n39575), .I0(n12088[18]), .I1(GND_net), 
            .CO(n39576));
    SB_LUT4 add_4846_20_lut (.I0(GND_net), .I1(n12088[17]), .I2(GND_net), 
            .I3(n39574), .O(n11119[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_20 (.CI(n39574), .I0(n12088[17]), .I1(GND_net), 
            .CO(n39575));
    SB_CARRY add_958_14 (.CI(n38276), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4236[12]), .CO(n38277));
    SB_CARRY mult_11_add_1225_12 (.CI(n39353), .I0(n10588[9]), .I1(n804_adj_4994), 
            .CO(n39354));
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4998));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_958_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4236[11]), .I3(n38275), .O(\PID_CONTROLLER.integral_23__N_3672 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4846_19_lut (.I0(GND_net), .I1(n12088[16]), .I2(GND_net), 
            .I3(n39573), .O(n11119[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_19 (.CI(n39573), .I0(n12088[16]), .I1(GND_net), 
            .CO(n39574));
    SB_LUT4 add_4846_18_lut (.I0(GND_net), .I1(n12088[15]), .I2(GND_net), 
            .I3(n39572), .O(n11119[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_13 (.CI(n38275), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4236[11]), .CO(n38276));
    SB_CARRY add_4846_18 (.CI(n39572), .I0(n12088[15]), .I1(GND_net), 
            .CO(n39573));
    SB_LUT4 add_4846_17_lut (.I0(GND_net), .I1(n12088[14]), .I2(GND_net), 
            .I3(n39571), .O(n11119[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_17 (.CI(n39571), .I0(n12088[14]), .I1(GND_net), 
            .CO(n39572));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10588[8]), .I2(n731_adj_4999), 
            .I3(n39352), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_3_lut (.I0(GND_net), .I1(n15969[0]), .I2(n168_adj_5000), 
            .I3(n39201), .O(n15425[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_5001));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5053_3 (.CI(n39201), .I0(n15969[0]), .I1(n168_adj_5000), 
            .CO(n39202));
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_5002));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4846_16_lut (.I0(GND_net), .I1(n12088[13]), .I2(n1099), 
            .I3(n39570), .O(n11119[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_16 (.CI(n39570), .I0(n12088[13]), .I1(n1099), .CO(n39571));
    SB_LUT4 add_4846_15_lut (.I0(GND_net), .I1(n12088[12]), .I2(n1026), 
            .I3(n39569), .O(n11119[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4846_15 (.CI(n39569), .I0(n12088[12]), .I1(n1026), .CO(n39570));
    SB_LUT4 add_4846_14_lut (.I0(GND_net), .I1(n12088[11]), .I2(n953), 
            .I3(n39568), .O(n11119[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n39352), .I0(n10588[8]), .I1(n731_adj_4999), 
            .CO(n39353));
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4894));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10588[7]), .I2(n658_adj_5003), 
            .I3(n39351), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5053_2_lut (.I0(GND_net), .I1(n26_adj_5004), .I2(n95_adj_5005), 
            .I3(GND_net), .O(n15425[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5053_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n39351), .I0(n10588[7]), .I1(n658_adj_5003), 
            .CO(n39352));
    SB_CARRY add_4846_14 (.CI(n39568), .I0(n12088[11]), .I1(n953), .CO(n39569));
    SB_LUT4 add_4846_13_lut (.I0(GND_net), .I1(n12088[10]), .I2(n880), 
            .I3(n39567), .O(n11119[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4236[10]), .I3(n38274), .O(\PID_CONTROLLER.integral_23__N_3672 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_13 (.CI(n39567), .I0(n12088[10]), .I1(n880), .CO(n39568));
    SB_LUT4 add_4846_12_lut (.I0(GND_net), .I1(n12088[9]), .I2(n807), 
            .I3(n39566), .O(n11119[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_12 (.CI(n39566), .I0(n12088[9]), .I1(n807), .CO(n39567));
    SB_LUT4 add_4846_11_lut (.I0(GND_net), .I1(n12088[8]), .I2(n734), 
            .I3(n39565), .O(n11119[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_11 (.CI(n39565), .I0(n12088[8]), .I1(n734), .CO(n39566));
    SB_CARRY add_5053_2 (.CI(GND_net), .I0(n26_adj_5004), .I1(n95_adj_5005), 
            .CO(n39201));
    SB_LUT4 add_4846_10_lut (.I0(GND_net), .I1(n12088[7]), .I2(n661_adj_5006), 
            .I3(n39564), .O(n11119[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_10 (.CI(n39564), .I0(n12088[7]), .I1(n661_adj_5006), 
            .CO(n39565));
    SB_LUT4 add_4846_9_lut (.I0(GND_net), .I1(n12088[6]), .I2(n588_adj_5007), 
            .I3(n39563), .O(n11119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10588[6]), .I2(n585_adj_5008), 
            .I3(n39350), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_9 (.CI(n39563), .I0(n12088[6]), .I1(n588_adj_5007), 
            .CO(n39564));
    SB_LUT4 add_5253_9_lut (.I0(GND_net), .I1(n18416[6]), .I2(n630_adj_5009), 
            .I3(n39200), .O(n18289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4846_8_lut (.I0(GND_net), .I1(n12088[5]), .I2(n515_adj_5010), 
            .I3(n39562), .O(n11119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n39350), .I0(n10588[6]), .I1(n585_adj_5008), 
            .CO(n39351));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10588[5]), .I2(n512_adj_5011), 
            .I3(n39349), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_8_lut (.I0(GND_net), .I1(n18416[5]), .I2(n557_adj_5012), 
            .I3(n39199), .O(n18289[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_8 (.CI(n39199), .I0(n18416[5]), .I1(n557_adj_5012), 
            .CO(n39200));
    SB_CARRY add_4846_8 (.CI(n39562), .I0(n12088[5]), .I1(n515_adj_5010), 
            .CO(n39563));
    SB_LUT4 add_4846_7_lut (.I0(GND_net), .I1(n12088[4]), .I2(n442_adj_5013), 
            .I3(n39561), .O(n11119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_7 (.CI(n39561), .I0(n12088[4]), .I1(n442_adj_5013), 
            .CO(n39562));
    SB_LUT4 add_4846_6_lut (.I0(GND_net), .I1(n12088[3]), .I2(n369_adj_5014), 
            .I3(n39560), .O(n11119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[23]), 
            .I3(n38402), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_6 (.CI(n39560), .I0(n12088[3]), .I1(n369_adj_5014), 
            .CO(n39561));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[22]), 
            .I3(n38401), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4846_5_lut (.I0(GND_net), .I1(n12088[2]), .I2(n296_adj_5017), 
            .I3(n39559), .O(n11119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_5 (.CI(n39559), .I0(n12088[2]), .I1(n296_adj_5017), 
            .CO(n39560));
    SB_LUT4 add_4846_4_lut (.I0(GND_net), .I1(n12088[1]), .I2(n223_adj_5018), 
            .I3(n39558), .O(n11119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n38401), .I0(GND_net), .I1(n1_adj_5147[22]), 
            .CO(n38402));
    SB_CARRY add_4846_4 (.CI(n39558), .I0(n12088[1]), .I1(n223_adj_5018), 
            .CO(n39559));
    SB_LUT4 add_4846_3_lut (.I0(GND_net), .I1(n12088[0]), .I2(n150_adj_5019), 
            .I3(n39557), .O(n11119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_3 (.CI(n39557), .I0(n12088[0]), .I1(n150_adj_5019), 
            .CO(n39558));
    SB_LUT4 add_4846_2_lut (.I0(GND_net), .I1(n8_adj_5020), .I2(n77_adj_5021), 
            .I3(GND_net), .O(n11119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_12 (.CI(n38274), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4236[10]), .CO(n38275));
    SB_CARRY add_4846_2 (.CI(GND_net), .I0(n8_adj_5020), .I1(n77_adj_5021), 
            .CO(n39557));
    SB_LUT4 add_4889_22_lut (.I0(GND_net), .I1(n12969[19]), .I2(GND_net), 
            .I3(n39556), .O(n12088[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_7_lut (.I0(GND_net), .I1(n18416[4]), .I2(n484_adj_5022), 
            .I3(n39198), .O(n18289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_21_lut (.I0(GND_net), .I1(n12969[18]), .I2(GND_net), 
            .I3(n39555), .O(n12088[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_21 (.CI(n39555), .I0(n12969[18]), .I1(GND_net), 
            .CO(n39556));
    SB_LUT4 add_4889_20_lut (.I0(GND_net), .I1(n12969[17]), .I2(GND_net), 
            .I3(n39554), .O(n12088[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_20 (.CI(n39554), .I0(n12969[17]), .I1(GND_net), 
            .CO(n39555));
    SB_LUT4 add_4889_19_lut (.I0(GND_net), .I1(n12969[16]), .I2(GND_net), 
            .I3(n39553), .O(n12088[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_19 (.CI(n39553), .I0(n12969[16]), .I1(GND_net), 
            .CO(n39554));
    SB_CARRY mult_11_add_1225_8 (.CI(n39349), .I0(n10588[5]), .I1(n512_adj_5011), 
            .CO(n39350));
    SB_LUT4 add_4889_18_lut (.I0(GND_net), .I1(n12969[15]), .I2(GND_net), 
            .I3(n39552), .O(n12088[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_7 (.CI(n39198), .I0(n18416[4]), .I1(n484_adj_5022), 
            .CO(n39199));
    SB_CARRY add_4889_18 (.CI(n39552), .I0(n12969[15]), .I1(GND_net), 
            .CO(n39553));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[21]), 
            .I3(n38400), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_17_lut (.I0(GND_net), .I1(n12969[14]), .I2(GND_net), 
            .I3(n39551), .O(n12088[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_17 (.CI(n39551), .I0(n12969[14]), .I1(GND_net), 
            .CO(n39552));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10588[4]), .I2(n439_adj_5024), 
            .I3(n39348), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5253_6_lut (.I0(GND_net), .I1(n18416[3]), .I2(n411_adj_5025), 
            .I3(n39197), .O(n18289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4236[9]), .I3(n38273), .O(\PID_CONTROLLER.integral_23__N_3672 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n38400), .I0(GND_net), .I1(n1_adj_5147[21]), 
            .CO(n38401));
    SB_CARRY mult_11_add_1225_7 (.CI(n39348), .I0(n10588[4]), .I1(n439_adj_5024), 
            .CO(n39349));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10588[3]), .I2(n366_adj_5026), 
            .I3(n39347), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n39347), .I0(n10588[3]), .I1(n366_adj_5026), 
            .CO(n39348));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10588[2]), .I2(n293_adj_5027), 
            .I3(n39346), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n39346), .I0(n10588[2]), .I1(n293_adj_5027), 
            .CO(n39347));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10588[1]), .I2(n220_adj_5028), 
            .I3(n39345), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[20]), 
            .I3(n38399), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_6 (.CI(n39197), .I0(n18416[3]), .I1(n411_adj_5025), 
            .CO(n39198));
    SB_CARRY mult_11_add_1225_4 (.CI(n39345), .I0(n10588[1]), .I1(n220_adj_5028), 
            .CO(n39346));
    SB_LUT4 add_5253_5_lut (.I0(GND_net), .I1(n18416[2]), .I2(n338_adj_5030), 
            .I3(n39196), .O(n18289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10588[0]), .I2(n147_adj_5031), 
            .I3(n39344), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_5 (.CI(n39196), .I0(n18416[2]), .I1(n338_adj_5030), 
            .CO(n39197));
    SB_LUT4 add_4889_16_lut (.I0(GND_net), .I1(n12969[13]), .I2(n1102_adj_5032), 
            .I3(n39550), .O(n12088[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_16 (.CI(n39550), .I0(n12969[13]), .I1(n1102_adj_5032), 
            .CO(n39551));
    SB_CARRY add_958_11 (.CI(n38273), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4236[9]), .CO(n38274));
    SB_LUT4 add_4889_15_lut (.I0(GND_net), .I1(n12969[12]), .I2(n1029_adj_5033), 
            .I3(n39549), .O(n12088[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_15 (.CI(n39549), .I0(n12969[12]), .I1(n1029_adj_5033), 
            .CO(n39550));
    SB_LUT4 add_4889_14_lut (.I0(GND_net), .I1(n12969[11]), .I2(n956_adj_5034), 
            .I3(n39548), .O(n12088[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n39344), .I0(n10588[0]), .I1(n147_adj_5031), 
            .CO(n39345));
    SB_CARRY add_4889_14 (.CI(n39548), .I0(n12969[11]), .I1(n956_adj_5034), 
            .CO(n39549));
    SB_LUT4 add_5253_4_lut (.I0(GND_net), .I1(n18416[1]), .I2(n265_adj_5035), 
            .I3(n39195), .O(n18289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_13_lut (.I0(GND_net), .I1(n12969[10]), .I2(n883_adj_5036), 
            .I3(n39547), .O(n12088[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4236[8]), .I3(n38272), .O(\PID_CONTROLLER.integral_23__N_3672 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_13 (.CI(n39547), .I0(n12969[10]), .I1(n883_adj_5036), 
            .CO(n39548));
    SB_LUT4 add_4889_12_lut (.I0(GND_net), .I1(n12969[9]), .I2(n810_adj_5037), 
            .I3(n39546), .O(n12088[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n38399), .I0(GND_net), .I1(n1_adj_5147[20]), 
            .CO(n38400));
    SB_CARRY add_4889_12 (.CI(n39546), .I0(n12969[9]), .I1(n810_adj_5037), 
            .CO(n39547));
    SB_LUT4 add_4889_11_lut (.I0(GND_net), .I1(n12969[8]), .I2(n737_adj_5038), 
            .I3(n39545), .O(n12088[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_4 (.CI(n39195), .I0(n18416[1]), .I1(n265_adj_5035), 
            .CO(n39196));
    SB_CARRY add_4889_11 (.CI(n39545), .I0(n12969[8]), .I1(n737_adj_5038), 
            .CO(n39546));
    SB_CARRY add_958_10 (.CI(n38272), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4236[8]), .CO(n38273));
    SB_LUT4 add_4889_10_lut (.I0(GND_net), .I1(n12969[7]), .I2(n664_adj_5039), 
            .I3(n39544), .O(n12088[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_10 (.CI(n39544), .I0(n12969[7]), .I1(n664_adj_5039), 
            .CO(n39545));
    SB_LUT4 add_4889_9_lut (.I0(GND_net), .I1(n12969[6]), .I2(n591_adj_5040), 
            .I3(n39543), .O(n12088[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[19]), 
            .I3(n38398), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_9 (.CI(n39543), .I0(n12969[6]), .I1(n591_adj_5040), 
            .CO(n39544));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n38398), .I0(GND_net), .I1(n1_adj_5147[19]), 
            .CO(n38399));
    SB_LUT4 add_4889_8_lut (.I0(GND_net), .I1(n12969[5]), .I2(n518_adj_5042), 
            .I3(n39542), .O(n12088[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_8 (.CI(n39542), .I0(n12969[5]), .I1(n518_adj_5042), 
            .CO(n39543));
    SB_LUT4 add_5253_3_lut (.I0(GND_net), .I1(n18416[0]), .I2(n192_adj_5043), 
            .I3(n39194), .O(n18289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[18]), 
            .I3(n38397), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5253_3 (.CI(n39194), .I0(n18416[0]), .I1(n192_adj_5043), 
            .CO(n39195));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_5045), .I2(n74_adj_5046), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_7_lut (.I0(GND_net), .I1(n12969[4]), .I2(n445_adj_5047), 
            .I3(n39541), .O(n12088[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_7 (.CI(n39541), .I0(n12969[4]), .I1(n445_adj_5047), 
            .CO(n39542));
    SB_LUT4 add_5253_2_lut (.I0(GND_net), .I1(n50_adj_5048), .I2(n119_adj_5049), 
            .I3(GND_net), .O(n18289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5253_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_5045), .I1(n74_adj_5046), 
            .CO(n39344));
    SB_LUT4 add_4823_23_lut (.I0(GND_net), .I1(n11605[20]), .I2(GND_net), 
            .I3(n39343), .O(n10588[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_22_lut (.I0(GND_net), .I1(n11605[19]), .I2(GND_net), 
            .I3(n39342), .O(n10588[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_22 (.CI(n39342), .I0(n11605[19]), .I1(GND_net), 
            .CO(n39343));
    SB_CARRY add_5253_2 (.CI(GND_net), .I0(n50_adj_5048), .I1(n119_adj_5049), 
            .CO(n39194));
    SB_LUT4 add_958_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4236[7]), .I3(n38271), .O(\PID_CONTROLLER.integral_23__N_3672 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_16_lut (.I0(GND_net), .I1(n16449[13]), .I2(n1120_adj_5050), 
            .I3(n39193), .O(n15969[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n38397), .I0(GND_net), .I1(n1_adj_5147[18]), 
            .CO(n38398));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[17]), 
            .I3(n38396), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_21_lut (.I0(GND_net), .I1(n11605[18]), .I2(GND_net), 
            .I3(n39341), .O(n10588[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n38396), .I0(GND_net), .I1(n1_adj_5147[17]), 
            .CO(n38397));
    SB_LUT4 add_5084_15_lut (.I0(GND_net), .I1(n16449[12]), .I2(n1047_adj_5052), 
            .I3(n39192), .O(n15969[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[16]), 
            .I3(n38395), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_9 (.CI(n38271), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4236[7]), .CO(n38272));
    SB_CARRY add_4823_21 (.CI(n39341), .I0(n11605[18]), .I1(GND_net), 
            .CO(n39342));
    SB_CARRY unary_minus_16_add_3_18 (.CI(n38395), .I0(GND_net), .I1(n1_adj_5147[16]), 
            .CO(n38396));
    SB_CARRY add_5084_15 (.CI(n39192), .I0(n16449[12]), .I1(n1047_adj_5052), 
            .CO(n39193));
    SB_LUT4 add_958_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4236[6]), .I3(n38270), .O(\PID_CONTROLLER.integral_23__N_3672 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_20_lut (.I0(GND_net), .I1(n11605[17]), .I2(GND_net), 
            .I3(n39340), .O(n10588[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_6_lut (.I0(GND_net), .I1(n12969[3]), .I2(n372_adj_5054), 
            .I3(n39540), .O(n12088[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_14_lut (.I0(GND_net), .I1(n16449[11]), .I2(n974_adj_5055), 
            .I3(n39191), .O(n15969[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_20 (.CI(n39340), .I0(n11605[17]), .I1(GND_net), 
            .CO(n39341));
    SB_CARRY add_5084_14 (.CI(n39191), .I0(n16449[11]), .I1(n974_adj_5055), 
            .CO(n39192));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[15]), 
            .I3(n38394), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n38394), .I0(GND_net), .I1(n1_adj_5147[15]), 
            .CO(n38395));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[14]), 
            .I3(n38393), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_6 (.CI(n39540), .I0(n12969[3]), .I1(n372_adj_5054), 
            .CO(n39541));
    SB_LUT4 add_4889_5_lut (.I0(GND_net), .I1(n12969[2]), .I2(n299_adj_5058), 
            .I3(n39539), .O(n12088[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n38393), .I0(GND_net), .I1(n1_adj_5147[14]), 
            .CO(n38394));
    SB_CARRY add_4889_5 (.CI(n39539), .I0(n12969[2]), .I1(n299_adj_5058), 
            .CO(n39540));
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_5059));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4893));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[13]), 
            .I3(n38392), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_19_lut (.I0(GND_net), .I1(n11605[16]), .I2(GND_net), 
            .I3(n39339), .O(n10588[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_19 (.CI(n39339), .I0(n11605[16]), .I1(GND_net), 
            .CO(n39340));
    SB_LUT4 add_4823_18_lut (.I0(GND_net), .I1(n11605[15]), .I2(GND_net), 
            .I3(n39338), .O(n10588[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_18 (.CI(n39338), .I0(n11605[15]), .I1(GND_net), 
            .CO(n39339));
    SB_LUT4 add_5084_13_lut (.I0(GND_net), .I1(n16449[10]), .I2(n901_adj_5061), 
            .I3(n39190), .O(n15969[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_13 (.CI(n39190), .I0(n16449[10]), .I1(n901_adj_5061), 
            .CO(n39191));
    SB_LUT4 add_4823_17_lut (.I0(GND_net), .I1(n11605[14]), .I2(GND_net), 
            .I3(n39337), .O(n10588[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n38392), .I0(GND_net), .I1(n1_adj_5147[13]), 
            .CO(n38393));
    SB_CARRY add_958_8 (.CI(n38270), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4236[6]), .CO(n38271));
    SB_LUT4 add_5084_12_lut (.I0(GND_net), .I1(n16449[9]), .I2(n828_adj_5062), 
            .I3(n39189), .O(n15969[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_17 (.CI(n39337), .I0(n11605[14]), .I1(GND_net), 
            .CO(n39338));
    SB_LUT4 add_4823_16_lut (.I0(GND_net), .I1(n11605[13]), .I2(n1099_adj_5063), 
            .I3(n39336), .O(n10588[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_12 (.CI(n39189), .I0(n16449[9]), .I1(n828_adj_5062), 
            .CO(n39190));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[12]), 
            .I3(n38391), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n38391), .I0(GND_net), .I1(n1_adj_5147[12]), 
            .CO(n38392));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[11]), 
            .I3(n38390), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n38390), .I0(GND_net), .I1(n1_adj_5147[11]), 
            .CO(n38391));
    SB_LUT4 add_5084_11_lut (.I0(GND_net), .I1(n16449[8]), .I2(n755_adj_5066), 
            .I3(n39188), .O(n15969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[10]), 
            .I3(n38389), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4236[5]), .I3(n38269), .O(\PID_CONTROLLER.integral_23__N_3672 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_11 (.CI(n39188), .I0(n16449[8]), .I1(n755_adj_5066), 
            .CO(n39189));
    SB_LUT4 add_5084_10_lut (.I0(GND_net), .I1(n16449[7]), .I2(n682_adj_5068), 
            .I3(n39187), .O(n15969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_16 (.CI(n39336), .I0(n11605[13]), .I1(n1099_adj_5063), 
            .CO(n39337));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n38389), .I0(GND_net), .I1(n1_adj_5147[10]), 
            .CO(n38390));
    SB_CARRY add_958_7 (.CI(n38269), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4236[5]), .CO(n38270));
    SB_LUT4 add_958_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4236[4]), .I3(n38268), .O(\PID_CONTROLLER.integral_23__N_3672 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_10 (.CI(n39187), .I0(n16449[7]), .I1(n682_adj_5068), 
            .CO(n39188));
    SB_LUT4 add_4823_15_lut (.I0(GND_net), .I1(n11605[12]), .I2(n1026_adj_5069), 
            .I3(n39335), .O(n10588[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_9_lut (.I0(GND_net), .I1(n16449[6]), .I2(n609_adj_5070), 
            .I3(n39186), .O(n15969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_9 (.CI(n39186), .I0(n16449[6]), .I1(n609_adj_5070), 
            .CO(n39187));
    SB_CARRY add_958_6 (.CI(n38268), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4236[4]), .CO(n38269));
    SB_CARRY add_4823_15 (.CI(n39335), .I0(n11605[12]), .I1(n1026_adj_5069), 
            .CO(n39336));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[9]), 
            .I3(n38388), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_4_lut (.I0(GND_net), .I1(n12969[1]), .I2(n226_adj_5072), 
            .I3(n39538), .O(n12088[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4236[3]), .I3(n38267), .O(\PID_CONTROLLER.integral_23__N_3672 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_4 (.CI(n39538), .I0(n12969[1]), .I1(n226_adj_5072), 
            .CO(n39539));
    SB_LUT4 add_4823_14_lut (.I0(GND_net), .I1(n11605[11]), .I2(n953_adj_5073), 
            .I3(n39334), .O(n10588[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_3_lut (.I0(GND_net), .I1(n12969[0]), .I2(n153_adj_5074), 
            .I3(n39537), .O(n12088[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_8_lut (.I0(GND_net), .I1(n16449[5]), .I2(n536_adj_5075), 
            .I3(n39185), .O(n15969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_8 (.CI(n39185), .I0(n16449[5]), .I1(n536_adj_5075), 
            .CO(n39186));
    SB_CARRY add_958_5 (.CI(n38267), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4236[3]), .CO(n38268));
    SB_CARRY add_4889_3 (.CI(n39537), .I0(n12969[0]), .I1(n153_adj_5074), 
            .CO(n39538));
    SB_LUT4 add_4889_2_lut (.I0(GND_net), .I1(n11_adj_5076), .I2(n80_adj_5077), 
            .I3(GND_net), .O(n12088[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_2 (.CI(GND_net), .I0(n11_adj_5076), .I1(n80_adj_5077), 
            .CO(n39537));
    SB_LUT4 add_4929_21_lut (.I0(GND_net), .I1(n13768[18]), .I2(GND_net), 
            .I3(n39536), .O(n12969[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_20_lut (.I0(GND_net), .I1(n13768[17]), .I2(GND_net), 
            .I3(n39535), .O(n12969[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n38388), .I0(GND_net), .I1(n1_adj_5147[9]), 
            .CO(n38389));
    SB_CARRY add_4823_14 (.CI(n39334), .I0(n11605[11]), .I1(n953_adj_5073), 
            .CO(n39335));
    SB_LUT4 add_958_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4236[2]), .I3(n38266), .O(\PID_CONTROLLER.integral_23__N_3672 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_20 (.CI(n39535), .I0(n13768[17]), .I1(GND_net), 
            .CO(n39536));
    SB_LUT4 add_4823_13_lut (.I0(GND_net), .I1(n11605[10]), .I2(n880_adj_5078), 
            .I3(n39333), .O(n10588[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_19_lut (.I0(GND_net), .I1(n13768[16]), .I2(GND_net), 
            .I3(n39534), .O(n12969[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_4 (.CI(n38266), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4236[2]), .CO(n38267));
    SB_CARRY add_4929_19 (.CI(n39534), .I0(n13768[16]), .I1(GND_net), 
            .CO(n39535));
    SB_LUT4 add_4929_18_lut (.I0(GND_net), .I1(n13768[15]), .I2(GND_net), 
            .I3(n39533), .O(n12969[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_13 (.CI(n39333), .I0(n11605[10]), .I1(n880_adj_5078), 
            .CO(n39334));
    SB_LUT4 add_4823_12_lut (.I0(GND_net), .I1(n11605[9]), .I2(n807_adj_5079), 
            .I3(n39332), .O(n10588[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_12 (.CI(n39332), .I0(n11605[9]), .I1(n807_adj_5079), 
            .CO(n39333));
    SB_LUT4 add_4823_11_lut (.I0(GND_net), .I1(n11605[8]), .I2(n734_adj_5080), 
            .I3(n39331), .O(n10588[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_18 (.CI(n39533), .I0(n13768[15]), .I1(GND_net), 
            .CO(n39534));
    SB_LUT4 add_5084_7_lut (.I0(GND_net), .I1(n16449[4]), .I2(n463_adj_5081), 
            .I3(n39184), .O(n15969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_17_lut (.I0(GND_net), .I1(n13768[14]), .I2(GND_net), 
            .I3(n39532), .O(n12969[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_17 (.CI(n39532), .I0(n13768[14]), .I1(GND_net), 
            .CO(n39533));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5084_7 (.CI(n39184), .I0(n16449[4]), .I1(n463_adj_5081), 
            .CO(n39185));
    SB_LUT4 add_4929_16_lut (.I0(GND_net), .I1(n13768[13]), .I2(n1105_adj_5083), 
            .I3(n39531), .O(n12969[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_16 (.CI(n39531), .I0(n13768[13]), .I1(n1105_adj_5083), 
            .CO(n39532));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[8]), 
            .I3(n38387), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_15_lut (.I0(GND_net), .I1(n13768[12]), .I2(n1032_adj_5059), 
            .I3(n39530), .O(n12969[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_15 (.CI(n39530), .I0(n13768[12]), .I1(n1032_adj_5059), 
            .CO(n39531));
    SB_CARRY add_4823_11 (.CI(n39331), .I0(n11605[8]), .I1(n734_adj_5080), 
            .CO(n39332));
    SB_LUT4 add_4929_14_lut (.I0(GND_net), .I1(n13768[11]), .I2(n959_adj_5002), 
            .I3(n39529), .O(n12969[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_14 (.CI(n39529), .I0(n13768[11]), .I1(n959_adj_5002), 
            .CO(n39530));
    SB_LUT4 add_4929_13_lut (.I0(GND_net), .I1(n13768[10]), .I2(n886_adj_5001), 
            .I3(n39528), .O(n12969[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_13 (.CI(n39528), .I0(n13768[10]), .I1(n886_adj_5001), 
            .CO(n39529));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n38387), .I0(GND_net), .I1(n1_adj_5147[8]), 
            .CO(n38388));
    SB_LUT4 add_4929_12_lut (.I0(GND_net), .I1(n13768[9]), .I2(n813_adj_4998), 
            .I3(n39527), .O(n12969[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_12 (.CI(n39527), .I0(n13768[9]), .I1(n813_adj_4998), 
            .CO(n39528));
    SB_LUT4 add_4929_11_lut (.I0(GND_net), .I1(n13768[8]), .I2(n740_adj_4990), 
            .I3(n39526), .O(n12969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_11 (.CI(n39526), .I0(n13768[8]), .I1(n740_adj_4990), 
            .CO(n39527));
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_5083));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4929_10_lut (.I0(GND_net), .I1(n13768[7]), .I2(n667_adj_4989), 
            .I3(n39525), .O(n12969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_5081));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4929_10 (.CI(n39525), .I0(n13768[7]), .I1(n667_adj_4989), 
            .CO(n39526));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[7]), 
            .I3(n38386), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_9_lut (.I0(GND_net), .I1(n13768[6]), .I2(n594_adj_4983), 
            .I3(n39524), .O(n12969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_9 (.CI(n39524), .I0(n13768[6]), .I1(n594_adj_4983), 
            .CO(n39525));
    SB_LUT4 add_4823_10_lut (.I0(GND_net), .I1(n11605[7]), .I2(n661), 
            .I3(n39330), .O(n10588[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_8_lut (.I0(GND_net), .I1(n13768[5]), .I2(n521_adj_4981), 
            .I3(n39523), .O(n12969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n38386), .I0(GND_net), .I1(n1_adj_5147[7]), 
            .CO(n38387));
    SB_CARRY add_4823_10 (.CI(n39330), .I0(n11605[7]), .I1(n661), .CO(n39331));
    SB_CARRY add_4929_8 (.CI(n39523), .I0(n13768[5]), .I1(n521_adj_4981), 
            .CO(n39524));
    SB_LUT4 add_4929_7_lut (.I0(GND_net), .I1(n13768[4]), .I2(n448_adj_4979), 
            .I3(n39522), .O(n12969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_9_lut (.I0(GND_net), .I1(n11605[6]), .I2(n588), .I3(n39329), 
            .O(n10588[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_9 (.CI(n39329), .I0(n11605[6]), .I1(n588), .CO(n39330));
    SB_CARRY add_4929_7 (.CI(n39522), .I0(n13768[4]), .I1(n448_adj_4979), 
            .CO(n39523));
    SB_LUT4 add_5084_6_lut (.I0(GND_net), .I1(n16449[3]), .I2(n390_adj_4974), 
            .I3(n39183), .O(n15969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_6_lut (.I0(GND_net), .I1(n13768[3]), .I2(n375_adj_4973), 
            .I3(n39521), .O(n12969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_6 (.CI(n39521), .I0(n13768[3]), .I1(n375_adj_4973), 
            .CO(n39522));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[6]), 
            .I3(n38385), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4929_5_lut (.I0(GND_net), .I1(n13768[2]), .I2(n302_adj_4971), 
            .I3(n39520), .O(n12969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_5 (.CI(n39520), .I0(n13768[2]), .I1(n302_adj_4971), 
            .CO(n39521));
    SB_LUT4 add_4929_4_lut (.I0(GND_net), .I1(n13768[1]), .I2(n229_adj_4970), 
            .I3(n39519), .O(n12969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_6 (.CI(n39183), .I0(n16449[3]), .I1(n390_adj_4974), 
            .CO(n39184));
    SB_LUT4 add_4823_8_lut (.I0(GND_net), .I1(n11605[5]), .I2(n515), .I3(n39328), 
            .O(n10588[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4236[1]), .I3(n38265), .O(\PID_CONTROLLER.integral_23__N_3672 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_8 (.CI(n39328), .I0(n11605[5]), .I1(n515), .CO(n39329));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n38385), .I0(GND_net), .I1(n1_adj_5147[6]), 
            .CO(n38386));
    SB_CARRY add_4929_4 (.CI(n39519), .I0(n13768[1]), .I1(n229_adj_4970), 
            .CO(n39520));
    SB_LUT4 add_4929_3_lut (.I0(GND_net), .I1(n13768[0]), .I2(n156_adj_4967), 
            .I3(n39518), .O(n12969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_3 (.CI(n39518), .I0(n13768[0]), .I1(n156_adj_4967), 
            .CO(n39519));
    SB_LUT4 add_4929_2_lut (.I0(GND_net), .I1(n14_adj_4966), .I2(n83_adj_4965), 
            .I3(GND_net), .O(n12969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4929_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4929_2 (.CI(GND_net), .I0(n14_adj_4966), .I1(n83_adj_4965), 
            .CO(n39518));
    SB_LUT4 add_4967_20_lut (.I0(GND_net), .I1(n14489[17]), .I2(GND_net), 
            .I3(n39517), .O(n13768[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4967_19_lut (.I0(GND_net), .I1(n14489[16]), .I2(GND_net), 
            .I3(n39516), .O(n13768[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_19 (.CI(n39516), .I0(n14489[16]), .I1(GND_net), 
            .CO(n39517));
    SB_LUT4 add_4967_18_lut (.I0(GND_net), .I1(n14489[15]), .I2(GND_net), 
            .I3(n39515), .O(n13768[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_18 (.CI(n39515), .I0(n14489[15]), .I1(GND_net), 
            .CO(n39516));
    SB_LUT4 add_4967_17_lut (.I0(GND_net), .I1(n14489[14]), .I2(GND_net), 
            .I3(n39514), .O(n13768[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_17 (.CI(n39514), .I0(n14489[14]), .I1(GND_net), 
            .CO(n39515));
    SB_LUT4 add_4967_16_lut (.I0(GND_net), .I1(n14489[13]), .I2(n1108_adj_4963), 
            .I3(n39513), .O(n13768[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_16 (.CI(n39513), .I0(n14489[13]), .I1(n1108_adj_4963), 
            .CO(n39514));
    SB_LUT4 add_4967_15_lut (.I0(GND_net), .I1(n14489[12]), .I2(n1035_adj_4962), 
            .I3(n39512), .O(n13768[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_15 (.CI(n39512), .I0(n14489[12]), .I1(n1035_adj_4962), 
            .CO(n39513));
    SB_LUT4 add_4967_14_lut (.I0(GND_net), .I1(n14489[11]), .I2(n962_adj_4961), 
            .I3(n39511), .O(n13768[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_14 (.CI(n39511), .I0(n14489[11]), .I1(n962_adj_4961), 
            .CO(n39512));
    SB_LUT4 add_4967_13_lut (.I0(GND_net), .I1(n14489[10]), .I2(n889_adj_4956), 
            .I3(n39510), .O(n13768[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_13 (.CI(n39510), .I0(n14489[10]), .I1(n889_adj_4956), 
            .CO(n39511));
    SB_LUT4 add_4967_12_lut (.I0(GND_net), .I1(n14489[9]), .I2(n816_adj_4955), 
            .I3(n39509), .O(n13768[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_12 (.CI(n39509), .I0(n14489[9]), .I1(n816_adj_4955), 
            .CO(n39510));
    SB_LUT4 add_4967_11_lut (.I0(GND_net), .I1(n14489[8]), .I2(n743_adj_4954), 
            .I3(n39508), .O(n13768[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_11 (.CI(n39508), .I0(n14489[8]), .I1(n743_adj_4954), 
            .CO(n39509));
    SB_LUT4 add_4967_10_lut (.I0(GND_net), .I1(n14489[7]), .I2(n670_adj_4953), 
            .I3(n39507), .O(n13768[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_10 (.CI(n39507), .I0(n14489[7]), .I1(n670_adj_4953), 
            .CO(n39508));
    SB_LUT4 add_4967_9_lut (.I0(GND_net), .I1(n14489[6]), .I2(n597_adj_4952), 
            .I3(n39506), .O(n13768[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_9 (.CI(n39506), .I0(n14489[6]), .I1(n597_adj_4952), 
            .CO(n39507));
    SB_LUT4 add_4967_8_lut (.I0(GND_net), .I1(n14489[5]), .I2(n524_adj_4951), 
            .I3(n39505), .O(n13768[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_8 (.CI(n39505), .I0(n14489[5]), .I1(n524_adj_4951), 
            .CO(n39506));
    SB_LUT4 add_4967_7_lut (.I0(GND_net), .I1(n14489[4]), .I2(n451_adj_4950), 
            .I3(n39504), .O(n13768[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_7 (.CI(n39504), .I0(n14489[4]), .I1(n451_adj_4950), 
            .CO(n39505));
    SB_LUT4 add_4967_6_lut (.I0(GND_net), .I1(n14489[3]), .I2(n378_adj_4949), 
            .I3(n39503), .O(n13768[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_6 (.CI(n39503), .I0(n14489[3]), .I1(n378_adj_4949), 
            .CO(n39504));
    SB_LUT4 add_4967_5_lut (.I0(GND_net), .I1(n14489[2]), .I2(n305_adj_4948), 
            .I3(n39502), .O(n13768[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_5 (.CI(n39502), .I0(n14489[2]), .I1(n305_adj_4948), 
            .CO(n39503));
    SB_LUT4 add_4967_4_lut (.I0(GND_net), .I1(n14489[1]), .I2(n232_adj_4947), 
            .I3(n39501), .O(n13768[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_4 (.CI(n39501), .I0(n14489[1]), .I1(n232_adj_4947), 
            .CO(n39502));
    SB_LUT4 add_4967_3_lut (.I0(GND_net), .I1(n14489[0]), .I2(n159_adj_4946), 
            .I3(n39500), .O(n13768[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_3 (.CI(n39500), .I0(n14489[0]), .I1(n159_adj_4946), 
            .CO(n39501));
    SB_LUT4 add_4967_2_lut (.I0(GND_net), .I1(n17_adj_4942), .I2(n86_adj_4940), 
            .I3(GND_net), .O(n13768[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4967_2 (.CI(GND_net), .I0(n17_adj_4942), .I1(n86_adj_4940), 
            .CO(n39500));
    SB_LUT4 add_5228_10_lut (.I0(GND_net), .I1(n18209[7]), .I2(n700_adj_4939), 
            .I3(n39499), .O(n18029[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_3 (.CI(n38265), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4236[1]), .CO(n38266));
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5080));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5079));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4823_7_lut (.I0(GND_net), .I1(n11605[4]), .I2(n442), .I3(n39327), 
            .O(n10588[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[5]), 
            .I3(n38384), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n38384), .I0(GND_net), .I1(n1_adj_5147[5]), 
            .CO(n38385));
    SB_LUT4 add_958_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4236[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3672 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5228_9_lut (.I0(GND_net), .I1(n18209[6]), .I2(n627_adj_4922), 
            .I3(n39498), .O(n18029[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_9 (.CI(n39498), .I0(n18209[6]), .I1(n627_adj_4922), 
            .CO(n39499));
    SB_LUT4 add_5228_8_lut (.I0(GND_net), .I1(n18209[5]), .I2(n554_adj_4921), 
            .I3(n39497), .O(n18029[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_8 (.CI(n39497), .I0(n18209[5]), .I1(n554_adj_4921), 
            .CO(n39498));
    SB_LUT4 add_5228_7_lut (.I0(GND_net), .I1(n18209[4]), .I2(n481_adj_4920), 
            .I3(n39496), .O(n18029[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_7 (.CI(n39496), .I0(n18209[4]), .I1(n481_adj_4920), 
            .CO(n39497));
    SB_LUT4 add_5228_6_lut (.I0(GND_net), .I1(n18209[3]), .I2(n408_adj_4919), 
            .I3(n39495), .O(n18029[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_6 (.CI(n39495), .I0(n18209[3]), .I1(n408_adj_4919), 
            .CO(n39496));
    SB_LUT4 add_5228_5_lut (.I0(GND_net), .I1(n18209[2]), .I2(n335_adj_4918), 
            .I3(n39494), .O(n18029[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_5 (.CI(n39494), .I0(n18209[2]), .I1(n335_adj_4918), 
            .CO(n39495));
    SB_LUT4 add_5228_4_lut (.I0(GND_net), .I1(n18209[1]), .I2(n262_adj_4917), 
            .I3(n39493), .O(n18029[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_4 (.CI(n39493), .I0(n18209[1]), .I1(n262_adj_4917), 
            .CO(n39494));
    SB_LUT4 add_5228_3_lut (.I0(GND_net), .I1(n18209[0]), .I2(n189_adj_4916), 
            .I3(n39492), .O(n18029[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_5078));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5228_3 (.CI(n39492), .I0(n18209[0]), .I1(n189_adj_4916), 
            .CO(n39493));
    SB_LUT4 add_5228_2_lut (.I0(GND_net), .I1(n47_adj_4915), .I2(n116_adj_4914), 
            .I3(GND_net), .O(n18029[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_7 (.CI(n39327), .I0(n11605[4]), .I1(n442), .CO(n39328));
    SB_CARRY add_5228_2 (.CI(GND_net), .I0(n47_adj_4915), .I1(n116_adj_4914), 
            .CO(n39492));
    SB_LUT4 add_5084_5_lut (.I0(GND_net), .I1(n16449[2]), .I2(n317_adj_4913), 
            .I3(n39182), .O(n15969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5003_19_lut (.I0(GND_net), .I1(n15136[16]), .I2(GND_net), 
            .I3(n39491), .O(n14489[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5003_18_lut (.I0(GND_net), .I1(n15136[15]), .I2(GND_net), 
            .I3(n39490), .O(n14489[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_18 (.CI(n39490), .I0(n15136[15]), .I1(GND_net), 
            .CO(n39491));
    SB_LUT4 add_5003_17_lut (.I0(GND_net), .I1(n15136[14]), .I2(GND_net), 
            .I3(n39489), .O(n14489[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_17 (.CI(n39489), .I0(n15136[14]), .I1(GND_net), 
            .CO(n39490));
    SB_LUT4 add_5003_16_lut (.I0(GND_net), .I1(n15136[13]), .I2(n1111_adj_4912), 
            .I3(n39488), .O(n14489[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_16 (.CI(n39488), .I0(n15136[13]), .I1(n1111_adj_4912), 
            .CO(n39489));
    SB_LUT4 add_5003_15_lut (.I0(GND_net), .I1(n15136[12]), .I2(n1038_adj_4911), 
            .I3(n39487), .O(n14489[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_15 (.CI(n39487), .I0(n15136[12]), .I1(n1038_adj_4911), 
            .CO(n39488));
    SB_LUT4 add_5003_14_lut (.I0(GND_net), .I1(n15136[11]), .I2(n965_adj_4910), 
            .I3(n39486), .O(n14489[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_14 (.CI(n39486), .I0(n15136[11]), .I1(n965_adj_4910), 
            .CO(n39487));
    SB_LUT4 add_5003_13_lut (.I0(GND_net), .I1(n15136[10]), .I2(n892_adj_4909), 
            .I3(n39485), .O(n14489[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_13 (.CI(n39485), .I0(n15136[10]), .I1(n892_adj_4909), 
            .CO(n39486));
    SB_LUT4 add_5003_12_lut (.I0(GND_net), .I1(n15136[9]), .I2(n819_adj_4908), 
            .I3(n39484), .O(n14489[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_12 (.CI(n39484), .I0(n15136[9]), .I1(n819_adj_4908), 
            .CO(n39485));
    SB_LUT4 add_5003_11_lut (.I0(GND_net), .I1(n15136[8]), .I2(n746_adj_4907), 
            .I3(n39483), .O(n14489[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_11 (.CI(n39483), .I0(n15136[8]), .I1(n746_adj_4907), 
            .CO(n39484));
    SB_LUT4 add_5003_10_lut (.I0(GND_net), .I1(n15136[7]), .I2(n673_adj_4905), 
            .I3(n39482), .O(n14489[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_10 (.CI(n39482), .I0(n15136[7]), .I1(n673_adj_4905), 
            .CO(n39483));
    SB_LUT4 add_5003_9_lut (.I0(GND_net), .I1(n15136[6]), .I2(n600_adj_4904), 
            .I3(n39481), .O(n14489[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_9 (.CI(n39481), .I0(n15136[6]), .I1(n600_adj_4904), 
            .CO(n39482));
    SB_CARRY add_5084_5 (.CI(n39182), .I0(n16449[2]), .I1(n317_adj_4913), 
            .CO(n39183));
    SB_CARRY add_958_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4236[0]), .CO(n38265));
    SB_LUT4 add_5003_8_lut (.I0(GND_net), .I1(n15136[5]), .I2(n527_adj_4903), 
            .I3(n39480), .O(n14489[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_8 (.CI(n39480), .I0(n15136[5]), .I1(n527_adj_4903), 
            .CO(n39481));
    SB_LUT4 add_5003_7_lut (.I0(GND_net), .I1(n15136[4]), .I2(n454_adj_4901), 
            .I3(n39479), .O(n14489[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_7 (.CI(n39479), .I0(n15136[4]), .I1(n454_adj_4901), 
            .CO(n39480));
    SB_LUT4 add_4823_6_lut (.I0(GND_net), .I1(n11605[3]), .I2(n369), .I3(n39326), 
            .O(n10588[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20589_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20589_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[4]), 
            .I3(n38383), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n38383), .I0(GND_net), .I1(n1_adj_5147[4]), 
            .CO(n38384));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[3]), 
            .I3(n38382), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n38382), .I0(GND_net), .I1(n1_adj_5147[3]), 
            .CO(n38383));
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n10612[0]), .I2(n10081[0]), 
            .I3(n38264), .O(duty_23__N_3772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[2]), 
            .I3(n38381), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5003_6_lut (.I0(GND_net), .I1(n15136[3]), .I2(n381_adj_4897), 
            .I3(n39478), .O(n14489[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_5077));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4823_6 (.CI(n39326), .I0(n11605[3]), .I1(n369), .CO(n39327));
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5076));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_5075));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_5074));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_5073));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20588_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20588_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n38263), .O(duty_23__N_3772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n38263), .I0(n106[22]), .I1(n155[22]), .CO(n38264));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n38381), .I0(GND_net), .I1(n1_adj_5147[2]), 
            .CO(n38382));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[1]), 
            .I3(n38380), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n38262), .O(duty_23__N_3772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n38262), .I0(n106[21]), .I1(n155[21]), .CO(n38263));
    SB_CARRY add_5003_6 (.CI(n39478), .I0(n15136[3]), .I1(n381_adj_4897), 
            .CO(n39479));
    SB_LUT4 add_4823_5_lut (.I0(GND_net), .I1(n11605[2]), .I2(n296), .I3(n39325), 
            .O(n10588[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_4_lut (.I0(GND_net), .I1(n16449[1]), .I2(n244_adj_4895), 
            .I3(n39181), .O(n15969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n38261), .O(duty_23__N_3772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n38380), .I0(GND_net), .I1(n1_adj_5147[1]), 
            .CO(n38381));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5147[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n38261), .I0(n106[20]), .I1(n155[20]), .CO(n38262));
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_5072));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n38260), .O(duty_23__N_3772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5147[0]), 
            .CO(n38380));
    SB_CARRY add_12_21 (.CI(n38260), .I0(n106[19]), .I1(n155[19]), .CO(n38261));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5146[23]), 
            .I3(n38379), .O(\PID_CONTROLLER.integral_23__N_3723 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_5146[22]), .I3(n38378), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n38378), .I0(GND_net), .I1(n1_adj_5146[22]), 
            .CO(n38379));
    SB_LUT4 add_5003_5_lut (.I0(GND_net), .I1(n15136[2]), .I2(n308), .I3(n39477), 
            .O(n14489[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_5 (.CI(n39325), .I0(n11605[2]), .I1(n296), .CO(n39326));
    SB_CARRY add_5084_4 (.CI(n39181), .I0(n16449[1]), .I1(n244_adj_4895), 
            .CO(n39182));
    SB_CARRY add_5003_5 (.CI(n39477), .I0(n15136[2]), .I1(n308), .CO(n39478));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_5146[21]), .I3(n38377), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_5070));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4823_4_lut (.I0(GND_net), .I1(n11605[1]), .I2(n223), .I3(n39324), 
            .O(n10588[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5084_3_lut (.I0(GND_net), .I1(n16449[0]), .I2(n171_adj_4885), 
            .I3(n39180), .O(n15969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_3 (.CI(n39180), .I0(n16449[0]), .I1(n171_adj_4885), 
            .CO(n39181));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n38377), .I0(GND_net), .I1(n1_adj_5146[21]), 
            .CO(n38378));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_5146[20]), .I3(n38376), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n38376), .I0(GND_net), .I1(n1_adj_5146[20]), 
            .CO(n38377));
    SB_CARRY add_4823_4 (.CI(n39324), .I0(n11605[1]), .I1(n223), .CO(n39325));
    SB_LUT4 add_5084_2_lut (.I0(GND_net), .I1(n29_adj_4883), .I2(n98_adj_4881), 
            .I3(GND_net), .O(n15969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5084_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5084_2 (.CI(GND_net), .I0(n29_adj_4883), .I1(n98_adj_4881), 
            .CO(n39180));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_5146[19]), .I3(n38375), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5113_15_lut (.I0(GND_net), .I1(n16869[12]), .I2(n1050), 
            .I3(n39179), .O(n16449[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n38375), .I0(GND_net), .I1(n1_adj_5146[19]), 
            .CO(n38376));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_5146[18]), .I3(n38374), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n38374), .I0(GND_net), .I1(n1_adj_5146[18]), 
            .CO(n38375));
    SB_LUT4 add_5003_4_lut (.I0(GND_net), .I1(n15136[1]), .I2(n235), .I3(n39476), 
            .O(n14489[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5113_14_lut (.I0(GND_net), .I1(n16869[11]), .I2(n977), 
            .I3(n39178), .O(n16449[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_3_lut (.I0(GND_net), .I1(n11605[0]), .I2(n150_adj_4874), 
            .I3(n39323), .O(n10588[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_5146[17]), .I3(n38373), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_5069));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5003_4 (.CI(n39476), .I0(n15136[1]), .I1(n235), .CO(n39477));
    SB_LUT4 add_5003_3_lut (.I0(GND_net), .I1(n15136[0]), .I2(n162), .I3(n39475), 
            .O(n14489[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_3 (.CI(n39323), .I0(n11605[0]), .I1(n150_adj_4874), 
            .CO(n39324));
    SB_LUT4 i20587_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20587_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4823_2_lut (.I0(GND_net), .I1(n8_adj_4869), .I2(n77), 
            .I3(GND_net), .O(n10588[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_2 (.CI(GND_net), .I0(n8_adj_4869), .I1(n77), .CO(n39323));
    SB_CARRY add_5003_3 (.CI(n39475), .I0(n15136[0]), .I1(n162), .CO(n39476));
    SB_LUT4 add_5003_2_lut (.I0(GND_net), .I1(n20_adj_4866), .I2(n89), 
            .I3(GND_net), .O(n14489[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5003_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5003_2 (.CI(GND_net), .I0(n20_adj_4866), .I1(n89), .CO(n39475));
    SB_LUT4 add_5037_18_lut (.I0(GND_net), .I1(n15713[15]), .I2(GND_net), 
            .I3(n39474), .O(n15136[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4868_22_lut (.I0(GND_net), .I1(n12529[19]), .I2(GND_net), 
            .I3(n39322), .O(n11605[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5113_14 (.CI(n39178), .I0(n16869[11]), .I1(n977), .CO(n39179));
    SB_LUT4 add_5037_17_lut (.I0(GND_net), .I1(n15713[14]), .I2(GND_net), 
            .I3(n39473), .O(n15136[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_17 (.CI(n39473), .I0(n15713[14]), .I1(GND_net), 
            .CO(n39474));
    SB_LUT4 add_5113_13_lut (.I0(GND_net), .I1(n16869[10]), .I2(n904_adj_4864), 
            .I3(n39177), .O(n16449[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5037_16_lut (.I0(GND_net), .I1(n15713[13]), .I2(n1114_adj_4863), 
            .I3(n39472), .O(n15136[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_16 (.CI(n39472), .I0(n15713[13]), .I1(n1114_adj_4863), 
            .CO(n39473));
    SB_LUT4 add_5037_15_lut (.I0(GND_net), .I1(n15713[12]), .I2(n1041_adj_4862), 
            .I3(n39471), .O(n15136[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n38259), .O(duty_23__N_3772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n38373), .I0(GND_net), .I1(n1_adj_5146[17]), 
            .CO(n38374));
    SB_CARRY add_12_20 (.CI(n38259), .I0(n106[18]), .I1(n155[18]), .CO(n38260));
    SB_CARRY add_5037_15 (.CI(n39471), .I0(n15713[12]), .I1(n1041_adj_4862), 
            .CO(n39472));
    SB_LUT4 add_4868_21_lut (.I0(GND_net), .I1(n12529[18]), .I2(GND_net), 
            .I3(n39321), .O(n11605[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4868_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_5146[16]), .I3(n38372), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5113_13 (.CI(n39177), .I0(n16869[10]), .I1(n904_adj_4864), 
            .CO(n39178));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n38258), .O(duty_23__N_3772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n38372), .I0(GND_net), .I1(n1_adj_5146[16]), 
            .CO(n38373));
    SB_CARRY add_12_19 (.CI(n38258), .I0(n106[17]), .I1(n155[17]), .CO(n38259));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_5146[15]), .I3(n38371), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n38371), .I0(GND_net), .I1(n1_adj_5146[15]), 
            .CO(n38372));
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_5068));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5037_14_lut (.I0(GND_net), .I1(n15713[11]), .I2(n968_adj_4859), 
            .I3(n39470), .O(n15136[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5037_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_5146[14]), .I3(n38370), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20586_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20586_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_5066));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5113_12_lut (.I0(GND_net), .I1(n16869[9]), .I2(n831), 
            .I3(n39176), .O(n16449[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5113_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5037_14 (.CI(n39470), .I0(n15713[11]), .I1(n968_adj_4859), 
            .CO(n39471));
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4891));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_5063));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_5062));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_5061));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24570_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_5084), 
            .I3(n18633[1]), .O(n6_adj_4749));   // verilog/motorControl.v(34[16:22])
    defparam i24570_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_5058));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1560 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n18633[1]), 
            .I3(n4_adj_5084), .O(n18584[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1560.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_5055));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5054));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20585_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20585_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_5052));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_5050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20584_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20584_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5049));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_5048));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_5047));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_5046));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5045));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_5043));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_5042));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4890));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_5040));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_5039));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_5038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1561 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n18633[0]), 
            .I3(n38050), .O(n18584[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1561.LUT_INIT = 16'h8778;
    SB_LUT4 i24562_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n38050), 
            .I3(n18633[0]), .O(n4_adj_5084));   // verilog/motorControl.v(34[16:22])
    defparam i24562_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_5037));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24549_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n18584[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24549_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20583_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20583_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_5036));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_5035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_5034));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_5033));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_5032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_5031));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5030));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24551_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n38050));   // verilog/motorControl.v(34[16:22])
    defparam i24551_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_5028));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_5027));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20582_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20582_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_5025));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5024));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5085));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_5022));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5086));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5087));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5088));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5089));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_5021));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5020));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5090));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5091));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_5019));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_5018));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5017));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5147[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_5014));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_5013));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_5012));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5092));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_5011));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5093));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5094));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5095));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5096));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_5010));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_5009));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5097));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5098));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_5008));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_5007));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_5006));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20581_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20581_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5099));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5100));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_5005));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5101));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5102));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_5004));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_5003));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5103));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24486_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n37968), 
            .I3(n18681[0]), .O(n4_adj_4772));   // verilog/motorControl.v(34[16:22])
    defparam i24486_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1562 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n18681[0]), 
            .I3(n37968), .O(n18664[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1562.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32313_4_lut (.I0(n21_adj_5103), .I1(n19_adj_5102), .I2(n17_adj_5101), 
            .I3(n9_adj_5100), .O(n47394));
    defparam i32313_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32306_4_lut (.I0(n27_adj_5099), .I1(n15_adj_5098), .I2(n13_adj_5097), 
            .I3(n11_adj_5096), .O(n47387));
    defparam i32306_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_5095), 
            .I3(GND_net), .O(n12_adj_5104));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_5097), 
            .I3(GND_net), .O(n10_adj_5105));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_5104), .I1(n257[17]), .I2(n35_adj_5092), 
            .I3(GND_net), .O(n30_adj_5106));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32569_4_lut (.I0(n13_adj_5097), .I1(n11_adj_5096), .I2(n9_adj_5100), 
            .I3(n47406), .O(n47650));
    defparam i32569_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32563_4_lut (.I0(n19_adj_5102), .I1(n17_adj_5101), .I2(n15_adj_5098), 
            .I3(n47650), .O(n47644));
    defparam i32563_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32890_4_lut (.I0(n25_adj_5094), .I1(n23_adj_5093), .I2(n21_adj_5103), 
            .I3(n47644), .O(n47971));
    defparam i32890_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32732_4_lut (.I0(n31_adj_5090), .I1(n29_adj_5089), .I2(n27_adj_5099), 
            .I3(n47971), .O(n47813));
    defparam i32732_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_5000));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32930_4_lut (.I0(n37_adj_5088), .I1(n35_adj_5092), .I2(n33_adj_5095), 
            .I3(n47813), .O(n48011));
    defparam i32930_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_5091), 
            .I3(GND_net), .O(n16_adj_5107));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32746_3_lut (.I0(n6_adj_4906), .I1(n257[10]), .I2(n21_adj_5103), 
            .I3(GND_net), .O(n47827));   // verilog/motorControl.v(38[19:35])
    defparam i32746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32747_3_lut (.I0(n47827), .I1(n257[11]), .I2(n23_adj_5093), 
            .I3(GND_net), .O(n47828));   // verilog/motorControl.v(38[19:35])
    defparam i32747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4999));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_5101), 
            .I3(GND_net), .O(n8_adj_5108));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_5107), .I1(n257[22]), .I2(n45_adj_5087), 
            .I3(GND_net), .O(n24_adj_5109));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32231_4_lut (.I0(n43_adj_5091), .I1(n25_adj_5094), .I2(n23_adj_5093), 
            .I3(n47394), .O(n47312));
    defparam i32231_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i20580_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20580_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20579_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20579_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32728_4_lut (.I0(n24_adj_5109), .I1(n8_adj_5108), .I2(n45_adj_5087), 
            .I3(n47310), .O(n47809));   // verilog/motorControl.v(38[19:35])
    defparam i32728_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32544_3_lut (.I0(n47828), .I1(n257[12]), .I2(n25_adj_5094), 
            .I3(GND_net), .O(n47625));   // verilog/motorControl.v(38[19:35])
    defparam i32544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(n257[1]), 
            .I2(duty_23__N_3772[1]), .I3(n257[0]), .O(n4_adj_5110));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i20578_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20578_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32742_3_lut (.I0(n4_adj_5110), .I1(n257[13]), .I2(n27_adj_5099), 
            .I3(GND_net), .O(n47823));   // verilog/motorControl.v(38[19:35])
    defparam i32742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32743_3_lut (.I0(n47823), .I1(n257[14]), .I2(n29_adj_5089), 
            .I3(GND_net), .O(n47824));   // verilog/motorControl.v(38[19:35])
    defparam i32743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4997));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32268_4_lut (.I0(n33_adj_5095), .I1(n31_adj_5090), .I2(n29_adj_5089), 
            .I3(n47387), .O(n47349));
    defparam i32268_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32948_4_lut (.I0(n30_adj_5106), .I1(n10_adj_5105), .I2(n35_adj_5092), 
            .I3(n47340), .O(n48029));   // verilog/motorControl.v(38[19:35])
    defparam i32948_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4996));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32546_3_lut (.I0(n47824), .I1(n257[15]), .I2(n31_adj_5090), 
            .I3(GND_net), .O(n47627));   // verilog/motorControl.v(38[19:35])
    defparam i32546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32986_4_lut (.I0(n47627), .I1(n48029), .I2(n35_adj_5092), 
            .I3(n47349), .O(n48067));   // verilog/motorControl.v(38[19:35])
    defparam i32986_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32987_3_lut (.I0(n48067), .I1(n257[18]), .I2(n37_adj_5088), 
            .I3(GND_net), .O(n48068));   // verilog/motorControl.v(38[19:35])
    defparam i32987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32977_3_lut (.I0(n48068), .I1(n257[19]), .I2(n39_adj_5086), 
            .I3(GND_net), .O(n48058));   // verilog/motorControl.v(38[19:35])
    defparam i32977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32234_4_lut (.I0(n43_adj_5091), .I1(n41_adj_5085), .I2(n39_adj_5086), 
            .I3(n48011), .O(n47315));
    defparam i32234_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32884_4_lut (.I0(n47625), .I1(n47809), .I2(n45_adj_5087), 
            .I3(n47312), .O(n47965));   // verilog/motorControl.v(38[19:35])
    defparam i32884_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32953_3_lut (.I0(n48058), .I1(n257[20]), .I2(n41_adj_5085), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(38[19:35])
    defparam i32953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32886_4_lut (.I0(n40), .I1(n47965), .I2(n45_adj_5087), .I3(n47315), 
            .O(n47967));   // verilog/motorControl.v(38[19:35])
    defparam i32886_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32887_3_lut (.I0(n47967), .I1(duty_23__N_3772[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4853));   // verilog/motorControl.v(38[19:35])
    defparam i32887_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3772[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5111));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4995));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4994));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3772[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5112));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3772[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5113));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4993));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3772[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5114));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5115));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4992));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4991));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3772[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5116));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3772[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5117));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i20577_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20577_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20576_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20576_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4988));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3772[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5118));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3772[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5119));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3772[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5120));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3772[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5121));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3772[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5122));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3772[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5123));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3772[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5124));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5125));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3772[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5126));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3772[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5127));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4986));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3772[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5128));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4985));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3772[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5129));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4984));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32349_4_lut (.I0(n21_adj_5129), .I1(n19_adj_5128), .I2(n17_adj_5127), 
            .I3(n9_adj_5126), .O(n47430));
    defparam i32349_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i20575_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20575_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4982));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1563 (.I0(n62), .I1(n131), .I2(n18664[0]), 
            .I3(n204), .O(n18633[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1563.LUT_INIT = 16'h8778;
    SB_LUT4 i32343_4_lut (.I0(n27_adj_5123), .I1(n15_adj_5124), .I2(n13_adj_5122), 
            .I3(n11_adj_5121), .O(n47424));
    defparam i32343_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_851_i12_3_lut (.I0(duty_23__N_3772[7]), .I1(duty_23__N_3772[16]), 
            .I2(n33_adj_5125), .I3(GND_net), .O(n12_adj_5130));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i10_3_lut (.I0(duty_23__N_3772[5]), .I1(duty_23__N_3772[6]), 
            .I2(n13_adj_5122), .I3(GND_net), .O(n10_adj_5131));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24516_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n18664[0]), 
            .O(n4_adj_4764));   // verilog/motorControl.v(34[16:22])
    defparam i24516_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 duty_23__I_851_i30_3_lut (.I0(n12_adj_5130), .I1(duty_23__N_3772[17]), 
            .I2(n35_adj_5120), .I3(GND_net), .O(n30_adj_5132));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32608_4_lut (.I0(n13_adj_5122), .I1(n11_adj_5121), .I2(n9_adj_5126), 
            .I3(n47440), .O(n47689));
    defparam i32608_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32604_4_lut (.I0(n19_adj_5128), .I1(n17_adj_5127), .I2(n15_adj_5124), 
            .I3(n47689), .O(n47685));
    defparam i32604_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32900_4_lut (.I0(n25_adj_5117), .I1(n23_adj_5116), .I2(n21_adj_5129), 
            .I3(n47685), .O(n47981));
    defparam i32900_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32756_4_lut (.I0(n31_adj_5119), .I1(n29_adj_5118), .I2(n27_adj_5123), 
            .I3(n47981), .O(n47837));
    defparam i32756_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32938_4_lut (.I0(n37_adj_5114), .I1(n35_adj_5120), .I2(n33_adj_5125), 
            .I3(n47837), .O(n48019));
    defparam i32938_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_851_i16_3_lut (.I0(duty_23__N_3772[9]), .I1(duty_23__N_3772[21]), 
            .I2(n43_adj_5115), .I3(GND_net), .O(n16_adj_5133));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20574_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20574_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24473_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n18664[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24473_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32830_3_lut (.I0(n6_adj_4902), .I1(duty_23__N_3772[10]), .I2(n21_adj_5129), 
            .I3(GND_net), .O(n47911));   // verilog/motorControl.v(36[10:25])
    defparam i32830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32831_3_lut (.I0(n47911), .I1(duty_23__N_3772[11]), .I2(n23_adj_5116), 
            .I3(GND_net), .O(n47912));   // verilog/motorControl.v(36[10:25])
    defparam i32831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4976));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4975));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4969));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20573_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20573_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4964));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20572_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20572_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24475_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n37968));   // verilog/motorControl.v(34[16:22])
    defparam i24475_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 duty_23__I_851_i8_3_lut (.I0(duty_23__N_3772[4]), .I1(duty_23__N_3772[8]), 
            .I2(n17_adj_5127), .I3(GND_net), .O(n8_adj_5134));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i24_3_lut (.I0(n16_adj_5133), .I1(duty_23__N_3772[22]), 
            .I2(n45_adj_5113), .I3(GND_net), .O(n24_adj_5135));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32329_4_lut (.I0(n43_adj_5115), .I1(n25_adj_5117), .I2(n23_adj_5116), 
            .I3(n47430), .O(n47410));
    defparam i32329_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32726_4_lut (.I0(n24_adj_5135), .I1(n8_adj_5134), .I2(n45_adj_5113), 
            .I3(n47408), .O(n47807));   // verilog/motorControl.v(36[10:25])
    defparam i32726_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i20571_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20571_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32534_3_lut (.I0(n47912), .I1(duty_23__N_3772[12]), .I2(n25_adj_5117), 
            .I3(GND_net), .O(n47615));   // verilog/motorControl.v(36[10:25])
    defparam i32534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(duty_23__N_3772[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_5136));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i32828_3_lut (.I0(n4_adj_5136), .I1(duty_23__N_3772[13]), .I2(n27_adj_5123), 
            .I3(GND_net), .O(n47909));   // verilog/motorControl.v(36[10:25])
    defparam i32828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32829_3_lut (.I0(n47909), .I1(duty_23__N_3772[14]), .I2(n29_adj_5118), 
            .I3(GND_net), .O(n47910));   // verilog/motorControl.v(36[10:25])
    defparam i32829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32339_4_lut (.I0(n33_adj_5125), .I1(n31_adj_5119), .I2(n29_adj_5118), 
            .I3(n47424), .O(n47420));
    defparam i32339_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32892_4_lut (.I0(n30_adj_5132), .I1(n10_adj_5131), .I2(n35_adj_5120), 
            .I3(n47418), .O(n47973));   // verilog/motorControl.v(36[10:25])
    defparam i32892_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32536_3_lut (.I0(n47910), .I1(duty_23__N_3772[15]), .I2(n31_adj_5119), 
            .I3(GND_net), .O(n47617));   // verilog/motorControl.v(36[10:25])
    defparam i32536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32974_4_lut (.I0(n47617), .I1(n47973), .I2(n35_adj_5120), 
            .I3(n47420), .O(n48055));   // verilog/motorControl.v(36[10:25])
    defparam i32974_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32975_3_lut (.I0(n48055), .I1(duty_23__N_3772[18]), .I2(n37_adj_5114), 
            .I3(GND_net), .O(n48056));   // verilog/motorControl.v(36[10:25])
    defparam i32975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32955_3_lut (.I0(n48056), .I1(duty_23__N_3772[19]), .I2(n39_adj_5111), 
            .I3(GND_net), .O(n48036));   // verilog/motorControl.v(36[10:25])
    defparam i32955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32331_4_lut (.I0(n43_adj_5115), .I1(n41_adj_5112), .I2(n39_adj_5111), 
            .I3(n48019), .O(n47412));
    defparam i32331_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32880_4_lut (.I0(n47615), .I1(n47807), .I2(n45_adj_5113), 
            .I3(n47410), .O(n47961));   // verilog/motorControl.v(36[10:25])
    defparam i32880_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i24503_2_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(\Kp[1] ), 
            .I3(n1[19]), .O(n18633[0]));   // verilog/motorControl.v(34[16:22])
    defparam i24503_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32542_3_lut (.I0(n48036), .I1(duty_23__N_3772[20]), .I2(n41_adj_5112), 
            .I3(GND_net), .O(n47623));   // verilog/motorControl.v(36[10:25])
    defparam i32542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32936_4_lut (.I0(n47623), .I1(n47961), .I2(n45_adj_5113), 
            .I3(n47412), .O(n48017));   // verilog/motorControl.v(36[10:25])
    defparam i32936_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32937_3_lut (.I0(n48017), .I1(PWMLimit[23]), .I2(duty_23__N_3772[23]), 
            .I3(GND_net), .O(duty_23__N_3771));   // verilog/motorControl.v(36[10:25])
    defparam i32937_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4960));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20570_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20570_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4958));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3772[0]), .I1(n257[0]), .I2(n256_adj_4853), 
            .I3(GND_net), .O(duty_23__N_3747[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3747[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4957));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20569_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20569_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_5137));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_5138));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_5139));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32432_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n47513));
    defparam i32432_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i32430_3_lut (.I0(n11_adj_5139), .I1(n9_adj_5138), .I2(n47513), 
            .I3(GND_net), .O(n47511));
    defparam i32430_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_376_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n49340));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_376_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32794_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n49340), 
            .I2(IntegralLimit[7]), .I3(n47511), .O(n47875));
    defparam i32794_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32668_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_5137), 
            .I2(IntegralLimit[9]), .I3(n47875), .O(n47749));
    defparam i32668_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_358_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n49322));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_358_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32666_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_5137), 
            .I2(IntegralLimit[9]), .I3(n9_adj_5138), .O(n47747));
    defparam i32666_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32664_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n49322), 
            .I2(IntegralLimit[11]), .I3(n47747), .O(n47745));
    defparam i32664_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_352_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n49316));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_352_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32381_4_lut (.I0(n27), .I1(n15_adj_4784), .I2(n13), .I3(n11_adj_4811), 
            .O(n47462));
    defparam i32381_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32387_4_lut (.I0(n21), .I1(n19_adj_4777), .I2(n17_adj_4781), 
            .I3(n9_adj_4813), .O(n47468));
    defparam i32387_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_5140));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32361_2_lut (.I0(n43), .I1(n19_adj_4777), .I2(GND_net), .I3(GND_net), 
            .O(n47442));
    defparam i32361_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4781), .I3(GND_net), 
            .O(n8));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_5140), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32397_2_lut (.I0(n7), .I1(n5_adj_4838), .I2(GND_net), .I3(GND_net), 
            .O(n47478));
    defparam i32397_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32640_4_lut (.I0(n13), .I1(n11_adj_4811), .I2(n9_adj_4813), 
            .I3(n47478), .O(n47721));
    defparam i32640_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32636_4_lut (.I0(n19_adj_4777), .I1(n17_adj_4781), .I2(n15_adj_4784), 
            .I3(n47721), .O(n47717));
    defparam i32636_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32910_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n47717), 
            .O(n47991));
    defparam i32910_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32772_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n47991), 
            .O(n47853));
    defparam i32772_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32942_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n47853), 
            .O(n48023));
    defparam i32942_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32670_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n49340), 
            .I2(IntegralLimit[7]), .I3(n11_adj_5139), .O(n47751));
    defparam i32670_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5146[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_345_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n49309));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_345_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32658_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n49309), 
            .I2(IntegralLimit[14]), .I3(n47751), .O(n47739));
    defparam i32658_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_340_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n49304));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_340_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_5141));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32410_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47491));
    defparam i32410_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4733));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4795));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_5141), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4732));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32858_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n49322), 
            .I2(IntegralLimit[11]), .I3(n47749), .O(n47939));
    defparam i32858_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32418_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n49316), 
            .I2(IntegralLimit[13]), .I3(n47939), .O(n47499));
    defparam i32418_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_343_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n49307));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_343_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32788_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n49307), 
            .I2(IntegralLimit[15]), .I3(n47499), .O(n47869));
    defparam i32788_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_369_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n49333));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_369_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32914_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n49333), 
            .I2(IntegralLimit[17]), .I3(n47869), .O(n47995));
    defparam i32914_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_334_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n49298));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_334_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32966_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n49298), 
            .I2(IntegralLimit[19]), .I3(n47995), .O(n48047));
    defparam i32966_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_331_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n49295));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_331_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_5142));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32399_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n47480));
    defparam i32399_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_327_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n49291));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_327_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_5142), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_5143));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i8_4_lut_adj_1564 (.I0(n6_adj_4945), .I1(n11_adj_4944), .I2(n8_adj_4943), 
            .I3(n12_adj_4941), .O(n18));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_5144));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32846_3_lut (.I0(n6_adj_5144), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n47927));   // verilog/motorControl.v(31[10:34])
    defparam i32846_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32847_3_lut (.I0(n47927), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n47928));   // verilog/motorControl.v(31[10:34])
    defparam i32847_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32401_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n49316), 
            .I2(IntegralLimit[21]), .I3(n47745), .O(n47482));
    defparam i32401_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i32722_4_lut (.I0(n24_adj_5143), .I1(n8_adj_4937), .I2(n49291), 
            .I3(n47480), .O(n47803));   // verilog/motorControl.v(31[10:34])
    defparam i32722_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32514_3_lut (.I0(n47928), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n47595));   // verilog/motorControl.v(31[10:34])
    defparam i32514_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3723 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4840), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_5145));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i32836_3_lut (.I0(n4_adj_5145), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n47917));   // verilog/motorControl.v(31[38:63])
    defparam i32836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32837_3_lut (.I0(n47917), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n47918));   // verilog/motorControl.v(31[38:63])
    defparam i32837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4794));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32373_2_lut (.I0(n33), .I1(n15_adj_4784), .I2(GND_net), .I3(GND_net), 
            .O(n47454));
    defparam i32373_2_lut.LUT_INIT = 16'heeee;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (b_prev, GND_net, a_new, direction_N_3907, 
            ENCODER0_B_N_keep, n1668, ENCODER0_A_N_keep, encoder0_position, 
            VCC_net, n28376, n1632) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3907;
    input ENCODER0_B_N_keep;
    input n1668;
    input ENCODER0_A_N_keep;
    output [31:0]encoder0_position;
    input VCC_net;
    input n28376;
    output n1632;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3910, debounce_cnt, a_prev;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_3913;
    wire [31:0]n133;
    
    wire direction_N_3906, n39086, n39085, n39084, n39083, n39082, 
        n39081, n39080, n39079, n39078, n39077, n39076, n39075, 
        n39074, n39073, n39072, n39071, n39070, n39069, n39068, 
        n39067, n39066, n39065, n39064, n39063, n39062, n39061, 
        n39060, n39059, n39058, n39057, n39056, n28375, n28374;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 i33021_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i33021_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2202_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[31]), .I3(n39086), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2202_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[30]), .I3(n39085), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_32 (.CI(n39085), .I0(direction_N_3906), 
            .I1(encoder0_position[30]), .CO(n39086));
    SB_LUT4 position_2202_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[29]), .I3(n39084), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_31 (.CI(n39084), .I0(direction_N_3906), 
            .I1(encoder0_position[29]), .CO(n39085));
    SB_LUT4 position_2202_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[28]), .I3(n39083), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_30 (.CI(n39083), .I0(direction_N_3906), 
            .I1(encoder0_position[28]), .CO(n39084));
    SB_LUT4 position_2202_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[27]), .I3(n39082), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_29 (.CI(n39082), .I0(direction_N_3906), 
            .I1(encoder0_position[27]), .CO(n39083));
    SB_LUT4 position_2202_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[26]), .I3(n39081), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_28 (.CI(n39081), .I0(direction_N_3906), 
            .I1(encoder0_position[26]), .CO(n39082));
    SB_LUT4 position_2202_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[25]), .I3(n39080), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_27 (.CI(n39080), .I0(direction_N_3906), 
            .I1(encoder0_position[25]), .CO(n39081));
    SB_LUT4 position_2202_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[24]), .I3(n39079), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_26 (.CI(n39079), .I0(direction_N_3906), 
            .I1(encoder0_position[24]), .CO(n39080));
    SB_LUT4 position_2202_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[23]), .I3(n39078), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_25 (.CI(n39078), .I0(direction_N_3906), 
            .I1(encoder0_position[23]), .CO(n39079));
    SB_LUT4 position_2202_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[22]), .I3(n39077), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_24 (.CI(n39077), .I0(direction_N_3906), 
            .I1(encoder0_position[22]), .CO(n39078));
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2202_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[21]), .I3(n39076), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_23 (.CI(n39076), .I0(direction_N_3906), 
            .I1(encoder0_position[21]), .CO(n39077));
    SB_LUT4 position_2202_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[20]), .I3(n39075), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY position_2202_add_4_22 (.CI(n39075), .I0(direction_N_3906), 
            .I1(encoder0_position[20]), .CO(n39076));
    SB_LUT4 position_2202_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[19]), .I3(n39074), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_21 (.CI(n39074), .I0(direction_N_3906), 
            .I1(encoder0_position[19]), .CO(n39075));
    SB_LUT4 position_2202_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[18]), .I3(n39073), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_20 (.CI(n39073), .I0(direction_N_3906), 
            .I1(encoder0_position[18]), .CO(n39074));
    SB_LUT4 position_2202_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[17]), .I3(n39072), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_19 (.CI(n39072), .I0(direction_N_3906), 
            .I1(encoder0_position[17]), .CO(n39073));
    SB_LUT4 position_2202_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[16]), .I3(n39071), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_18 (.CI(n39071), .I0(direction_N_3906), 
            .I1(encoder0_position[16]), .CO(n39072));
    SB_LUT4 position_2202_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[15]), .I3(n39070), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_17 (.CI(n39070), .I0(direction_N_3906), 
            .I1(encoder0_position[15]), .CO(n39071));
    SB_LUT4 position_2202_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[14]), .I3(n39069), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_16 (.CI(n39069), .I0(direction_N_3906), 
            .I1(encoder0_position[14]), .CO(n39070));
    SB_LUT4 position_2202_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[13]), .I3(n39068), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_15 (.CI(n39068), .I0(direction_N_3906), 
            .I1(encoder0_position[13]), .CO(n39069));
    SB_LUT4 position_2202_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[12]), .I3(n39067), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_14 (.CI(n39067), .I0(direction_N_3906), 
            .I1(encoder0_position[12]), .CO(n39068));
    SB_LUT4 position_2202_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[11]), .I3(n39066), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_13 (.CI(n39066), .I0(direction_N_3906), 
            .I1(encoder0_position[11]), .CO(n39067));
    SB_LUT4 position_2202_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[10]), .I3(n39065), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_12 (.CI(n39065), .I0(direction_N_3906), 
            .I1(encoder0_position[10]), .CO(n39066));
    SB_LUT4 position_2202_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[9]), .I3(n39064), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_11 (.CI(n39064), .I0(direction_N_3906), 
            .I1(encoder0_position[9]), .CO(n39065));
    SB_LUT4 position_2202_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[8]), .I3(n39063), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_10 (.CI(n39063), .I0(direction_N_3906), 
            .I1(encoder0_position[8]), .CO(n39064));
    SB_LUT4 position_2202_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[7]), .I3(n39062), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_9 (.CI(n39062), .I0(direction_N_3906), 
            .I1(encoder0_position[7]), .CO(n39063));
    SB_LUT4 position_2202_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[6]), .I3(n39061), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_8 (.CI(n39061), .I0(direction_N_3906), 
            .I1(encoder0_position[6]), .CO(n39062));
    SB_LUT4 position_2202_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[5]), .I3(n39060), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_7 (.CI(n39060), .I0(direction_N_3906), 
            .I1(encoder0_position[5]), .CO(n39061));
    SB_LUT4 position_2202_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[4]), .I3(n39059), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_6 (.CI(n39059), .I0(direction_N_3906), 
            .I1(encoder0_position[4]), .CO(n39060));
    SB_LUT4 position_2202_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[3]), .I3(n39058), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_5 (.CI(n39058), .I0(direction_N_3906), 
            .I1(encoder0_position[3]), .CO(n39059));
    SB_LUT4 position_2202_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[2]), .I3(n39057), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_4 (.CI(n39057), .I0(direction_N_3906), 
            .I1(encoder0_position[2]), .CO(n39058));
    SB_LUT4 position_2202_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[1]), .I3(n39056), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_3 (.CI(n39056), .I0(direction_N_3906), 
            .I1(encoder0_position[1]), .CO(n39057));
    SB_LUT4 position_2202_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n39056));
    SB_DFFE position_2202__i31 (.Q(encoder0_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i30 (.Q(encoder0_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i29 (.Q(encoder0_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i28 (.Q(encoder0_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i27 (.Q(encoder0_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i26 (.Q(encoder0_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i25 (.Q(encoder0_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i24 (.Q(encoder0_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i23 (.Q(encoder0_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i22 (.Q(encoder0_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i21 (.Q(encoder0_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i20 (.Q(encoder0_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i19 (.Q(encoder0_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i18 (.Q(encoder0_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i17 (.Q(encoder0_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i16 (.Q(encoder0_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i15 (.Q(encoder0_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i14 (.Q(encoder0_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i13 (.Q(encoder0_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i12 (.Q(encoder0_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i11 (.Q(encoder0_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i10 (.Q(encoder0_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i9 (.Q(encoder0_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i8 (.Q(encoder0_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i7 (.Q(encoder0_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i6 (.Q(encoder0_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i5 (.Q(encoder0_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i4 (.Q(encoder0_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i3 (.Q(encoder0_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i2 (.Q(encoder0_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i1 (.Q(encoder0_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i0 (.Q(encoder0_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1632), .C(n1668), .D(n28376));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n28375));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n28374));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i14864_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n28375));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14863_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n28374));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14863_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n28234, \data_out_frame[13] , CLK_c, n28233, n26879, 
            n28232, \data_out_frame[14] , n28231, n28230, GND_net, 
            n28229, n28228, n28227, n28226, n28225, \data_out_frame[6] , 
            \data_out_frame[7] , \data_out_frame[4] , \data_out_frame[5] , 
            \FRAME_MATCHER.state , \data_out_frame[16] , \data_out_frame[17] , 
            \data_out_frame[18] , \data_out_frame[19] , \data_out_frame[22] , 
            \data_out_frame[23] , \data_out_frame[20] , \data_out_frame[21][4] , 
            \data_out_frame[25] , \data_out_frame[15] , \data_out_frame[24] , 
            rx_data_ready, n28224, n28223, \data_out_frame[10] , n27595, 
            \data_out_frame[12] , \data_out_frame[21][2] , n9, n3813, 
            n4452, n23534, n29908, \FRAME_MATCHER.i_31__N_2626 , \data_in[0] , 
            \data_in[1] , \data_in[2] , \data_in[3] , n28222, n28221, 
            n3303, n63, \FRAME_MATCHER.i_31__N_2624 , \FRAME_MATCHER.i_31__N_2622 , 
            \data_out_frame[8] , \data_out_frame[9] , \data_out_frame[11] , 
            setpoint, n28220, n28219, n28218, n28217, n28216, n28215, 
            n28214, n28213, n28212, n28211, n28210, n28209, n28208, 
            n28207, n27596, n28206, \data_in_frame[5] , n28205, \data_out_frame[21][1] , 
            \data_in_frame[3] , n28204, \data_in_frame[2] , n28203, 
            n28202, \data_out_frame[21][0] , \data_in_frame[1] , \data_out_frame[21][3] , 
            tx_active, n28200, n36539, n28199, n28198, n28197, n28196, 
            n28195, n28194, n28193, n28192, n28191, n28190, n28189, 
            n28188, n28187, n28186, n28185, n28184, n28183, n28182, 
            n28181, n28180, \data_out_frame[27][1] , ID, n28179, n28178, 
            rx_data, \data_in_frame[8] , \data_in_frame[11] , \data_in_frame[13] , 
            \data_in_frame[9] , n122, n5, n49229, \data_in_frame[10] , 
            \data_in_frame[4] , n28177, \data_in_frame[6] , n28176, 
            n28175, n28715, n28714, n28713, n28712, n28711, n28710, 
            neopxl_color, n28709, n28708, n28707, n28706, n28705, 
            n28704, n28703, n28702, n28701, n28700, n28699, n28698, 
            n28697, n28696, n28695, n28694, n28693, n28692, n28691, 
            n28690, n28689, n28688, n28687, n28686, n28685, n28684, 
            n28683, n28174, n28173, n28172, n28171, n28170, n28169, 
            n28168, n28167, n28166, n28165, n28164, n28163, n28162, 
            n28161, n28160, n28156, n28152, n28151, n42180, n28149, 
            PWMLimit, n28148, control_mode, n28146, n28145, \Ki[0] , 
            n28144, \Kp[0] , n28143, DE_c, LED_c, n28682, n28681, 
            n28680, n28662, n28661, \Kp[1] , \data_in_frame[12] , 
            n28638, n28637, n28636, n28635, \Kp[2] , n28634, n28633, 
            n28632, n49000, n28630, n28629, n28109, IntegralLimit, 
            n28106, n28105, n28104, n28103, n28102, n28101, n28100, 
            n28099, n28098, n28097, n28095, n28094, n28093, n28092, 
            n4, n7, n28091, n27804, n28090, n28089, n28088, n28545, 
            \Kp[3] , n28544, \Kp[4] , n28534, \Kp[5] , n28516, n28515, 
            n28514, n28513, n28512, n28511, n28510, n28509, n28452, 
            \data_in_frame[21] , n28451, n28450, n28449, n28448, n28447, 
            n28446, n28445, n28438, n28437, n28433, n28432, n28431, 
            n28430, n28429, n28428, n28426, n28425, n28424, n28423, 
            n28422, n28421, n28420, n28416, \Kp[6] , n28415, n28414, 
            n28413, n28412, n28411, n28410, n28409, n28408, n28407, 
            \Kp[7] , n28406, \Kp[8] , n28405, \Kp[9] , n28404, \Kp[10] , 
            n28403, \Kp[11] , n28402, \Kp[12] , n28401, \Kp[13] , 
            n28400, \Kp[14] , n28399, \Kp[15] , n28398, \Ki[1] , 
            n28397, \Ki[2] , n28396, \Ki[3] , n28395, \Ki[4] , n28394, 
            \Ki[5] , n28393, \Ki[6] , n28392, \Ki[7] , n28391, \Ki[8] , 
            n28390, \Ki[9] , n28389, \Ki[10] , n28388, \Ki[11] , 
            n28387, \Ki[12] , n28386, \Ki[13] , n28385, \Ki[14] , 
            n28384, \Ki[15] , n28383, n28382, n28381, n28380, n28379, 
            n28378, n28377, n28373, n28361, n28360, n28359, n28358, 
            n28357, n28356, n28355, n28354, n28353, n28352, n28351, 
            n28350, n28349, n28348, n28347, n28346, n28345, n28344, 
            n28343, n28342, n28341, n28340, n28339, n28338, n28337, 
            n28336, n28335, n28329, n28328, n28327, n28326, n28325, 
            n28324, n28323, n28322, n28321, n28320, n28319, n28318, 
            n28317, n28316, n28315, n28314, n28313, n28312, n28311, 
            n28310, n28309, n28308, n28307, n28306, n28305, n28304, 
            n28303, n28302, n28301, n28300, n28299, n28298, n28297, 
            n42822, n28296, n28295, n28294, n28293, n28292, n28291, 
            n28290, n28289, n28288, n28287, n28286, n28285, n28284, 
            n28283, n28282, n28281, n28280, n28279, n28278, n28277, 
            n28276, n28275, n28274, n28273, n28272, n28271, n28270, 
            n28269, n28268, n28267, n28266, n28262, n28261, n28260, 
            n28258, n28257, n42836, n28256, n28255, n28254, n28253, 
            n28252, n28251, n42843, n28250, n28249, n28248, n28247, 
            n28246, n28245, n28243, n28242, n28241, n28240, n28239, 
            n28087, n28238, n28237, n28236, n28235, n43608, n42830, 
            n23568, \state[0] , \state[3] , \state[2] , n7233, \r_SM_Main_2__N_3613[1] , 
            r_SM_Main, n18940, \r_Bit_Index[0] , tx_o, n27763, n28054, 
            VCC_net, n48986, n28365, n28159, n4_adj_10, tx_enable, 
            \r_Bit_Index[0]_adj_11 , n27767, r_SM_Main_adj_18, n28056, 
            \r_SM_Main_2__N_3542[2] , r_Rx_Data, n26339, n26334, n33899, 
            RX_N_10, n28368, n42422, n28142, n28141, n28140, n28139, 
            n28138, n28128, n28127, n42722, n4_adj_15, n4_adj_16, 
            n4_adj_17, n28372) /* synthesis syn_module_defined=1 */ ;
    input n28234;
    output [7:0]\data_out_frame[13] ;
    input CLK_c;
    input n28233;
    output n26879;
    input n28232;
    output [7:0]\data_out_frame[14] ;
    input n28231;
    input n28230;
    input GND_net;
    input n28229;
    input n28228;
    input n28227;
    input n28226;
    input n28225;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output [31:0]\FRAME_MATCHER.state ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output \data_out_frame[21][4] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[24] ;
    output rx_data_ready;
    input n28224;
    input n28223;
    output [7:0]\data_out_frame[10] ;
    output n27595;
    output [7:0]\data_out_frame[12] ;
    output \data_out_frame[21][2] ;
    input n9;
    output n3813;
    output n4452;
    output n23534;
    output n29908;
    output \FRAME_MATCHER.i_31__N_2626 ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    input n28222;
    input n28221;
    output n3303;
    output n63;
    output \FRAME_MATCHER.i_31__N_2624 ;
    output \FRAME_MATCHER.i_31__N_2622 ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[11] ;
    output [23:0]setpoint;
    input n28220;
    input n28219;
    input n28218;
    input n28217;
    input n28216;
    input n28215;
    input n28214;
    input n28213;
    input n28212;
    input n28211;
    input n28210;
    input n28209;
    input n28208;
    input n28207;
    output n27596;
    input n28206;
    output [7:0]\data_in_frame[5] ;
    input n28205;
    output \data_out_frame[21][1] ;
    output [7:0]\data_in_frame[3] ;
    input n28204;
    output [7:0]\data_in_frame[2] ;
    input n28203;
    input n28202;
    output \data_out_frame[21][0] ;
    output [7:0]\data_in_frame[1] ;
    output \data_out_frame[21][3] ;
    output tx_active;
    input n28200;
    output n36539;
    input n28199;
    input n28198;
    input n28197;
    input n28196;
    input n28195;
    input n28194;
    input n28193;
    input n28192;
    input n28191;
    input n28190;
    input n28189;
    input n28188;
    input n28187;
    input n28186;
    input n28185;
    input n28184;
    input n28183;
    input n28182;
    input n28181;
    input n28180;
    output \data_out_frame[27][1] ;
    input [7:0]ID;
    input n28179;
    input n28178;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[9] ;
    output n122;
    output n5;
    output n49229;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[4] ;
    input n28177;
    output [7:0]\data_in_frame[6] ;
    input n28176;
    input n28175;
    input n28715;
    input n28714;
    input n28713;
    input n28712;
    input n28711;
    input n28710;
    output [23:0]neopxl_color;
    input n28709;
    input n28708;
    input n28707;
    input n28706;
    input n28705;
    input n28704;
    input n28703;
    input n28702;
    input n28701;
    input n28700;
    input n28699;
    input n28698;
    input n28697;
    input n28696;
    input n28695;
    input n28694;
    input n28693;
    input n28692;
    input n28691;
    input n28690;
    input n28689;
    input n28688;
    input n28687;
    input n28686;
    input n28685;
    input n28684;
    input n28683;
    input n28174;
    input n28173;
    input n28172;
    input n28171;
    input n28170;
    input n28169;
    input n28168;
    input n28167;
    input n28166;
    input n28165;
    input n28164;
    input n28163;
    input n28162;
    input n28161;
    input n28160;
    input n28156;
    input n28152;
    input n28151;
    input n42180;
    input n28149;
    output [23:0]PWMLimit;
    input n28148;
    output [7:0]control_mode;
    input n28146;
    input n28145;
    output \Ki[0] ;
    input n28144;
    output \Kp[0] ;
    input n28143;
    output DE_c;
    output LED_c;
    input n28682;
    input n28681;
    input n28680;
    input n28662;
    input n28661;
    output \Kp[1] ;
    output [7:0]\data_in_frame[12] ;
    input n28638;
    input n28637;
    input n28636;
    input n28635;
    output \Kp[2] ;
    input n28634;
    input n28633;
    input n28632;
    input n49000;
    input n28630;
    input n28629;
    input n28109;
    output [23:0]IntegralLimit;
    input n28106;
    input n28105;
    input n28104;
    input n28103;
    input n28102;
    input n28101;
    input n28100;
    input n28099;
    input n28098;
    input n28097;
    input n28095;
    input n28094;
    input n28093;
    input n28092;
    output n4;
    output n7;
    input n28091;
    output n27804;
    input n28090;
    input n28089;
    input n28088;
    input n28545;
    output \Kp[3] ;
    input n28544;
    output \Kp[4] ;
    input n28534;
    output \Kp[5] ;
    input n28516;
    input n28515;
    input n28514;
    input n28513;
    input n28512;
    input n28511;
    input n28510;
    input n28509;
    input n28452;
    output [7:0]\data_in_frame[21] ;
    input n28451;
    input n28450;
    input n28449;
    input n28448;
    input n28447;
    input n28446;
    input n28445;
    input n28438;
    input n28437;
    input n28433;
    input n28432;
    input n28431;
    input n28430;
    input n28429;
    input n28428;
    input n28426;
    input n28425;
    input n28424;
    input n28423;
    input n28422;
    input n28421;
    input n28420;
    input n28416;
    output \Kp[6] ;
    input n28415;
    input n28414;
    input n28413;
    input n28412;
    input n28411;
    input n28410;
    input n28409;
    input n28408;
    input n28407;
    output \Kp[7] ;
    input n28406;
    output \Kp[8] ;
    input n28405;
    output \Kp[9] ;
    input n28404;
    output \Kp[10] ;
    input n28403;
    output \Kp[11] ;
    input n28402;
    output \Kp[12] ;
    input n28401;
    output \Kp[13] ;
    input n28400;
    output \Kp[14] ;
    input n28399;
    output \Kp[15] ;
    input n28398;
    output \Ki[1] ;
    input n28397;
    output \Ki[2] ;
    input n28396;
    output \Ki[3] ;
    input n28395;
    output \Ki[4] ;
    input n28394;
    output \Ki[5] ;
    input n28393;
    output \Ki[6] ;
    input n28392;
    output \Ki[7] ;
    input n28391;
    output \Ki[8] ;
    input n28390;
    output \Ki[9] ;
    input n28389;
    output \Ki[10] ;
    input n28388;
    output \Ki[11] ;
    input n28387;
    output \Ki[12] ;
    input n28386;
    output \Ki[13] ;
    input n28385;
    output \Ki[14] ;
    input n28384;
    output \Ki[15] ;
    input n28383;
    input n28382;
    input n28381;
    input n28380;
    input n28379;
    input n28378;
    input n28377;
    input n28373;
    input n28361;
    input n28360;
    input n28359;
    input n28358;
    input n28357;
    input n28356;
    input n28355;
    input n28354;
    input n28353;
    input n28352;
    input n28351;
    input n28350;
    input n28349;
    input n28348;
    input n28347;
    input n28346;
    input n28345;
    input n28344;
    input n28343;
    input n28342;
    input n28341;
    input n28340;
    input n28339;
    input n28338;
    input n28337;
    input n28336;
    input n28335;
    input n28329;
    input n28328;
    input n28327;
    input n28326;
    input n28325;
    input n28324;
    input n28323;
    input n28322;
    input n28321;
    input n28320;
    input n28319;
    input n28318;
    input n28317;
    input n28316;
    input n28315;
    input n28314;
    input n28313;
    input n28312;
    input n28311;
    input n28310;
    input n28309;
    input n28308;
    input n28307;
    input n28306;
    input n28305;
    input n28304;
    input n28303;
    input n28302;
    input n28301;
    input n28300;
    input n28299;
    input n28298;
    input n28297;
    output n42822;
    input n28296;
    input n28295;
    input n28294;
    input n28293;
    input n28292;
    input n28291;
    input n28290;
    input n28289;
    input n28288;
    input n28287;
    input n28286;
    input n28285;
    input n28284;
    input n28283;
    input n28282;
    input n28281;
    input n28280;
    input n28279;
    input n28278;
    input n28277;
    input n28276;
    input n28275;
    input n28274;
    input n28273;
    input n28272;
    input n28271;
    input n28270;
    input n28269;
    input n28268;
    input n28267;
    input n28266;
    input n28262;
    input n28261;
    input n28260;
    input n28258;
    input n28257;
    output n42836;
    input n28256;
    input n28255;
    input n28254;
    input n28253;
    input n28252;
    input n28251;
    output n42843;
    input n28250;
    input n28249;
    input n28248;
    input n28247;
    input n28246;
    input n28245;
    input n28243;
    input n28242;
    input n28241;
    input n28240;
    input n28239;
    input n28087;
    input n28238;
    input n28237;
    input n28236;
    input n28235;
    input n43608;
    output n42830;
    output n23568;
    input \state[0] ;
    input \state[3] ;
    input \state[2] ;
    output n7233;
    output \r_SM_Main_2__N_3613[1] ;
    output [2:0]r_SM_Main;
    output n18940;
    output \r_Bit_Index[0] ;
    output tx_o;
    output n27763;
    output n28054;
    input VCC_net;
    input n48986;
    input n28365;
    input n28159;
    output n4_adj_10;
    output tx_enable;
    output \r_Bit_Index[0]_adj_11 ;
    output n27767;
    output [2:0]r_SM_Main_adj_18;
    output n28056;
    output \r_SM_Main_2__N_3542[2] ;
    output r_Rx_Data;
    output n26339;
    output n26334;
    output n33899;
    input RX_N_10;
    input n28368;
    input n42422;
    input n28142;
    input n28141;
    input n28140;
    input n28139;
    input n28138;
    input n28128;
    input n28127;
    input n42722;
    output n4_adj_15;
    output n4_adj_16;
    output n4_adj_17;
    input n28372;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n57, n59, n58, n60, n69, n61, n68, n62;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3846, n3, n2, n3_adj_4435, n2_adj_4436, n3_adj_4437, n3_adj_4438;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n46314, n46315, n46313, n141, n43606, n34377, n45195, 
        n7001, n23743, n3_adj_4439, n4_c;
    wire [31:0]\FRAME_MATCHER.state_31__N_2724 ;
    
    wire n16, n4_adj_4440, n34628, n44876, n48951, n47240, n46308, 
        n46309, n46307, n48957, n47249, n46391, n46392, n46332, 
        n46331, n46281, n46280, n48981, n47236, n40416, n40271, 
        n42861, n6, n44663, n41102, n6_adj_4441, n45100, n43263, 
        n6_adj_4442, n44071, n27326, n43290, n41232, n12, n43450, 
        n43435, n42871, n44066, n43168, n27031, n27010, n43395, 
        n10, n2134, n43154, n40935, n44246, n43438, n43197, n43266, 
        n44073, n41175, n40257, n6_adj_4443, n44687, \FRAME_MATCHER.rx_data_ready_prev , 
        n161, n43368, n6_adj_4444, n45206, n45042, n43190, n6_adj_4445, 
        n41236, n14, n41104, n10_adj_4446, n44272, n40830, n43514;
    wire [7:0]n8825;
    
    wire n27621, n28080, n43407, n45249, n41137, n14_adj_4447, n43362, 
        n43074, n15, n41109, n41208, n43999, n27241, n43199, n12_adj_4448, 
        n43411, n40829, n44713, n40210, n40307, n44637, n41135, 
        n41204, n6_adj_4449, n44012, n26801, n43462, n14_adj_4450, 
        n130, n110, n2_adj_4451, n43305, n1516, n15_adj_4452, n10_adj_4453, 
        n43209, n14_adj_4454, n43187, n27484, n40355, n41177, n43206, 
        n42944, n43278, n43441, n10_adj_4455, n43216, n43420, n10_adj_4456, 
        n40347, n43254, n1, n42849, n81, n8, n43600, n10_adj_4457;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(112[11:16])
    
    wire n21657, n7_c, n34544, n19789, tx_transmit_N_3513, n29859, 
        n26449, n3065, n11, n8_adj_4458, n26350, n7_adj_4459, n5_c, 
        n771, \FRAME_MATCHER.i_31__N_2620 , n14_adj_4460, n26425, n15_adj_4461, 
        n26245, n16_adj_4462, n17, n26347, n10_adj_4463, n10_adj_4464, 
        n14_adj_4465, n26422, n18, n20, n15_adj_4466, n63_c, n16_adj_4467, 
        n17_adj_4468, n63_adj_4469, n44, n42, n43, n41, n40, n39, 
        n50, n2_adj_4470, n45, n26232, n8_adj_4471, n20_adj_4472, 
        n1_adj_4473, n19, n46207;
    wire [31:0]n92;
    
    wire n5_adj_4475, n46187, n42122, n39751, n1_adj_4476, n48985, 
        n2_adj_4477, n46451, n46452, n46341, n46340, n46343, n46344, 
        n46434, n46433, n3_adj_4478, n46352, n3_adj_4479, n46353, 
        n3_adj_4480, n46428, n46427, n46379, n3_adj_4481, n46380, 
        n46410, n46409, n3_adj_4482, n46385, n46386, n46374, n46373, 
        n46394, n46395, n2_adj_4483, n3_adj_4484, n2_adj_4485, n3_adj_4486, 
        n2_adj_4487, n3_adj_4488, n2_adj_4489, n3_adj_4490, n46296, 
        n2_adj_4491, n3_adj_4492, n46295, n2_adj_4493, n3_adj_4494, 
        n2_adj_4495, n3_adj_4496, n2_adj_4497, n3_adj_4498, n2_adj_4499, 
        n3_adj_4500;
    wire [0:0]n4888;
    wire [2:0]r_SM_Main_2__N_3616;
    
    wire n43770, n2_adj_4501, n3_adj_4502, n2_adj_4503, n3_adj_4504, 
        n7002, n27605, n2_adj_4505, n3_adj_4506, n2_adj_4507, n3_adj_4508, 
        n2_adj_4509, n3_adj_4510, n2_adj_4511, n3_adj_4512, n2_adj_4513, 
        n3_adj_4514, n2_adj_4515, n3_adj_4516, n2_adj_4517, n3_adj_4518, 
        n2_adj_4519, n3_adj_4520, n10_adj_4521, n2_adj_4522, n3_adj_4523, 
        n2_adj_4524, n3_adj_4525, n2_adj_4526, n3_adj_4527, n46397, 
        n46398, n2_adj_4528, n3_adj_4529, n2_adj_4530, n2_adj_4531, 
        n2_adj_4532, n2_adj_4533, n12_adj_4534, n42707, n4_adj_4535, 
        n42854, n133, n31, n43499, n44262, n10_adj_4536, n2_adj_4537, 
        n43350;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n43117, n8_adj_4538, n43269;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n7003, n41115, n7004, n7005, n7006, n7007, n7008, n7009;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n7010, n7011, n7012, n7013, n10_adj_4539, n7014, n7015, 
        n7016, n7017, n43080, n43353, n6_adj_4540;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n7018, n42174, n7019, n7020, n7021;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire Kp_23__N_969, n42941, n7022, n7023, n43068, n7024, n7025, 
        n43088, n27122, n12_adj_4541, n43248, n43365, n25950, n44678, 
        n43383, n14_adj_4542, n43493, n15_adj_4543, n27090, n26855, 
        n4_adj_4544, n53, n42978, n6_adj_4545, n46302, n48963, n47254, 
        n46275, n20_adj_4546, n43196, n46301, n48783, n46276, n46413, 
        n7_adj_4547, n48831, n46412;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n48969, n47227, n46455, n20_adj_4548, n26832, n27522, n33792, 
        n46294, n46292, n48867, n46456, n46407, n7_adj_4549, n48837, 
        n46406, n43423, n1191, n43302, n15_adj_4550, n14_adj_4551, 
        n38241, n48975, n47229, n46446, n42858, n20_adj_4552, n46288, 
        n46286, n48861, n46447, n46404, n7_adj_4553, n48801, n46403, 
        n43090, n27288, n26950, n42888, n44677, n38240, n26840, 
        n46272, n46271, n38239, n43323, n43401, n40261, n34624;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n48978, n48972, n48966, n48960, n48954, n48948, n48942, 
        n48945, n48936, n12_adj_4554, n42838, n28592, n10_adj_4555, 
        n11_adj_4556, n28593, n28594, n9_adj_4557, n46355, n46356, 
        n48939, n46431, n46430, n38238, n43045, n43343, Kp_23__N_1330, 
        n43511, n43225, n42867;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n18_adj_4558, n27050, n16_adj_4559, n46448, n46449, n28595, 
        n46443, n46442, n20_adj_4560, n26557, n43432, n41082, n43123, 
        n27189, n12_adj_4561, n38237, n26744, n43377, n44609, n40284, 
        n38236, n28596, n1510, n25928, n28597, n40393, n27041, 
        n41122, n43241, n43386, n43487;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n8_adj_4562, n27056, n28598, n43340;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n12_adj_4563, n43174, n28599, n38235, n43162, n40582, n8_adj_4565, 
        n44811, n43293, n14_adj_4566, n43468, n43453, n15_adj_4567, 
        n42949, n27103, n27174, n42878, n43508, n43039, n10_adj_4568, 
        n42984, n6_adj_4569, n40326, n44005, n26676, n43417, n4_adj_4570, 
        n41149, n43484, n43398, n38234, n38233, n40244, n15_adj_4571, 
        n27234, n14_adj_4572, n43257, n46382, n26860, n42864, n26083, 
        n46383, n46389, n38232, n46388, n43183, n6_adj_4573, n41182, 
        n10_adj_4574, n27145, n26735, n43035, n6_adj_4575, n43474, 
        n1168, n43145, n48849, n48924, n48807, n7_adj_4576, n48918, 
        n47663, n48912, n48825, n7_adj_4577, n27053, n41096, n18_adj_4578, 
        n43334, n41094, n19_adj_4579, n43171, n43281, n42891, n26637, 
        n10_adj_4580, n43120, n46327, n46325, n42907, n6_adj_4581, 
        n6_adj_4582, n17_adj_4583, n41169, n38231, n42963, n43099, 
        n42915, n24, n43505, n43011, n40197, n22, n43374, n18_adj_4584, 
        n42928, n26, n43177, n43102, Kp_23__N_936, n40225, n47248, 
        Kp_23__N_1096, n27377, n46320, Kp_23__N_1099, Kp_23__N_1195, 
        n43523, n46321, n43496, n10_adj_4585, n48873, n48906, n46319, 
        n42957, n42955, n40294, n44813, n26504, n44105, n47247, 
        n9_adj_4586, n42925, n10_adj_4587, n9_adj_4588, n8_adj_4589, 
        n8_adj_4590, n28583, n46361, n46362, n28584, n28585, n43202, 
        n28147, n46368, n46367, n42222, n28586, n42220, n34718, 
        n28587, n38230, n28589, n75, n28590, n28591, n7_adj_4591, 
        n42218, n48819, n7_adj_4592, n10_adj_4593, n42810, n28535, 
        n28543, n28679, n28678, n28677, n28676, n28675, n42975, 
        n8_adj_4594, n28674, n28673, n28672, n28671, n28670, n28669, 
        n28668, n28667, n28666, n28665, n28664, n28663, n28660, 
        n28659, n28658, n28657, n28656, n28655, n28654, n28653, 
        n38229, n43077, n26656, n43459, n16_adj_4595, n28652, n43299, 
        n27425, n43049, n17_adj_4596, n46349, n46350, n48900, n43526, 
        n42216, n41242, n26843, n43429, n28546, n28578, n46347, 
        n46346, n47638, n28579, n28651, n28650, n43471, n43328, 
        n15_adj_4597, n28580, n28649, n43222, n40336, n41098, n42292, 
        n14_adj_4598, n27262, n28581, n28582, n43284, n12_adj_4599, 
        n48894, n28648, n43447, n47640, n28647, n28646, n48888, 
        n28645, n48813, n7_adj_4600, n28644, n28643, n41230, n43065, 
        n48882, n28642, n48855, n7_adj_4601, n28641, n28640, n28639, 
        n48870, n43108, n10_adj_4602, n48864, n48858, n28628, n48852, 
        n28627, n28626, n28625, Kp_23__N_1306, n10_adj_4603, n16_adj_4604, 
        n48846, n28624, n40205, n43083, n11_adj_4605, n48834, n26717, 
        n42995, n43520, n24464, n27306, n12_adj_4606, n43142, n42938, 
        n28611, n25962, n43105, n43003, n43052, n28610, n28609, 
        n42298, n26702, n8_adj_4607, n43004, n6_adj_4608, n40675, 
        n41193, n27149, n4_adj_4609, n27047, n43480, n26755, n40699, 
        n42302, n14_adj_4610, n10_adj_4611, n43093, n28608, n43251, 
        n32, n28607, n28606, n43132, n31_adj_4612, n35, n43015, 
        n42987, n10_adj_4613, n43311, n43151, n34, n6_adj_4614, 
        n43021, n10_adj_4615, n39_adj_4616, n43318, n44_adj_4617, 
        n38, n42268, n42168, n43502, n33, n32_adj_4618, n43008, 
        n44_adj_4619, n42969, n42_adj_4620, n27296, n43314, n43_adj_4621, 
        n43031, n43371, n42_adj_4622, n43456, n43517, n43_adj_4623, 
        n28604, n43165, n41_adj_4624, n43308, n43490, n40_adj_4625, 
        n50_adj_4626, n45_adj_4627, n43356, n41_adj_4628, n38228, 
        n41117, n40922, n44527, n43444, n43158, n40_adj_4629, n26915, 
        n39_adj_4630, n10_adj_4631, n50_adj_4632, n43296, n6_adj_4633, 
        n38227, n38226, n43359, n34442, n26456, n45_adj_4636, n28603, 
        n27421, n28602, n43287, n14_adj_4637, n9_adj_4638, n42932, 
        n41143, n41113, n41184, n26747, n6_adj_4639, n6_adj_4640;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n5_adj_4641, n42921, n38225, Kp_23__N_1189, n13, n18_adj_4642, 
        n1247, n27360, n16_adj_4643, n27403, n38224, n27078, n42966, 
        n43071, n17_adj_4644, n7_adj_4645, n26593, n26599, n27072, 
        n38223, n26604, n42960, n27253, n26545, n1513, n42881, 
        n26580, n27500, n27059, n26905, n43426, n27258, n10_adj_4646, 
        n4_adj_4647, n27062, n26730, n24669, n6_adj_4648, n8_adj_4649, 
        n10_adj_4650, Kp_23__N_1186, n26624, n38222, n8_adj_4651, 
        n8_adj_4652, n28525, n27152, n28526, n28527, n28528, n38221, 
        n43245, n16_adj_4653, n43238, n17_adj_4654, n28530, n28531, 
        n38220, n43465, n43392, n43331, n26662, n43028, n14_adj_4655, 
        n4_adj_4656, n41086, n44882, n28532, n28533, n43193, n38219, 
        n42816, n38218, n27139, n10_adj_4657, n48828, n44237, Kp_23__N_1093, 
        Kp_23__N_1090, n14_adj_4658, n48822, n12_adj_4659, n27186, 
        n41188, n38217, n11_adj_4660, n26050, n6_adj_4661, n42991, 
        n38216, n48816, n48810, n38215, n48804, n48798, n38214, 
        n26863, n43042, n43148, n27354, n40238, n28601, n43114, 
        n43126, n8_adj_4662, n28517, n28518, n28519, n7_adj_4663, 
        n28520, n28521, n28522, n7_adj_4664, n42190, n42312, n42204, 
        n33802, n42206, n42310, n42208, n42308, n42210, n42248, 
        n34417, n42306, n42212, n7_adj_4665, n8_adj_4666, n39601, 
        n42164, n42244, n34415, n7_adj_4667, n34413, n42304, n42214, 
        n7_adj_4668, n34411, n42286, n42224, n42284, n42226, n7_adj_4669, 
        n8_adj_4670, n42282, n42182, n42228, n42276, n42230, n42274, 
        n34409, n42272, n42232, n42270, n42176, n42178, n27469, 
        n42918, n12_adj_4671, n28523, n28524, n44659, n5_adj_4672, 
        n14_adj_4673, Kp_23__N_1301, n10_adj_4674, n28600, n38213, 
        n38212, n38211, n38210, n38209, n42896, n20_adj_4675, n19_adj_4676, 
        n21, n42912, n28501, n28502, n38208, n38207, n28503, n28504, 
        n28505, n28506, n28507, n28508, n38206, n42902, n38205, 
        n38204, n43055, n10_adj_4677, n43347, n8_adj_4678, n28493, 
        n28494, n28495, n28496, n28497, n28498, n28499, n28500, 
        n42832, n28485, n28486, n28487, n28488, n28489, n28490, 
        n28491, n14_adj_4679, n28492, n28477, n28478, n28479, n28480, 
        n28481, n42952, n28482, n28483, n28484, n28469, n28470, 
        n28471, n28472, n28473, n28474, n28475, n28476, n28461, 
        n28462, n28463, n28464, n28465, n28468, n28467, n28466, 
        n28460, n28459, n28458, n28457, n28456, n28455, n28454, 
        n28453, n28, n43275, n42884, n42899, n32_adj_4680, n43272, 
        n30, n31_adj_4681, n41090, n27357, n29, n26667, n2_adj_4682, 
        n43111, n6_adj_4683, n24_adj_4684, n22_adj_4685, n26_adj_4686, 
        n42981, n12_adj_4687, n44479, n41145, n16_adj_4688, n17_adj_4689, 
        n45310, n12_adj_4690, n8_adj_4691, n44982, n44432, n1130, 
        n44899, n45108, n10_adj_4692, n44441, n44205, n44203, n34626, 
        n44641, n49063, n12_adj_4693, n44064, n8_adj_4694, n44594, 
        n20_adj_4695, n18_adj_4696, n19_adj_4697, n17_adj_4698, n6_adj_4699, 
        n22_adj_4700, n28_adj_4701, n21_adj_4702, n29_adj_4703, n43180, 
        n6_adj_4704, n12_adj_4705, n46303, n24_adj_4706, n24791, n46282, 
        n26_adj_4707, n43235, n26491, n29_adj_4708, n46147, n12_adj_4709, 
        n28_adj_4710, n43414, n6_adj_4711, n32_adj_4712, n44251, n46149, 
        n12_adj_4713, n8_adj_4714, n12_adj_4715, n48, n48780, n43006, 
        n56, n55, n63_adj_4716, n34434;
    
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n28234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n28233));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33_4_lut (.I0(n57), .I1(n59), .I2(n58), .I3(n60), .O(n69));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35_4_lut (.I0(n69), .I1(n61), .I2(n68), .I3(n62), .O(n26879));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n28232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n28231));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n28230));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_658_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n28229));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n28228));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n28227));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2), .S(n3_adj_4435));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4436), .S(n3_adj_4437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n28226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n28225));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4438));
    defparam select_658_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31233_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46314));
    defparam i31233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31234_4_lut (.I0(n46314), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n46315));
    defparam i31234_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i31232_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46313));
    defparam i31232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33689_3_lut (.I0(n141), .I1(n43606), .I2(n34377), .I3(GND_net), 
            .O(n45195));
    defparam i33689_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_4_lut (.I0(n7001), .I1(\FRAME_MATCHER.state [1]), .I2(n23743), 
            .I3(n3_adj_4439), .O(n4_c));
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 i1_4_lut_adj_884 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n4_c), .I3(\FRAME_MATCHER.state_31__N_2724 [3]), .O(n16));
    defparam i1_4_lut_adj_884.LUT_INIT = 16'ha0e4;
    SB_LUT4 i33322_4_lut (.I0(n16), .I1(n4_adj_4440), .I2(\FRAME_MATCHER.state [0]), 
            .I3(n34628), .O(n44876));
    defparam i33322_4_lut.LUT_INIT = 16'h3133;
    SB_LUT4 i32201_2_lut (.I0(n48951), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47240));
    defparam i32201_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31227_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46308));
    defparam i31227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31228_4_lut (.I0(n46308), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n46309));
    defparam i31228_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i31226_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46307));
    defparam i31226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32249_2_lut (.I0(n48957), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47249));
    defparam i32249_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31310_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46391));
    defparam i31310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31311_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46392));
    defparam i31311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31251_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46332));
    defparam i31251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31250_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21][4] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46331));
    defparam i31250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31200_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46281));
    defparam i31200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31199_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46280));
    defparam i31199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32188_2_lut (.I0(n48981), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47236));
    defparam i32188_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut (.I0(n40416), .I1(n40271), .I2(n42861), .I3(n6), 
            .O(n44663));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_885 (.I0(n40271), .I1(\data_out_frame[25] [7]), 
            .I2(n41102), .I3(n6_adj_4441), .O(n45100));
    defparam i4_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_886 (.I0(n40416), .I1(\data_out_frame[23] [6]), 
            .I2(n43263), .I3(n6_adj_4442), .O(n44071));
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut (.I0(n27326), .I1(n43290), .I2(n41232), .I3(\data_out_frame[15] [2]), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[19] [4]), .I1(n12), .I2(n43450), 
            .I3(\data_out_frame[19] [3]), .O(n40416));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43263));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_887 (.I0(n40416), .I1(\data_out_frame[23] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41102));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n41102), .I1(n43435), .I2(n43263), .I3(n42871), 
            .O(n44066));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_888 (.I0(n43168), .I1(n27031), .I2(n27010), .I3(n43395), 
            .O(n10));
    defparam i4_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[19] [5]), .I1(n10), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n2134));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_889 (.I0(\data_out_frame[24] [2]), .I1(n2134), 
            .I2(GND_net), .I3(GND_net), .O(n43435));
    defparam i1_2_lut_adj_889.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_out_frame[22] [0]), .I1(n43154), 
            .I2(n40935), .I3(n44246), .O(n43438));
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_891 (.I0(n43197), .I1(n43438), .I2(n43435), .I3(n43266), 
            .O(n44073));
    defparam i3_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_out_frame[24] [3]), .I1(n41175), 
            .I2(GND_net), .I3(GND_net), .O(n43266));
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_893 (.I0(\data_out_frame[22] [3]), .I1(n40257), 
            .I2(n42871), .I3(n6_adj_4443), .O(n44687));
    defparam i4_4_lut_adj_893.LUT_INIT = 16'h9669;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_894 (.I0(n43368), .I1(n40257), .I2(n41175), .I3(n6_adj_4444), 
            .O(n45206));
    defparam i4_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_out_frame[20] [1]), .I1(n45042), 
            .I2(GND_net), .I3(GND_net), .O(n43368));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_896 (.I0(\data_out_frame[17] [5]), .I1(n27326), 
            .I2(n43190), .I3(n6_adj_4445), .O(n41175));
    defparam i4_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_897 (.I0(n43368), .I1(\data_out_frame[24] [6]), 
            .I2(n41236), .I3(\data_out_frame[24] [5]), .O(n14));
    defparam i6_4_lut_adj_897.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut (.I0(n41104), .I1(n14), .I2(n10_adj_4446), .I3(n40257), 
            .O(n44272));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_898 (.I0(n26879), .I1(n40830), .I2(GND_net), 
            .I3(GND_net), .O(n41104));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n28224));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_out_frame[15] [4]), .I1(n43514), 
            .I2(GND_net), .I3(GND_net), .O(n43190));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n27621), .D(n8825[1]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n27621), .D(n8825[2]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n27621), .D(n8825[3]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n27621), .D(n8825[4]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n27621), .D(n8825[5]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n27621), .D(n8825[6]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n27621), .D(n8825[7]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_900 (.I0(\data_out_frame[17] [6]), .I1(n27031), 
            .I2(n43190), .I3(n43407), .O(n45249));
    defparam i3_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n28223));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_adj_901 (.I0(n41137), .I1(\data_out_frame[24] [7]), 
            .I2(n45042), .I3(GND_net), .O(n14_adj_4447));
    defparam i5_3_lut_adj_901.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_902 (.I0(n43362), .I1(\data_out_frame[25] [0]), 
            .I2(n40257), .I3(n43074), .O(n15));
    defparam i6_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n41109), .I2(n14_adj_4447), .I3(n41208), 
            .O(n40830));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_903 (.I0(n43999), .I1(n40830), .I2(GND_net), 
            .I3(GND_net), .O(n27241));
    defparam i1_2_lut_adj_903.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_904 (.I0(\data_out_frame[20] [5]), .I1(n43199), 
            .I2(\data_out_frame[24] [7]), .I3(n41236), .O(n12_adj_4448));
    defparam i5_4_lut_adj_904.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_905 (.I0(\data_out_frame[18] [1]), .I1(n12_adj_4448), 
            .I2(n43411), .I3(\data_out_frame[20] [3]), .O(n43999));
    defparam i6_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[25] [2]), .I1(n40829), .I2(n43999), 
            .I3(GND_net), .O(n44713));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_906 (.I0(n40210), .I1(\data_out_frame[25] [3]), 
            .I2(n40307), .I3(GND_net), .O(n44637));
    defparam i2_3_lut_adj_906.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_907 (.I0(n41135), .I1(n41204), .I2(\data_out_frame[23] [2]), 
            .I3(n6_adj_4449), .O(n40307));
    defparam i4_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n40307), .I1(n44012), .I2(GND_net), 
            .I3(GND_net), .O(n26801));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_909 (.I0(\data_out_frame[10] [4]), .I1(n43462), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n14_adj_4450));   // verilog/coms.v(73[16:42])
    defparam i5_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_910 (.I0(n130), .I1(n3_adj_4439), .I2(n110), 
            .I3(GND_net), .O(n27595));
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h0202;
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4451), .S(n3_adj_4438));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_911 (.I0(\data_out_frame[6] [2]), .I1(n43305), 
            .I2(\data_out_frame[14] [6]), .I3(n1516), .O(n15_adj_4452));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_912 (.I0(n15_adj_4452), .I1(\data_out_frame[12] [5]), 
            .I2(n14_adj_4450), .I3(\data_out_frame[12] [4]), .O(n27010));   // verilog/coms.v(73[16:42])
    defparam i8_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4453));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_913 (.I0(n43209), .I1(\data_out_frame[16] [6]), 
            .I2(n27010), .I3(\data_out_frame[17] [0]), .O(n14_adj_4454));
    defparam i6_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_914 (.I0(\data_out_frame[21][2] ), .I1(n14_adj_4454), 
            .I2(n10_adj_4453), .I3(\data_out_frame[19] [0]), .O(n41135));
    defparam i7_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_915 (.I0(\data_out_frame[17] [2]), .I1(n43187), 
            .I2(n27484), .I3(n40355), .O(n41177));
    defparam i3_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_916 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(n43206), .I3(n42944), .O(n41232));
    defparam i3_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_917 (.I0(n43278), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(n43441), .O(n10_adj_4455));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_918 (.I0(n43216), .I1(n41137), .I2(n40271), .I3(n43420), 
            .O(n10_adj_4456));
    defparam i4_4_lut_adj_918.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_919 (.I0(\data_out_frame[23] [3]), .I1(n10_adj_4456), 
            .I2(n40347), .I3(GND_net), .O(n44012));
    defparam i5_3_lut_adj_919.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_920 (.I0(n41177), .I1(n41135), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n43254));
    defparam i2_3_lut_adj_920.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n1), .I2(n42849), 
            .I3(GND_net), .O(n81));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_4_lut_adj_921 (.I0(\FRAME_MATCHER.state_31__N_2724 [3]), .I1(n81), 
            .I2(n8), .I3(n43600), .O(n10_adj_4457));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_921.LUT_INIT = 16'hccec;
    SB_LUT4 i2_4_lut (.I0(\FRAME_MATCHER.state_c [8]), .I1(n21657), .I2(n1), 
            .I3(n9), .O(n7_c));
    defparam i2_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i33683_2_lut (.I0(n34544), .I1(n19789), .I2(GND_net), .I3(GND_net), 
            .O(tx_transmit_N_3513));
    defparam i33683_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i16348_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n29859));   // verilog/coms.v(112[11:16])
    defparam i16348_3_lut.LUT_INIT = 16'hc9c9;
    SB_LUT4 i2_4_lut_adj_922 (.I0(n26449), .I1(n29859), .I2(n3065), .I3(n11), 
            .O(n3813));
    defparam i2_4_lut_adj_922.LUT_INIT = 16'h0a08;
    SB_LUT4 i20491_4_lut (.I0(n8_adj_4458), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26350), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i20491_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_4_lut_adj_923 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n23534), 
            .I2(n1), .I3(n9), .O(n7_adj_4459));
    defparam i2_4_lut_adj_923.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\FRAME_MATCHER.state [1]), .I1(n29908), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2626 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h8888;
    SB_LUT4 i20487_4_lut (.I0(n5_c), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i20487_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\FRAME_MATCHER.state [1]), .I1(n29908), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2620 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h4444;
    SB_LUT4 i5_3_lut_adj_926 (.I0(\data_in[0] [3]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4460));
    defparam i5_3_lut_adj_926.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_927 (.I0(\data_in[0] [6]), .I1(n26425), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4461));
    defparam i6_4_lut_adj_927.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_928 (.I0(n15_adj_4461), .I1(\data_in[3] [0]), .I2(n14_adj_4460), 
            .I3(\data_in[2] [2]), .O(n26245));
    defparam i8_4_lut_adj_928.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_929 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4462));
    defparam i6_4_lut_adj_929.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_930 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_930.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in[1] [6]), .I2(n16_adj_4462), 
            .I3(\data_in[3] [7]), .O(n26347));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_931 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4463));
    defparam i4_4_lut_adj_931.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_932 (.I0(\data_in[3] [4]), .I1(n10_adj_4463), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n26425));
    defparam i5_3_lut_adj_932.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut_adj_933 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4464));
    defparam i2_2_lut_adj_933.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_934 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4465));
    defparam i6_4_lut_adj_934.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_935 (.I0(\data_in[3] [6]), .I1(n14_adj_4465), .I2(n10_adj_4464), 
            .I3(\data_in[2] [1]), .O(n26422));
    defparam i7_4_lut_adj_935.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_936 (.I0(\data_in[2] [4]), .I1(n26422), .I2(\data_in[1] [5]), 
            .I3(n26425), .O(n18));
    defparam i7_4_lut_adj_936.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_937 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n26347), .O(n20));
    defparam i9_4_lut_adj_937.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4466));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4466), .I1(n20), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_c));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_938 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n26245), .O(n16_adj_4467));
    defparam i6_4_lut_adj_938.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_939 (.I0(n26347), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_4468));
    defparam i7_4_lut_adj_939.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_940 (.I0(n17_adj_4468), .I1(\data_in[3] [5]), .I2(n16_adj_4467), 
            .I3(\data_in[3] [1]), .O(n63_adj_4469));
    defparam i9_4_lut_adj_940.LUT_INIT = 16'hfbff;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n28222));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_941 (.I0(n2_adj_4470), .I1(\FRAME_MATCHER.i_31__N_2620 ), 
            .I2(n771), .I3(n23534), .O(n42849));
    defparam i1_4_lut_adj_941.LUT_INIT = 16'haeaa;
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n28221));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n26350));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_942 (.I0(\FRAME_MATCHER.i [4]), .I1(n26350), .I2(GND_net), 
            .I3(GND_net), .O(n26232));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_942.LUT_INIT = 16'heeee;
    SB_LUT4 i20490_4_lut (.I0(n8_adj_4471), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26232), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i20490_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i8_4_lut_adj_943 (.I0(n26422), .I1(\data_in[1] [3]), .I2(n26245), 
            .I3(\data_in[1] [2]), .O(n20_adj_4472));
    defparam i8_4_lut_adj_943.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_944 (.I0(n21657), .I1(n3813), .I2(GND_net), .I3(GND_net), 
            .O(n1_adj_4473));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_945 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_945.LUT_INIT = 16'hfeff;
    SB_LUT4 i31184_4_lut (.I0(\data_in[3] [2]), .I1(\data_in[0] [5]), .I2(\data_in[2] [0]), 
            .I3(\data_in[2] [5]), .O(n46207));
    defparam i31184_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n46207), .I1(n19), .I2(n20_adj_4472), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 select_686_Select_1_i5_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2624 ), 
            .I2(n3303), .I3(n92[1]), .O(n5_adj_4475));
    defparam select_686_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n1_adj_4473), 
            .I2(n46187), .I3(n2_adj_4470), .O(n42122));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_3_lut_adj_947 (.I0(n92[1]), .I1(n9), .I2(n63), .I3(GND_net), 
            .O(n39751));
    defparam i1_3_lut_adj_947.LUT_INIT = 16'h8c8c;
    SB_LUT4 i3_4_lut_adj_948 (.I0(\FRAME_MATCHER.i_31__N_2622 ), .I1(n39751), 
            .I2(n1_adj_4476), .I3(n5_adj_4475), .O(n48985));
    defparam i3_4_lut_adj_948.LUT_INIT = 16'hfffe;
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4477), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31370_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46451));
    defparam i31370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31371_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46452));
    defparam i31371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31260_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46341));
    defparam i31260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31259_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46340));
    defparam i31259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31262_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46343));
    defparam i31262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31263_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46344));
    defparam i31263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31353_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46434));
    defparam i31353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31352_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46433));
    defparam i31352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4478));
    defparam select_658_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31271_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46352));
    defparam i31271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4479));
    defparam select_658_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31272_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46353));
    defparam i31272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4480));
    defparam select_658_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31347_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46428));
    defparam i31347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31346_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46427));
    defparam i31346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31298_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46379));
    defparam i31298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4481));
    defparam select_658_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31299_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46380));
    defparam i31299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31329_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46410));
    defparam i31329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31328_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46409));
    defparam i31328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4482));
    defparam select_658_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31304_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46385));
    defparam i31304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31305_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46386));
    defparam i31305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31293_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46374));
    defparam i31293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31292_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46373));
    defparam i31292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31313_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46394));
    defparam i31313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31314_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46395));
    defparam i31314_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4483), .S(n3_adj_4484));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4485), .S(n3_adj_4486));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2_adj_4487), .S(n3_adj_4488));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4489), .S(n3_adj_4490));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31215_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46296));
    defparam i31215_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4491), .S(n3_adj_4492));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31214_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46295));
    defparam i31214_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4493), .S(n3_adj_4494));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4495), .S(n3_adj_4496));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4497), .S(n3_adj_4498));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4499), .S(n3_adj_4500));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3616[0]), .C(CLK_c), .D(n4888[0]), 
            .R(n43770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4501), .S(n3_adj_4502));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4503), .S(n3_adj_4504));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n27605), .D(n7002));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4505), .S(n3_adj_4506));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4507), .S(n3_adj_4508));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4509), .S(n3_adj_4510));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4511), .S(n3_adj_4512));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4513), .S(n3_adj_4514));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4515), .S(n3_adj_4516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n28220));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4517), .S(n3_adj_4518));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4519), .S(n3_adj_4520));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_949 (.I0(\FRAME_MATCHER.state_c [29]), .I1(\FRAME_MATCHER.state_c [30]), 
            .I2(\FRAME_MATCHER.state_c [13]), .I3(\FRAME_MATCHER.state_c [21]), 
            .O(n10_adj_4521));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_949.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n28219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n28218));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4522), .S(n3_adj_4523));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4524), .S(n3_adj_4525));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4526), .S(n3_adj_4527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n28217));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31316_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46397));
    defparam i31316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31317_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46398));
    defparam i31317_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4528), .S(n3_adj_4529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n28216));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n28215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n28214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n28213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n28212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n28211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n28210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n28209));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4530), .S(n3_adj_4482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n28208));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4531), .S(n3_adj_4481));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_950 (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(n3303), 
            .I2(n23534), .I3(GND_net), .O(n2_adj_4470));   // verilog/coms.v(115[11:12])
    defparam i1_3_lut_adj_950.LUT_INIT = 16'h2020;
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n28207));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_951 (.I0(n63_c), .I1(n63), .I2(n63_adj_4469), 
            .I3(GND_net), .O(n21657));   // verilog/coms.v(157[6] 159[9])
    defparam i2_3_lut_adj_951.LUT_INIT = 16'h8080;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4532), .S(n3_adj_4480));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4533), .S(n3_adj_4479));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_952 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n12_adj_4534), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(\FRAME_MATCHER.state_c [11]), 
            .O(n42707));   // verilog/coms.v(127[12] 300[6])
    defparam i6_4_lut_adj_952.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_953 (.I0(n42707), .I1(\FRAME_MATCHER.state_c [14]), 
            .I2(n10_adj_4521), .I3(\FRAME_MATCHER.state_c [19]), .O(n4_adj_4535));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_954 (.I0(\FRAME_MATCHER.state_c [7]), .I1(\FRAME_MATCHER.state_c [5]), 
            .I2(\FRAME_MATCHER.state_c [6]), .I3(GND_net), .O(n42854));
    defparam i2_3_lut_adj_954.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n133));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h2222;
    SB_LUT4 select_658_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4529));
    defparam select_658_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_956 (.I0(n110), .I1(n31), .I2(n133), .I3(\FRAME_MATCHER.state [2]), 
            .O(n27596));
    defparam i3_4_lut_adj_956.LUT_INIT = 16'h1000;
    SB_LUT4 i4_4_lut_adj_957 (.I0(\data_out_frame[18] [7]), .I1(n43499), 
            .I2(\data_out_frame[16] [0]), .I3(n44262), .O(n10_adj_4536));
    defparam i4_4_lut_adj_957.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4537), .S(n3_adj_4478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n28206));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4527));
    defparam select_658_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[5] [5]), 
            .I2(n43350), .I3(\data_in_frame[7] [6]), .O(n43117));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n28205));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_958 (.I0(\data_out_frame[21][1] ), .I1(\data_out_frame[19] [0]), 
            .I2(n8_adj_4538), .I3(n43269), .O(n43420));
    defparam i1_4_lut_adj_958.LUT_INIT = 16'h9669;
    SB_LUT4 mux_2022_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7003));
    defparam mux_2022_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_959 (.I0(\data_out_frame[18] [3]), .I1(n41115), 
            .I2(\data_out_frame[20] [5]), .I3(GND_net), .O(n43362));
    defparam i2_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 mux_2022_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7004));
    defparam mux_2022_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7005));
    defparam mux_2022_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43411));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2022_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7006));
    defparam mux_2022_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n28204));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_2022_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7007));
    defparam mux_2022_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7008));
    defparam mux_2022_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7009));
    defparam mux_2022_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7010));
    defparam mux_2022_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7011));
    defparam mux_2022_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7012));
    defparam mux_2022_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7013));
    defparam mux_2022_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_961 (.I0(n43362), .I1(\data_out_frame[22] [7]), 
            .I2(\data_out_frame[23] [2]), .I3(n43420), .O(n10_adj_4539));
    defparam i4_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7014));
    defparam mux_2022_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7015));
    defparam mux_2022_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7016));
    defparam mux_2022_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n28203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n28202));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_2022_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7017));
    defparam mux_2022_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_962 (.I0(\data_out_frame[21][0] ), .I1(n43080), 
            .I2(n43353), .I3(n6_adj_4540), .O(n40829));
    defparam i4_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7018));
    defparam mux_2022_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
            .D(n42174), .S(n48985));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_2022_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7019));
    defparam mux_2022_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7020));
    defparam mux_2022_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7021));
    defparam mux_2022_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_969), 
            .I2(GND_net), .I3(GND_net), .O(n42941));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42861));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2022_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7022));
    defparam mux_2022_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7023));
    defparam mux_2022_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_965 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43068));
    defparam i1_2_lut_adj_965.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2022_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7024));
    defparam mux_2022_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7025));
    defparam mux_2022_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_966 (.I0(\data_out_frame[25] [3]), .I1(n40829), 
            .I2(\data_out_frame[25] [2]), .I3(n40210), .O(n43088));
    defparam i3_4_lut_adj_966.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_967 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[21][4] ), .I3(n27122), .O(n12_adj_4541));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_968 (.I0(\data_out_frame[17] [0]), .I1(n12_adj_4541), 
            .I2(\data_out_frame[19] [2]), .I3(\data_out_frame[19] [3]), 
            .O(n43187));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43248));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43365));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_971 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [4]), .I3(GND_net), .O(n43080));
    defparam i2_3_lut_adj_971.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\data_out_frame[15] [1]), .I1(n25950), 
            .I2(GND_net), .I3(GND_net), .O(n40355));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4525));
    defparam select_658_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4523));
    defparam select_658_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_973 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n44678));
    defparam i2_3_lut_adj_973.LUT_INIT = 16'h8080;
    SB_LUT4 i5_3_lut_adj_974 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[20] [1]), 
            .I2(n43383), .I3(GND_net), .O(n14_adj_4542));
    defparam i5_3_lut_adj_974.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_975 (.I0(n43493), .I1(\data_out_frame[17] [5]), 
            .I2(n42944), .I3(n43450), .O(n15_adj_4543));
    defparam i6_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_976 (.I0(n15_adj_4543), .I1(n43154), .I2(n14_adj_4542), 
            .I3(\data_out_frame[19] [5]), .O(n44246));
    defparam i8_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_977 (.I0(n27090), .I1(\data_out_frame[22] [1]), 
            .I2(n44246), .I3(GND_net), .O(n42871));
    defparam i2_3_lut_adj_977.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_978 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[24] [6]), 
            .I2(\data_out_frame[22] [7]), .I3(GND_net), .O(n43074));
    defparam i2_3_lut_adj_978.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43168));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_980 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43216));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[21][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n43278));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_982 (.I0(n26855), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(\data_out_frame[17] [4]), 
            .O(n43383));
    defparam i3_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_983 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n4_adj_4544), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/coms.v(151[5:27])
    defparam i2_2_lut_adj_983.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_out_frame[13] [0]), .I1(n42978), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4545));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i31221_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46302));
    defparam i31221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32244_2_lut (.I0(n48963), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47254));
    defparam i32244_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31194_4_lut (.I0(byte_transmit_counter[0]), .I1(n47254), .I2(byte_transmit_counter[3]), 
            .I3(\data_out_frame[20] [5]), .O(n46275));
    defparam i31194_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i20_3_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\data_out_frame[23] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4546));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_985 (.I0(n43383), .I1(n25950), .I2(\data_out_frame[19] [6]), 
            .I3(n6_adj_4545), .O(n40935));
    defparam i4_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n27621), .D(n8825[0]), .R(n28080));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_out_frame[20] [0]), .I1(n40935), 
            .I2(GND_net), .I3(GND_net), .O(n43196));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i31220_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46301));
    defparam i31220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31332_4_lut (.I0(n48783), .I1(n46276), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n46413));
    defparam i31332_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 select_658_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4520));
    defparam select_658_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31331_3_lut (.I0(n7_adj_4547), .I1(n48831), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n46412));
    defparam i31331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31333_3_lut (.I0(n46412), .I1(n46413), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[5]));
    defparam i31333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32241_2_lut (.I0(n48969), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47227));
    defparam i32241_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31374_4_lut (.I0(byte_transmit_counter[0]), .I1(n47227), .I2(byte_transmit_counter[3]), 
            .I3(\data_out_frame[20] [6]), .O(n46455));
    defparam i31374_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i20_3_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\data_out_frame[23] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4548));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_987 (.I0(n26832), .I1(n27522), .I2(\data_out_frame[14] [7]), 
            .I3(GND_net), .O(n42944));
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h9696;
    SB_LUT4 i20302_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), .I2(GND_net), 
            .I3(GND_net), .O(n33792));
    defparam i20302_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i31213_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n46294));
    defparam i31213_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31211_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46292));
    defparam i31211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31326_4_lut (.I0(n48867), .I1(n46456), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n46407));
    defparam i31326_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31325_3_lut (.I0(n7_adj_4549), .I1(n48837), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n46406));
    defparam i31325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31327_3_lut (.I0(n46406), .I1(n46407), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[6]));
    defparam i31327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_988 (.I0(n43423), .I1(n1191), .I2(\data_out_frame[12] [6]), 
            .I3(n43302), .O(n15_adj_4550));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4518));
    defparam select_658_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut_adj_989 (.I0(n15_adj_4550), .I1(\data_out_frame[4] [1]), 
            .I2(n14_adj_4551), .I3(\data_out_frame[10] [4]), .O(n25950));   // verilog/coms.v(75[16:43])
    defparam i8_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n38241), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n28200));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i32239_2_lut (.I0(n48975), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47229));
    defparam i32239_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_658_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4516));
    defparam select_658_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31365_4_lut (.I0(byte_transmit_counter[0]), .I1(n47229), .I2(byte_transmit_counter[3]), 
            .I3(\data_out_frame[20] [7]), .O(n46446));
    defparam i31365_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42858));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i20_3_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\data_out_frame[23] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4552));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_991 (.I0(n44678), .I1(n36539), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n26449));   // verilog/coms.v(212[5:16])
    defparam i2_3_lut_adj_991.LUT_INIT = 16'hfdfd;
    SB_LUT4 i31207_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n46288));
    defparam i31207_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31205_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46286));
    defparam i31205_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n28199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n28198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n28197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n28196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n28195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n28194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n28193));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31323_4_lut (.I0(n48861), .I1(n46447), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n46404));
    defparam i31323_4_lut.LUT_INIT = 16'hccca;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n28192));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31322_3_lut (.I0(n7_adj_4553), .I1(n48801), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n46403));
    defparam i31322_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n28191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n28190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n28189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n28188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n28187));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n28186));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_992 (.I0(n43197), .I1(\data_out_frame[24] [5]), 
            .I2(\data_out_frame[24] [4]), .I3(GND_net), .O(n43090));
    defparam i2_3_lut_adj_992.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_993 (.I0(n25950), .I1(n42944), .I2(GND_net), 
            .I3(GND_net), .O(n43290));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i31324_3_lut (.I0(n46403), .I1(n46404), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[7]));
    defparam i31324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14574_2_lut (.I0(\FRAME_MATCHER.i_31__N_2622 ), .I1(n26449), 
            .I2(GND_net), .I3(GND_net), .O(n28080));   // verilog/coms.v(127[12] 300[6])
    defparam i14574_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n28185));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_994 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[12] [1]), 
            .I2(n27288), .I3(\data_out_frame[12] [2]), .O(n26950));
    defparam i3_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n28184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n28183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n28182));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4514));
    defparam select_658_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_out_frame[16] [4]), .I1(n26950), 
            .I2(GND_net), .I3(GND_net), .O(n42888));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4512));
    defparam select_658_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4510));
    defparam select_658_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4437));
    defparam select_658_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_996 (.I0(\data_out_frame[18] [5]), .I1(n42888), 
            .I2(n44677), .I3(\data_out_frame[16] [3]), .O(n40347));
    defparam i3_4_lut_adj_996.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n28181));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_997 (.I0(n41204), .I1(n40347), .I2(GND_net), 
            .I3(GND_net), .O(n41109));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h9999;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n38240), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n28180));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_998 (.I0(n26840), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n43269));
    defparam i2_3_lut_adj_998.LUT_INIT = 16'h9696;
    SB_LUT4 i31191_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46272));
    defparam i31191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33680_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n141));
    defparam i33680_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\FRAME_MATCHER.state [0]), .I1(n36539), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_999.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1000 (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(n29908), 
            .I2(GND_net), .I3(GND_net), .O(n3065));
    defparam i2_2_lut_adj_1000.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(n3065), .I1(n11), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n141), .O(n3846));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'h5455;
    SB_LUT4 i31190_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46271));
    defparam i31190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4435));
    defparam select_658_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4508));
    defparam select_658_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1002 (.I0(n27484), .I1(n43209), .I2(\data_out_frame[20] [7]), 
            .I3(GND_net), .O(n41137));
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_8 (.CI(n38240), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n38241));
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n38239), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1003 (.I0(n43323), .I1(n43401), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n40261));
    defparam i2_3_lut_adj_1003.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n34377), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n4_adj_4440));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i21115_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n34377), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n34624));
    defparam i21115_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n48978));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48978_bdd_4_lut (.I0(n48978), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48981));
    defparam n48978_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33861 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48972));
    defparam byte_transmit_counter_0__bdd_4_lut_33861.LUT_INIT = 16'he4aa;
    SB_LUT4 n48972_bdd_4_lut (.I0(n48972), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48975));
    defparam n48972_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33856 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48966));
    defparam byte_transmit_counter_0__bdd_4_lut_33856.LUT_INIT = 16'he4aa;
    SB_LUT4 n48966_bdd_4_lut (.I0(n48966), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48969));
    defparam n48966_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33851 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48960));
    defparam byte_transmit_counter_0__bdd_4_lut_33851.LUT_INIT = 16'he4aa;
    SB_LUT4 n48960_bdd_4_lut (.I0(n48960), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48963));
    defparam n48960_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33846 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48954));
    defparam byte_transmit_counter_0__bdd_4_lut_33846.LUT_INIT = 16'he4aa;
    SB_LUT4 n48954_bdd_4_lut (.I0(n48954), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48957));
    defparam n48954_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33841 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48948));
    defparam byte_transmit_counter_0__bdd_4_lut_33841.LUT_INIT = 16'he4aa;
    SB_LUT4 n48948_bdd_4_lut (.I0(n48948), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48951));
    defparam n48948_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33836 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48942));
    defparam byte_transmit_counter_0__bdd_4_lut_33836.LUT_INIT = 16'he4aa;
    SB_LUT4 n48942_bdd_4_lut (.I0(n48942), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48945));
    defparam n48942_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33831 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27][1] ), 
            .I3(byte_transmit_counter[1]), .O(n48936));
    defparam byte_transmit_counter_0__bdd_4_lut_33831.LUT_INIT = 16'he4aa;
    SB_LUT4 select_658_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4506));
    defparam select_658_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28587_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43606));
    defparam i28587_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1004 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4554));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1004.LUT_INIT = 16'h7bde;
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n28179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n28178));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15081_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n28592));
    defparam i15081_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1005 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4555));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1005.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1006 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4556));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1006.LUT_INIT = 16'h7bde;
    SB_CARRY add_3971_7 (.CI(n38239), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n38240));
    SB_LUT4 i15082_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n28593));
    defparam i15082_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15083_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n28594));
    defparam i15083_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_4557));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'h7bde;
    SB_LUT4 i31274_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46355));
    defparam i31274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31275_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46356));
    defparam i31275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n48936_bdd_4_lut (.I0(n48936), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n48939));
    defparam n48936_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i31350_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46431));
    defparam i31350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31349_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21][0] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46430));
    defparam i31349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1008 (.I0(n9_adj_4557), .I1(n11_adj_4556), .I2(n10_adj_4555), 
            .I3(n12_adj_4554), .O(n23743));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1008.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n38238), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(n43045), .I1(n43343), .I2(Kp_23__N_1330), 
            .I3(GND_net), .O(n43511));
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1010 (.I0(\data_in_frame[18] [0]), .I1(n43225), 
            .I2(n42867), .I3(\data_in_frame[15] [6]), .O(n18_adj_4558));   // verilog/coms.v(73[16:42])
    defparam i7_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(\data_in_frame[11] [4]), .I1(n27050), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4559));   // verilog/coms.v(73[16:42])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31367_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46448));
    defparam i31367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31368_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46449));
    defparam i31368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15084_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n28595));
    defparam i15084_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31362_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46443));
    defparam i31362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31361_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46442));
    defparam i31361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1011 (.I0(\data_in_frame[11] [3]), .I1(n18_adj_4558), 
            .I2(Kp_23__N_1330), .I3(\data_in_frame[13] [4]), .O(n20_adj_4560));   // verilog/coms.v(73[16:42])
    defparam i9_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1012 (.I0(n26557), .I1(n20_adj_4560), .I2(n16_adj_4559), 
            .I3(\data_in_frame[9] [2]), .O(n43432));   // verilog/coms.v(73[16:42])
    defparam i10_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1013 (.I0(n41082), .I1(n43123), .I2(\data_in_frame[19] [0]), 
            .I3(n27189), .O(n12_adj_4561));
    defparam i5_4_lut_adj_1013.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_6 (.CI(n38238), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n38239));
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n38237), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1014 (.I0(n26744), .I1(n12_adj_4561), .I2(n43377), 
            .I3(n44609), .O(n40284));
    defparam i6_4_lut_adj_1014.LUT_INIT = 16'h9669;
    SB_CARRY add_3971_5 (.CI(n38237), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n38238));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n38236), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15085_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n28596));
    defparam i15085_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(n1510), .I1(n25928), .I2(GND_net), 
            .I3(GND_net), .O(n27288));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i15086_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n28597));
    defparam i15086_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(n40393), .I1(n27041), .I2(GND_net), 
            .I3(GND_net), .O(n41122));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1017 (.I0(n43241), .I1(n43386), .I2(n41122), 
            .I3(GND_net), .O(n43487));
    defparam i2_3_lut_adj_1017.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [7]), 
            .I2(n8_adj_4562), .I3(n27056), .O(n43045));   // verilog/coms.v(72[16:41])
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h9669;
    SB_LUT4 i15087_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n28598));
    defparam i15087_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1019 (.I0(n26557), .I1(n43340), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[16] [1]), .O(n12_adj_4563));   // verilog/coms.v(72[16:41])
    defparam i5_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1020 (.I0(\data_in_frame[13] [4]), .I1(n12_adj_4563), 
            .I2(\data_in_frame[18] [2]), .I3(n43045), .O(n43174));   // verilog/coms.v(72[16:41])
    defparam i6_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i20355_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), .I2(n63_adj_4469), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i20355_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i15088_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n28599));
    defparam i15088_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3971_4 (.CI(n38236), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n38237));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n38235), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43162));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 select_686_Select_2_i5_4_lut (.I0(n122), .I1(\FRAME_MATCHER.i_31__N_2624 ), 
            .I2(n3303), .I3(n63), .O(n5));
    defparam select_686_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_CARRY add_3971_3 (.CI(n38235), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n38236));
    SB_LUT4 i3_4_lut_adj_1022 (.I0(\data_in_frame[19] [7]), .I1(n40582), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[19] [1]), .O(n8_adj_4565));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3513), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1023 (.I0(\data_in_frame[19] [3]), .I1(n8_adj_4565), 
            .I2(n43162), .I3(\data_in_frame[19] [2]), .O(n43241));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1024 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n43305));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1024.LUT_INIT = 16'h9696;
    SB_LUT4 i20345_rep_265_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n49229));   // verilog/coms.v(142[4] 144[7])
    defparam i20345_rep_265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33674_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n34377), .I3(\FRAME_MATCHER.state [2]), .O(n44811));
    defparam i33674_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1025 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n130));
    defparam i1_2_lut_3_lut_adj_1025.LUT_INIT = 16'h1010;
    SB_LUT4 i20650_2_lut_3_lut (.I0(n63_adj_4469), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(139[4] 141[7])
    defparam i20650_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5_3_lut_adj_1026 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[10] [7]), 
            .I2(n43293), .I3(GND_net), .O(n14_adj_4566));
    defparam i5_3_lut_adj_1026.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1027 (.I0(n43468), .I1(\data_in_frame[17] [3]), 
            .I2(\data_in_frame[14] [7]), .I3(n43453), .O(n15_adj_4567));
    defparam i6_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1028 (.I0(n15_adj_4567), .I1(n42949), .I2(n14_adj_4566), 
            .I3(n27103), .O(n27174));
    defparam i8_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[17] [1]), .I1(n27174), 
            .I2(GND_net), .I3(GND_net), .O(n42878));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1030 (.I0(\data_in_frame[18] [3]), .I1(n43508), 
            .I2(n43039), .I3(\data_in_frame[16] [1]), .O(n10_adj_4568));
    defparam i4_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1031 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(n42984), .I3(n6_adj_4569), .O(n26832));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[16] [1]), .I1(n40326), .I2(n44005), 
            .I3(n26676), .O(n43417));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4570));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1033 (.I0(\data_in_frame[16] [4]), .I1(n4_adj_4570), 
            .I2(n41149), .I3(\data_in_frame[14] [2]), .O(n43377));
    defparam i2_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1034 (.I0(\data_out_frame[16] [1]), .I1(n40326), 
            .I2(n43484), .I3(n43398), .O(n41115));
    defparam i2_3_lut_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3513), 
            .CO(n38235));
    SB_LUT4 add_43_33_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n38234), .O(n2_adj_4526)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n38233), .O(n2_adj_4524)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1035 (.I0(n40244), .I1(\data_out_frame[10] [0]), 
            .I2(n26832), .I3(\data_out_frame[11] [0]), .O(n15_adj_4571));
    defparam i6_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_CARRY add_43_32 (.CI(n38233), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n38234));
    SB_LUT4 i8_4_lut_adj_1036 (.I0(n15_adj_4571), .I1(n27234), .I2(n14_adj_4572), 
            .I3(n1516), .O(n43257));
    defparam i8_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i31301_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46382));
    defparam i31301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1037 (.I0(n26860), .I1(n43257), .I2(n42864), 
            .I3(n26083), .O(n44677));
    defparam i3_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i31302_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46383));
    defparam i31302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31308_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46389));
    defparam i31308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_31_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n38232), .O(n2_adj_4522)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n38232), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n38233));
    SB_LUT4 i31307_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21][3] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46388));
    defparam i31307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1038 (.I0(\data_out_frame[11] [3]), .I1(n43183), 
            .I2(n43257), .I3(n6_adj_4573), .O(n41182));
    defparam i4_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1039 (.I0(n26840), .I1(\data_out_frame[18] [4]), 
            .I2(n41182), .I3(n44677), .O(n10_adj_4574));
    defparam i4_4_lut_adj_1039.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1040 (.I0(n27145), .I1(n26735), .I2(n43035), 
            .I3(n6_adj_4575), .O(n43474));
    defparam i4_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_out_frame[5] [0]), .I1(n1168), .I2(\data_out_frame[4] [5]), 
            .I3(\data_out_frame[6] [7]), .O(n43145));   // verilog/coms.v(85[17:70])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n48849), .I2(n47236), .I3(byte_transmit_counter[4]), .O(n48924));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48924_bdd_4_lut (.I0(n48924), .I1(n48807), .I2(n7_adj_4576), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n48924_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n46331), .I2(n46332), .I3(byte_transmit_counter[2]), .O(n48918));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48918_bdd_4_lut (.I0(n48918), .I1(n46392), .I2(n46391), .I3(byte_transmit_counter[2]), 
            .O(n47663));
    defparam n48918_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33816 (.I0(byte_transmit_counter[3]), 
            .I1(n47663), .I2(n47249), .I3(byte_transmit_counter[4]), .O(n48912));
    defparam byte_transmit_counter_3__bdd_4_lut_33816.LUT_INIT = 16'he4aa;
    SB_LUT4 n48912_bdd_4_lut (.I0(n48912), .I1(n48825), .I2(n7_adj_4577), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n48912_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1041 (.I0(\data_in_frame[13] [7]), .I1(n27053), 
            .I2(\data_in_frame[8] [2]), .I3(n41096), .O(n18_adj_4578));
    defparam i7_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1042 (.I0(n43334), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[9] [1]), .I3(n41094), .O(n19_adj_4579));
    defparam i8_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1043 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n43171));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1043.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1044 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n43281), .I3(GND_net), .O(n1168));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(n43353), .I1(n41115), .I2(\data_out_frame[18] [3]), 
            .I3(GND_net), .O(n42891));
    defparam i3_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(n26637), .I2(\data_in_frame[2] [6]), 
            .I3(n10_adj_4580), .O(n43120));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27122));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 i31246_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n46327));
    defparam i31246_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i31244_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46325));
    defparam i31244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut (.I0(n63_adj_4469), .I1(n63_c), .I2(n63), .I3(GND_net), 
            .O(n23534));   // verilog/coms.v(139[4] 141[7])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1046 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[3] [2]), .O(n43350));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1047 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n42907));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1048 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[4] [3]), .I3(GND_net), .O(n6_adj_4581));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1049 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n6_adj_4582));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1049.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n28177));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1050 (.I0(\data_in_frame[14] [1]), .I1(n19_adj_4579), 
            .I2(n17_adj_4583), .I3(n18_adj_4578), .O(n41169));
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_30_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n38231), .O(n2_adj_4519)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10_4_lut_adj_1051 (.I0(n43474), .I1(n42963), .I2(n43099), 
            .I3(n42915), .O(n24));
    defparam i10_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1052 (.I0(n43505), .I1(n43011), .I2(\data_in_frame[6] [5]), 
            .I3(n40197), .O(n22));
    defparam i8_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n43374), .I1(n24), .I2(n18_adj_4584), .I3(n42928), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1053 (.I0(\data_in_frame[3] [5]), .I1(n43177), 
            .I2(n43102), .I3(\data_in_frame[1] [6]), .O(Kp_23__N_936));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n38231), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n38232));
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[6] [0]), .I1(n26), .I2(n22), 
            .I3(n40225), .O(n41149));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32248_2_lut (.I0(n48939), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47248));
    defparam i32248_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n28176));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_out_frame[15] [4]), .I1(n43407), 
            .I2(GND_net), .I3(GND_net), .O(n43499));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1055 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_1096), 
            .I2(\data_in_frame[8] [5]), .I3(n27145), .O(n27377));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i31239_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46320));
    defparam i31239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1056 (.I0(\data_in_frame[6] [4]), .I1(Kp_23__N_1096), 
            .I2(\data_in_frame[6] [5]), .I3(Kp_23__N_1099), .O(Kp_23__N_1195));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1057 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [4]), .I3(GND_net), .O(n43523));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1057.LUT_INIT = 16'h9696;
    SB_LUT4 i31240_4_lut (.I0(n46320), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n46321));
    defparam i31240_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i4_4_lut_adj_1058 (.I0(n43496), .I1(n43395), .I2(n26676), 
            .I3(n43499), .O(n10_adj_4585));
    defparam i4_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33806 (.I0(byte_transmit_counter[3]), 
            .I1(n48873), .I2(n47240), .I3(byte_transmit_counter[4]), .O(n48906));
    defparam byte_transmit_counter_3__bdd_4_lut_33806.LUT_INIT = 16'he4aa;
    SB_LUT4 i31238_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46319));
    defparam i31238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1059 (.I0(\data_in_frame[5] [5]), .I1(n42957), 
            .I2(n42955), .I3(GND_net), .O(n40294));
    defparam i1_2_lut_3_lut_adj_1059.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1060 (.I0(n41149), .I1(n41169), .I2(\data_in_frame[14] [2]), 
            .I3(GND_net), .O(n44813));
    defparam i2_3_lut_adj_1060.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1061 (.I0(n26504), .I1(n44813), .I2(\data_in_frame[18] [4]), 
            .I3(\data_in_frame[11] [4]), .O(n43343));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(n44105), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43123));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n28175));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i32376_2_lut (.I0(n48945), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n47247));
    defparam i32376_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1063 (.I0(\data_in_frame[5] [5]), .I1(n42957), 
            .I2(\data_in_frame[10] [2]), .I3(GND_net), .O(n9_adj_4586));
    defparam i1_2_lut_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1064 (.I0(\data_in_frame[5] [5]), .I1(n42957), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n43035));
    defparam i1_2_lut_3_lut_adj_1064.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n28715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n28714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n28713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n28712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i218 (.Q(\data_out_frame[27][1] ), .C(CLK_c), 
           .D(n28711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n28710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n28709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n28708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n28707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n28706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n28705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n28704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n28703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n28702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n28701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n28700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n28699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n28698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n28697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n28696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n28695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n28694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n28693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n28692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n28691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n28690));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1065 (.I0(\data_out_frame[10] [5]), .I1(n42925), 
            .I2(\data_out_frame[13] [1]), .I3(\data_out_frame[12] [7]), 
            .O(n10_adj_4587));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1065.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n28689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n28688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n28687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n28686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n28685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n28684));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1066 (.I0(n9_adj_4588), .I1(n43123), .I2(n8_adj_4589), 
            .I3(\data_in_frame[16] [5]), .O(n44609));
    defparam i5_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i15072_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n28583));
    defparam i15072_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31280_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46361));
    defparam i31280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31281_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46362));
    defparam i31281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15073_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n28584));
    defparam i15073_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n28683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n28174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n28173));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15074_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n28585));
    defparam i15074_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n28172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n28171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21][0] ), .C(CLK_c), 
           .D(n28170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21][1] ), .C(CLK_c), 
           .D(n28169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21][2] ), .C(CLK_c), 
           .D(n28168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21][3] ), .C(CLK_c), 
           .D(n28167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21][4] ), .C(CLK_c), 
           .D(n28166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(CLK_c), 
           .D(n28165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(CLK_c), 
           .D(n28164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(CLK_c), 
           .D(n28163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(CLK_c), 
           .D(n28162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(CLK_c), 
           .D(n28161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(CLK_c), 
           .D(n28160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(CLK_c), 
           .D(n28156));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[18] [7]), .I1(n44609), 
            .I2(GND_net), .I3(GND_net), .O(n43202));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(CLK_c), 
           .D(n28152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n28151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
           .D(n42180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27522));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n28148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n28147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n28146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n28145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n28144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n28143));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31287_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46368));
    defparam i31287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31286_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21][2] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46367));
    defparam i31286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n23534), .I1(n42849), .I2(n3813), .I3(\FRAME_MATCHER.state_c [13]), 
            .O(n42222));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hec00;
    SB_LUT4 i15075_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n28586));
    defparam i15075_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1069 (.I0(n23534), .I1(n42849), .I2(n3813), 
            .I3(\FRAME_MATCHER.state_c [14]), .O(n42220));
    defparam i1_2_lut_4_lut_adj_1069.LUT_INIT = 16'hec00;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n44811), .D(n141), 
            .R(n34718));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15076_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n28587));
    defparam i15076_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_29_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n38230), .O(n2_adj_4517)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15078_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n28589));
    defparam i15078_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n44876), .D(n75), .R(n45195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n28682));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15079_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n28590));
    defparam i15079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15080_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n28591));
    defparam i15080_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1070 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4591));   // verilog/coms.v(85[17:63])
    defparam i2_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1071 (.I0(n23534), .I1(n42849), .I2(n3813), 
            .I3(\FRAME_MATCHER.state_c [15]), .O(n42218));
    defparam i1_2_lut_4_lut_adj_1071.LUT_INIT = 16'hec00;
    SB_LUT4 n48906_bdd_4_lut (.I0(n48906), .I1(n48819), .I2(n7_adj_4592), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n48906_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15024_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n28535));
    defparam i15024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15032_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n28543));
    defparam i15032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_29 (.CI(n38230), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n38231));
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n28681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n28680));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n28679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n28678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n28677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n28676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n28675));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1072 (.I0(n43302), .I1(n42975), .I2(n7_adj_4591), 
            .I3(n8_adj_4594), .O(n42925));   // verilog/coms.v(85[17:63])
    defparam i2_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n28674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n28673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n28672));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n28671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n28670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n28669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n28668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n28667));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n28666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n28665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n28664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n28663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n28662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n28661));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n28660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n28659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n28658));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n28657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n28656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n28655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n28654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n28653));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_28_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n38229), .O(n2_adj_4513)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1073 (.I0(\data_out_frame[14] [1]), .I1(n43077), 
            .I2(n26656), .I3(n43459), .O(n16_adj_4595));
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n28652));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1074 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n43293));
    defparam i2_3_lut_adj_1074.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1075 (.I0(n42925), .I1(n43299), .I2(n27425), 
            .I3(n43049), .O(n17_adj_4596));
    defparam i7_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33811 (.I0(byte_transmit_counter[1]), 
            .I1(n46349), .I2(n46350), .I3(byte_transmit_counter[2]), .O(n48900));
    defparam byte_transmit_counter_1__bdd_4_lut_33811.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43526));
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1077 (.I0(n23534), .I1(n42849), .I2(n3813), 
            .I3(\FRAME_MATCHER.state_c [16]), .O(n42216));
    defparam i1_2_lut_4_lut_adj_1077.LUT_INIT = 16'hec00;
    SB_LUT4 i9_4_lut_adj_1078 (.I0(n17_adj_4596), .I1(n41242), .I2(n16_adj_4595), 
            .I3(n26843), .O(n43429));
    defparam i9_4_lut_adj_1078.LUT_INIT = 16'h9669;
    SB_LUT4 i15035_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n28546));
    defparam i15035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43299));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i15067_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n28578));
    defparam i15067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n48900_bdd_4_lut (.I0(n48900), .I1(n46347), .I2(n46346), .I3(byte_transmit_counter[2]), 
            .O(n47638));
    defparam n48900_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42975));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'h6666;
    SB_LUT4 i15068_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n28579));
    defparam i15068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_in_frame[12] [6]), .I1(n27377), 
            .I2(GND_net), .I3(GND_net), .O(n43453));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n28651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n28650));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1082 (.I0(n43471), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[8] [6]), .I3(n43328), .O(n15_adj_4597));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i15069_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n28580));
    defparam i15069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n28649));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1083 (.I0(n40225), .I1(n43222), .I2(GND_net), 
            .I3(GND_net), .O(n41094));
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(\data_in_frame[11] [6]), .I1(n41094), 
            .I2(n40336), .I3(n41098), .O(n43505));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1085 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(n27050), .I3(GND_net), .O(n43340));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27053));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1087 (.I0(n23534), .I1(n1), .I2(n9), .I3(\FRAME_MATCHER.state_c [13]), 
            .O(n42292));
    defparam i1_2_lut_4_lut_adj_1087.LUT_INIT = 16'hec00;
    SB_LUT4 i8_4_lut_adj_1088 (.I0(n15_adj_4597), .I1(n42975), .I2(n14_adj_4598), 
            .I3(n27262), .O(n27031));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i15070_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n28581));
    defparam i15070_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15071_3_lut_4_lut (.I0(n10_adj_4593), .I1(n42810), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n28582));
    defparam i15071_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1089 (.I0(n42928), .I1(n43284), .I2(\data_in_frame[4] [5]), 
            .I3(\data_in_frame[6] [6]), .O(n12_adj_4599));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_out_frame[13] [7]), .I1(n43429), 
            .I2(GND_net), .I3(GND_net), .O(n42864));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33796 (.I0(byte_transmit_counter[1]), 
            .I1(n46367), .I2(n46368), .I3(byte_transmit_counter[2]), .O(n48894));
    defparam byte_transmit_counter_1__bdd_4_lut_33796.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n28648));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1091 (.I0(\data_in_frame[7] [0]), .I1(n12_adj_4599), 
            .I2(n43447), .I3(\data_in_frame[7] [1]), .O(Kp_23__N_1330));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 n48894_bdd_4_lut (.I0(n48894), .I1(n46362), .I2(n46361), .I3(byte_transmit_counter[2]), 
            .O(n47640));
    defparam n48894_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n28647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n28646));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33801 (.I0(byte_transmit_counter[3]), 
            .I1(n47640), .I2(n47247), .I3(byte_transmit_counter[4]), .O(n48888));
    defparam byte_transmit_counter_3__bdd_4_lut_33801.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n28645));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48888_bdd_4_lut (.I0(n48888), .I1(n48813), .I2(n7_adj_4600), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n48888_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n28644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n28643));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1092 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n41230), .I3(GND_net), .O(n43065));
    defparam i2_3_lut_adj_1092.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33786 (.I0(byte_transmit_counter[3]), 
            .I1(n47638), .I2(n47248), .I3(byte_transmit_counter[4]), .O(n48882));
    defparam byte_transmit_counter_3__bdd_4_lut_33786.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n28642));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48882_bdd_4_lut (.I0(n48882), .I1(n48855), .I2(n7_adj_4601), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n48882_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n28641));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n28640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n28639));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n28638));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n28637));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33791 (.I0(byte_transmit_counter[1]), 
            .I1(n46388), .I2(n46389), .I3(byte_transmit_counter[2]), .O(n48870));
    defparam byte_transmit_counter_1__bdd_4_lut_33791.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n28636));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48870_bdd_4_lut (.I0(n48870), .I1(n46383), .I2(n46382), .I3(byte_transmit_counter[2]), 
            .O(n48873));
    defparam n48870_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n28635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n28634));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1093 (.I0(n43108), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[13] [3]), .I3(n43145), .O(n10_adj_4602));
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33826 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48864));
    defparam byte_transmit_counter_0__bdd_4_lut_33826.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n28633));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48864_bdd_4_lut (.I0(n48864), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48867));
    defparam n48864_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n28632));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n49000));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33768 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48858));
    defparam byte_transmit_counter_0__bdd_4_lut_33768.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n28630));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48858_bdd_4_lut (.I0(n48858), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48861));
    defparam n48858_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n28629));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n28628));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33773 (.I0(byte_transmit_counter[1]), 
            .I1(n46442), .I2(n46443), .I3(byte_transmit_counter[2]), .O(n48852));
    defparam byte_transmit_counter_1__bdd_4_lut_33773.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n28627));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48852_bdd_4_lut (.I0(n48852), .I1(n46449), .I2(n46448), .I3(byte_transmit_counter[2]), 
            .O(n48855));
    defparam n48852_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n28626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n28625));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1094 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[13] [3]), 
            .I2(Kp_23__N_1306), .I3(n10_adj_4603), .O(n16_adj_4604));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33758 (.I0(byte_transmit_counter[1]), 
            .I1(n46430), .I2(n46431), .I3(byte_transmit_counter[2]), .O(n48846));
    defparam byte_transmit_counter_1__bdd_4_lut_33758.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n28624));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1095 (.I0(\data_in_frame[9] [3]), .I1(n40205), 
            .I2(n43083), .I3(\data_in_frame[10] [7]), .O(n11_adj_4605));   // verilog/coms.v(74[16:43])
    defparam i2_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 n48846_bdd_4_lut (.I0(n48846), .I1(n46356), .I2(n46355), .I3(byte_transmit_counter[2]), 
            .O(n48849));
    defparam n48846_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33753 (.I0(byte_transmit_counter[1]), 
            .I1(n46271), .I2(n46272), .I3(byte_transmit_counter[2]), .O(n48834));
    defparam byte_transmit_counter_1__bdd_4_lut_33753.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1096 (.I0(n26717), .I1(n42995), .I2(\data_in_frame[8] [6]), 
            .I3(\data_in_frame[8] [7]), .O(n43520));
    defparam i2_3_lut_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43049));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1098 (.I0(n26083), .I1(n24464), .I2(n43429), 
            .I3(GND_net), .O(n6_adj_4573));
    defparam i1_2_lut_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1099 (.I0(\data_out_frame[7] [5]), .I1(n43049), 
            .I2(n27306), .I3(\data_out_frame[8] [0]), .O(n12_adj_4606));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1100 (.I0(\data_out_frame[9] [6]), .I1(n12_adj_4606), 
            .I2(n43142), .I3(\data_out_frame[5] [6]), .O(n1510));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1101 (.I0(\data_out_frame[14] [4]), .I1(n1510), 
            .I2(\data_out_frame[12] [2]), .I3(GND_net), .O(n42938));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1101.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n28611));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_1102 (.I0(n11_adj_4605), .I1(n16_adj_4604), .I2(n25962), 
            .I3(n43105), .O(n43003));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1103 (.I0(n26557), .I1(n43065), .I2(Kp_23__N_1330), 
            .I3(GND_net), .O(n43052));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n28610));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n28609));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1104 (.I0(n23534), .I1(n1), .I2(n9), .I3(\FRAME_MATCHER.state_c [15]), 
            .O(n42298));
    defparam i1_2_lut_4_lut_adj_1104.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_3_lut_adj_1105 (.I0(n26702), .I1(n8_adj_4607), .I2(\data_in_frame[9] [1]), 
            .I3(GND_net), .O(n26557));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[15] [5]), .I1(n43003), 
            .I2(GND_net), .I3(GND_net), .O(n43004));
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43105));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1108 (.I0(\data_in_frame[17] [7]), .I1(n43004), 
            .I2(n43052), .I3(n6_adj_4608), .O(n40675));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1108.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(n41193), .I1(n26656), .I2(GND_net), 
            .I3(GND_net), .O(n41242));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1110 (.I0(n27149), .I1(n4_adj_4609), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n27047));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1111 (.I0(n27149), .I1(n4_adj_4609), .I2(\data_in_frame[16] [2]), 
            .I3(GND_net), .O(n43480));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1112 (.I0(n27149), .I1(n4_adj_4609), 
            .I2(n26755), .I3(n40699), .O(n43083));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1113 (.I0(n23534), .I1(n1), .I2(n9), .I3(\FRAME_MATCHER.state_c [16]), 
            .O(n42302));
    defparam i1_2_lut_4_lut_adj_1113.LUT_INIT = 16'hec00;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43328));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1115 (.I0(n43340), .I1(\data_in_frame[11] [5]), 
            .I2(n43065), .I3(n40393), .O(n14_adj_4610));
    defparam i6_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1116 (.I0(\data_in_frame[18] [0]), .I1(n14_adj_4610), 
            .I2(n10_adj_4611), .I3(\data_in_frame[11] [4]), .O(n40582));
    defparam i7_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(n40582), .I1(n40675), .I2(GND_net), 
            .I3(GND_net), .O(n43093));
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n28608));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1118 (.I0(\data_in_frame[11] [2]), .I1(n43251), 
            .I2(n43505), .I3(\data_in_frame[10] [1]), .O(n32));
    defparam i12_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 equal_286_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4590));   // verilog/coms.v(154[7:23])
    defparam equal_286_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i3_3_lut_4_lut (.I0(n40699), .I1(n26755), .I2(\data_in_frame[13] [6]), 
            .I3(\data_in_frame[11] [6]), .O(n8_adj_4562));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n28607));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n28606));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31265_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46346));
    defparam i31265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31266_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46347));
    defparam i31266_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_28 (.CI(n38229), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n38230));
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[12] [5]), 
            .I2(n43453), .I3(n43132), .O(n31_adj_4612));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31269_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46350));
    defparam i31269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_4_lut_adj_1119 (.I0(\data_in_frame[10] [2]), .I1(n40699), 
            .I2(\data_in_frame[11] [0]), .I3(n41230), .O(n35));
    defparam i15_4_lut_adj_1119.LUT_INIT = 16'h9669;
    SB_LUT4 i31268_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21][1] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n46349));
    defparam i31268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43015));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1121 (.I0(n42987), .I1(n10_adj_4613), .I2(n27103), 
            .I3(\data_in_frame[15] [4]), .O(n42867));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1122 (.I0(n43311), .I1(n27047), .I2(n43151), 
            .I3(\data_in_frame[10] [3]), .O(n34));
    defparam i14_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43471));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n28109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n28106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n28105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n28104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n28103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n28102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n28101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n28100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n28099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n28098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n28097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n28095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n28094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n28093));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1124 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n43459));
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1125 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[10] [1]), .I3(n6_adj_4614), .O(n43021));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1126 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n10_adj_4615));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_adj_1126.LUT_INIT = 16'hfbfb;
    SB_LUT4 i13_2_lut_4_lut (.I0(n42987), .I1(n10_adj_4613), .I2(n27103), 
            .I3(\data_in_frame[18] [2]), .O(n39_adj_4616));   // verilog/coms.v(75[16:43])
    defparam i13_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n27605), .D(n7025));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i18_4_lut_adj_1127 (.I0(\data_out_frame[8] [3]), .I1(n43318), 
            .I2(n43471), .I3(n43171), .O(n44_adj_4617));
    defparam i18_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n27605), .D(n7024));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n27605), .D(n7023));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n27605), .D(n7022));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n27605), .D(n7021));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n27605), .D(n7020));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n27605), .D(n7019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n27605), .D(n7018));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n27605), .D(n7017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n27605), .D(n7016));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n27605), .D(n7015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n27605), .D(n7014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n27605), .D(n7013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n27605), .D(n7012));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n27605), .D(n7011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n27605), .D(n7010));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n27605), .D(n7009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n27605), .D(n7008));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n27605), .D(n7007));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n27605), .D(n7006));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n27605), .D(n7005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n27605), .D(n7004));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n27605), .D(n7003));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i18_3_lut (.I0(n35), .I1(n31_adj_4612), .I2(n32), .I3(GND_net), 
            .O(n38));
    defparam i18_3_lut.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(CLK_c), 
            .D(n42268), .S(n42168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n28092));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13_4_lut_adj_1128 (.I0(\data_in_frame[11] [3]), .I1(n43526), 
            .I2(\data_in_frame[11] [4]), .I3(n43502), .O(n33));
    defparam i13_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1129 (.I0(\data_in_frame[15] [3]), .I1(n33), .I2(n38), 
            .I3(n34), .O(n32_adj_4618));
    defparam i6_4_lut_adj_1129.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1130 (.I0(n43293), .I1(n43039), .I2(n43202), 
            .I3(n43008), .O(n44_adj_4619));
    defparam i18_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1131 (.I0(\data_out_frame[9] [7]), .I1(n43462), 
            .I2(n42969), .I3(n1191), .O(n42_adj_4620));
    defparam i16_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1132 (.I0(n27296), .I1(\data_out_frame[8] [0]), 
            .I2(n43314), .I3(\data_out_frame[7] [6]), .O(n43_adj_4621));
    defparam i17_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1133 (.I0(\data_in_frame[18] [1]), .I1(n32_adj_4618), 
            .I2(n43031), .I3(n43371), .O(n42_adj_4622));
    defparam i16_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 n48834_bdd_4_lut (.I0(n48834), .I1(n46398), .I2(n46397), .I3(byte_transmit_counter[2]), 
            .O(n48837));
    defparam n48834_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i17_4_lut_adj_1134 (.I0(n43004), .I1(n43456), .I2(n43517), 
            .I3(n43343), .O(n43_adj_4623));
    defparam i17_4_lut_adj_1134.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n28604));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1135 (.I0(n43165), .I1(n27041), .I2(\data_in_frame[14] [0]), 
            .I3(n43377), .O(n41_adj_4624));
    defparam i15_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1136 (.I0(n43308), .I1(n43003), .I2(\data_in_frame[13] [7]), 
            .I3(n43490), .O(n40_adj_4625));
    defparam i14_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1137 (.I0(n41_adj_4624), .I1(n43_adj_4623), .I2(n42_adj_4622), 
            .I3(n44_adj_4619), .O(n50_adj_4626));
    defparam i24_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1138 (.I0(n42878), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[14] [1]), .I3(\data_in_frame[14] [2]), .O(n45_adj_4627));
    defparam i19_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 equal_287_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4471));   // verilog/coms.v(154[7:23])
    defparam equal_287_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1139 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [1]), 
            .I2(n43356), .I3(\data_out_frame[9] [0]), .O(n41_adj_4628));
    defparam i15_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_27_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n38228), .O(n2_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i25_4_lut_adj_1140 (.I0(n45_adj_4627), .I1(n50_adj_4626), .I2(n39_adj_4616), 
            .I3(n40_adj_4625), .O(n41117));
    defparam i25_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n40922), .I1(\data_in_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43456));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1378_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n44527), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n34624), .O(n4888[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_1378_i1_3_lut_4_lut.LUT_INIT = 16'h333a;
    SB_LUT4 i14_4_lut_adj_1142 (.I0(\data_out_frame[9] [5]), .I1(n43444), 
            .I2(n43158), .I3(\data_out_frame[8] [2]), .O(n40_adj_4629));
    defparam i14_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i13_2_lut_adj_1143 (.I0(n26915), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4630));
    defparam i13_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1144 (.I0(\data_out_frame[22] [6]), .I1(n10_adj_4631), 
            .I2(n41204), .I3(n40347), .O(n41208));
    defparam i5_3_lut_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1145 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[12] [2]), .I3(GND_net), .O(n43151));
    defparam i2_3_lut_adj_1145.LUT_INIT = 16'h9696;
    SB_LUT4 i24_4_lut_adj_1146 (.I0(n41_adj_4628), .I1(n43_adj_4621), .I2(n42_adj_4620), 
            .I3(n44_adj_4617), .O(n50_adj_4632));
    defparam i24_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_CARRY add_43_27 (.CI(n38228), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n38229));
    SB_LUT4 i1_2_lut_adj_1147 (.I0(n40699), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41098));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1148 (.I0(n41098), .I1(n40225), .I2(n43296), 
            .I3(n6_adj_4633), .O(n44105));
    defparam i4_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_26_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n38227), .O(n2_adj_4509)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut_4_lut (.I0(n63), .I1(n771), .I2(\FRAME_MATCHER.i_31__N_2620 ), 
            .I3(n4), .O(n7));   // verilog/coms.v(157[6] 159[9])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'haa20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1149 (.I0(\data_out_frame[23] [1]), .I1(n41137), 
            .I2(\data_out_frame[22] [6]), .I3(\data_out_frame[23] [0]), 
            .O(n6_adj_4540));
    defparam i1_2_lut_3_lut_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 select_686_Select_1_i1_3_lut_4_lut (.I0(n63), .I1(n771), .I2(\FRAME_MATCHER.i_31__N_2620 ), 
            .I3(n92[1]), .O(n1_adj_4476));   // verilog/coms.v(157[6] 159[9])
    defparam select_686_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'hf0d0;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43371));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1151 (.I0(n42854), .I1(n4_adj_4535), 
            .I2(\FRAME_MATCHER.state_c [4]), .I3(n4_adj_4544), .O(n36539));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1151.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_26 (.CI(n38227), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n38228));
    SB_LUT4 add_43_25_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n38226), .O(n2_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1152 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n43359));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i20938_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n34442));
    defparam i20938_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i19_4_lut_adj_1153 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[7] [1]), .I3(n26456), .O(n45_adj_4636));
    defparam i19_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n28603));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1154 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(\data_out_frame[7] [0]), .O(n27421));
    defparam i1_2_lut_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n28602));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_25 (.CI(n38226), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n38227));
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n43287), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[15] [3]), .I3(\data_in_frame[15] [2]), .O(n14_adj_4637));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1156 (.I0(n9_adj_4638), .I1(n14_adj_4637), .I2(n42932), 
            .I3(n41143), .O(n27041));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(n27041), .I1(n41113), .I2(GND_net), 
            .I3(GND_net), .O(n41184));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i25_4_lut_adj_1158 (.I0(n45_adj_4636), .I1(n50_adj_4632), .I2(n39_adj_4630), 
            .I3(n40_adj_4629), .O(n41193));
    defparam i25_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(n26747), .I1(n26755), .I2(GND_net), 
            .I3(GND_net), .O(n43132));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1160 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[18] [7]), 
            .I2(n44609), .I3(GND_net), .O(n6_adj_4639));
    defparam i1_2_lut_3_lut_adj_1160.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[17] [1]), 
            .I2(n27174), .I3(GND_net), .O(n6_adj_4640));
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1162 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[17] [7]), .I3(\data_in_frame[17] [6]), .O(n5_adj_4641));
    defparam i1_3_lut_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1163 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n42921));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1164 (.I0(n41193), .I1(n43021), .I2(GND_net), 
            .I3(GND_net), .O(n40244));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1164.LUT_INIT = 16'h9999;
    SB_LUT4 add_43_24_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n38225), .O(n2_adj_4505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut_4_lut_adj_1165 (.I0(Kp_23__N_1189), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_1195), .I3(\data_in_frame[8] [6]), .O(n13));
    defparam i3_3_lut_4_lut_adj_1165.LUT_INIT = 16'h6ff6;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(\data_in_frame[4] [3]), .I3(GND_net), .O(n18_adj_4642));   // verilog/coms.v(74[16:43])
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_out_frame[8] [5]), .I1(n1247), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n43356));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1167 (.I0(n43356), .I1(n27360), .I2(\data_out_frame[11] [7]), 
            .I3(n40244), .O(n16_adj_4643));
    defparam i6_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_CARRY add_43_24 (.CI(n38225), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n38226));
    SB_LUT4 i2_3_lut_4_lut_adj_1168 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[1] [4]), .O(n27403));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_23_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n38224), .O(n2_adj_4499)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1169 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [1]), .O(n27078));
    defparam i1_2_lut_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1170 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n42966));
    defparam i1_2_lut_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_CARRY add_43_23 (.CI(n38224), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n38225));
    SB_LUT4 i7_4_lut_adj_1171 (.I0(\data_out_frame[5] [5]), .I1(n43071), 
            .I2(\data_out_frame[7] [6]), .I3(n41242), .O(n17_adj_4644));
    defparam i7_4_lut_adj_1171.LUT_INIT = 16'h9669;
    SB_LUT4 equal_285_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4645));   // verilog/coms.v(154[7:23])
    defparam equal_285_i7_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_adj_1172 (.I0(n26593), .I1(\data_in_frame[4] [4]), 
            .I2(n26599), .I3(GND_net), .O(n27072));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1172.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_22_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n38223), .O(n2_adj_4497)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1173 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [7]), .I3(GND_net), .O(n26604));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1173.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1174 (.I0(n17_adj_4644), .I1(n43021), .I2(n16_adj_4643), 
            .I3(\data_out_frame[10] [0]), .O(n25928));
    defparam i9_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1175 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(n42960), .I3(\data_in_frame[3] [0]), .O(n27253));
    defparam i2_3_lut_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_CARRY add_43_22 (.CI(n38223), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n38224));
    SB_LUT4 i1_2_lut_3_lut_adj_1176 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[5] [5]), 
            .I2(n43350), .I3(GND_net), .O(n26545));
    defparam i1_2_lut_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1177 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[12] [3]), 
            .I2(n1513), .I3(n42938), .O(n42881));
    defparam i1_2_lut_3_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1178 (.I0(n26580), .I1(\data_in_frame[4] [7]), 
            .I2(n27500), .I3(GND_net), .O(n27059));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1178.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1179 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5] [3]), 
            .I2(n26905), .I3(GND_net), .O(n43426));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1179.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1180 (.I0(n26580), .I1(n42928), .I2(n43011), 
            .I3(n27258), .O(n4_adj_4609));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[11] [6]), .I3(\data_out_frame[12] [1]), 
            .O(n10_adj_4646));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4647));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1182 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n27062));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43077));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1184 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n26593));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1185 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26580));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1185.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1186 (.I0(\data_in_frame[10] [3]), .I1(\data_in_frame[8] [1]), 
            .I2(n26730), .I3(n24669), .O(n27189));
    defparam i1_2_lut_3_lut_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1187 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n6_adj_4648));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43142));
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1189 (.I0(\data_out_frame[4] [3]), .I1(n42969), 
            .I2(n10_adj_4587), .I3(n26915), .O(n27326));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1190 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[16] [7]), 
            .I2(n8_adj_4649), .I3(\data_in_frame[10] [4]), .O(n9_adj_4588));
    defparam i3_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1191 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(n26702), .I3(n26747), .O(n10_adj_4650));
    defparam i2_2_lut_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1192 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_1186), 
            .I2(n27377), .I3(GND_net), .O(n26624));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1192.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1193 (.I0(\data_out_frame[4] [3]), .I1(n42969), 
            .I2(\data_out_frame[8] [7]), .I3(n27421), .O(n43108));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_21_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n38222), .O(n2_adj_4495)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1194 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(n26702), .I3(GND_net), .O(n43334));
    defparam i1_2_lut_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1195 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n42963));
    defparam i1_2_lut_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1196 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[9] [5]), .I3(GND_net), .O(n43296));
    defparam i1_2_lut_3_lut_adj_1196.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1197 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(n26747), .I3(GND_net), .O(n43374));
    defparam i1_2_lut_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1198 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[10] [6]), .I3(GND_net), .O(n43311));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 equal_289_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4651));
    defparam equal_289_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i15014_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n28525));
    defparam i15014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1199 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [4]), 
            .I2(n40699), .I3(n27149), .O(n27056));
    defparam i1_2_lut_3_lut_4_lut_adj_1199.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1200 (.I0(n27152), .I1(n27377), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[10] [6]), .O(n43490));
    defparam i2_3_lut_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i15015_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n28526));
    defparam i15015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15016_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n28527));
    defparam i15016_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(n40922), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n41082));
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i15017_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n28528));
    defparam i15017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_21 (.CI(n38222), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n38223));
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n27425));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1203 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n27262));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1203.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_20_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n38221), .O(n2_adj_4493)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_1186), 
            .I2(n42949), .I3(\data_in_frame[17] [0]), .O(n8_adj_4649));
    defparam i3_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1205 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n27234));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1206 (.I0(\data_in_frame[12] [2]), .I1(Kp_23__N_1306), 
            .I2(n43132), .I3(\data_in_frame[10] [0]), .O(n43517));
    defparam i1_2_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43251));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1208 (.I0(n26604), .I1(\data_in_frame[10] [1]), 
            .I2(n43245), .I3(n42966), .O(n16_adj_4653));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1209 (.I0(\data_in_frame[8] [0]), .I1(n43238), 
            .I2(n43426), .I3(\data_in_frame[3] [1]), .O(n17_adj_4654));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1210 (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n9_adj_4638));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1210.LUT_INIT = 16'h9696;
    SB_LUT4 equal_292_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_4652));   // verilog/coms.v(154[7:23])
    defparam equal_292_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i9_4_lut_adj_1211 (.I0(n17_adj_4654), .I1(\data_in_frame[7] [7]), 
            .I2(n16_adj_4653), .I3(\data_in_frame[9] [7]), .O(n40922));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1212 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[12] [2]), .I3(n43456), .O(n6_adj_4633));
    defparam i1_2_lut_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i15019_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n28530));
    defparam i15019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15020_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n28531));
    defparam i15020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1213 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_1195), 
            .I2(n43520), .I3(n43526), .O(n6_adj_4575));
    defparam i1_2_lut_3_lut_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1214 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_1195), 
            .I2(n43520), .I3(\data_in_frame[11] [2]), .O(n27050));
    defparam i1_2_lut_3_lut_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1215 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n43158));   // verilog/coms.v(75[16:27])
    defparam i2_2_lut_3_lut_adj_1215.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1216 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[10] [3]), 
            .O(n6_adj_4614));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43165));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43287));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1219 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[4] [0]), .O(n26456));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1220 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[11] [3]), 
            .I2(n41117), .I3(GND_net), .O(n10_adj_4611));
    defparam i2_2_lut_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1221 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(n43225), .I3(GND_net), .O(n6_adj_4608));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_CARRY add_43_20 (.CI(n38221), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n38222));
    SB_LUT4 add_43_19_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n38220), .O(n2_adj_4491)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1222 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n42969));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1223 (.I0(n26702), .I1(n8_adj_4607), 
            .I2(Kp_23__N_1189), .I3(\data_in_frame[8] [4]), .O(n43465));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26735));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1225 (.I0(Kp_23__N_1189), .I1(Kp_23__N_1186), .I2(n26735), 
            .I3(\data_in_frame[12] [5]), .O(n43392));
    defparam i3_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1226 (.I0(n43331), .I1(n26662), .I2(n43028), 
            .I3(n40294), .O(n14_adj_4655));
    defparam i6_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1227 (.I0(n26083), .I1(n24464), .I2(\data_out_frame[11] [5]), 
            .I3(\data_out_frame[11] [4]), .O(n4_adj_4656));
    defparam i1_2_lut_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_CARRY add_43_19 (.CI(n38220), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n38221));
    SB_LUT4 i7_4_lut_adj_1228 (.I0(n9_adj_4586), .I1(n14_adj_4655), .I2(n43117), 
            .I3(n41086), .O(n44882));
    defparam i7_4_lut_adj_1228.LUT_INIT = 16'h9669;
    SB_LUT4 i15021_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n28532));
    defparam i15021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15022_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n28533));
    defparam i15022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1229 (.I0(\data_in_frame[12] [4]), .I1(n44882), 
            .I2(GND_net), .I3(GND_net), .O(n43193));
    defparam i1_2_lut_adj_1229.LUT_INIT = 16'h9999;
    SB_LUT4 add_43_18_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n38219), .O(n2_adj_4489)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2898_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4458));
    defparam i2898_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i15154_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n28665));
    defparam i15154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15155_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n28666));
    defparam i15155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1230 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[9] [4]), .I3(n41096), .O(n10_adj_4603));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1230.LUT_INIT = 16'h9669;
    SB_CARRY add_43_18 (.CI(n38219), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n38220));
    SB_LUT4 equal_2186_i8_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n42995), .I3(\data_in_frame[8] [7]), .O(n8_adj_4607));
    defparam equal_2186_i8_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_17_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n38218), .O(n2_adj_4485)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1231 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[8] [5]), .I3(n1247), .O(n27139));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(\data_in_frame[9] [4]), .I1(n40699), 
            .I2(n27149), .I3(GND_net), .O(n41230));
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1233 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[11] [1]), 
            .O(n14_adj_4598));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i15156_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n28667));
    defparam i15156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1234 (.I0(\data_in_frame[11] [5]), .I1(n26557), 
            .I2(n43065), .I3(Kp_23__N_1330), .O(n43039));
    defparam i1_2_lut_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(\data_out_frame[8] [5]), .I1(n1247), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n43302));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_CARRY add_43_17 (.CI(n38218), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n38219));
    SB_LUT4 i2_2_lut_adj_1236 (.I0(n43392), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4657));
    defparam i2_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33743 (.I0(byte_transmit_counter[1]), 
            .I1(n46295), .I2(n46296), .I3(byte_transmit_counter[2]), .O(n48828));
    defparam byte_transmit_counter_1__bdd_4_lut_33743.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1237 (.I0(n44237), .I1(\data_out_frame[15] [7]), 
            .I2(n10_adj_4585), .I3(n43323), .O(n44262));
    defparam i5_3_lut_4_lut_adj_1237.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1238 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(Kp_23__N_1093), .I3(Kp_23__N_1090), .O(Kp_23__N_1189));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 n48828_bdd_4_lut (.I0(n48828), .I1(n46395), .I2(n46394), .I3(byte_transmit_counter[2]), 
            .O(n48831));
    defparam n48828_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1239 (.I0(n43490), .I1(\data_in_frame[12] [7]), 
            .I2(n43287), .I3(\data_in_frame[15] [0]), .O(n14_adj_4658));
    defparam i6_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33738 (.I0(byte_transmit_counter[1]), 
            .I1(n46373), .I2(n46374), .I3(byte_transmit_counter[2]), .O(n48822));
    defparam byte_transmit_counter_1__bdd_4_lut_33738.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1240 (.I0(\data_in_frame[15] [1]), .I1(n14_adj_4658), 
            .I2(n10_adj_4657), .I3(n43193), .O(n41113));
    defparam i7_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1241 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[16] [6]), .I3(\data_out_frame[16] [4]), 
            .O(n43496));
    defparam i2_3_lut_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 n48822_bdd_4_lut (.I0(n48822), .I1(n46386), .I2(n46385), .I3(byte_transmit_counter[2]), 
            .O(n48825));
    defparam n48822_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1242 (.I0(\data_in_frame[14] [7]), .I1(n43165), 
            .I2(n41082), .I3(\data_in_frame[12] [6]), .O(n12_adj_4659));
    defparam i5_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1243 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(n27186), .O(n43331));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1244 (.I0(\data_in_frame[16] [7]), .I1(n12_adj_4659), 
            .I2(n43392), .I3(\data_in_frame[14] [5]), .O(n41188));
    defparam i6_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_16_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n38217), .O(n2_adj_4483)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[6] [3]), 
            .I2(\data_in_frame[6] [2]), .I3(\data_in_frame[6] [4]), .O(n18_adj_4584));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_out_frame[6] [6]), .I1(n43145), 
            .I2(GND_net), .I3(GND_net), .O(n27296));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(n26083), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[15] [7]), .I3(GND_net), .O(n43398));
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1247 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[1] [0]), 
            .I2(n42960), .I3(\data_in_frame[0] [5]), .O(n26905));
    defparam i1_2_lut_3_lut_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1248 (.I0(\data_in_frame[16] [6]), .I1(n27189), 
            .I2(\data_in_frame[17] [1]), .I3(n43193), .O(n11_adj_4660));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1248.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1249 (.I0(n11_adj_4660), .I1(n9_adj_4588), .I2(n41188), 
            .I3(n26744), .O(n26050));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1249.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1250 (.I0(n26050), .I1(n41188), .I2(n41113), 
            .I3(\data_in_frame[17] [1]), .O(n43386));
    defparam i3_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1251 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(n43117), .O(n26747));
    defparam i1_2_lut_3_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1252 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(n27078), .O(n42957));
    defparam i1_2_lut_3_lut_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_CARRY add_43_16 (.CI(n38217), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n38218));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1253 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(n42915), .O(n6_adj_4661));
    defparam i1_2_lut_3_lut_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1254 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[4] [7]), .O(n43318));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42991));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1256 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n27050), .I3(GND_net), .O(n43308));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1256.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_15_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n38216), .O(n2_adj_4477)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33733 (.I0(byte_transmit_counter[1]), 
            .I1(n46409), .I2(n46410), .I3(byte_transmit_counter[2]), .O(n48816));
    defparam byte_transmit_counter_1__bdd_4_lut_33733.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27103));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 n48816_bdd_4_lut (.I0(n48816), .I1(n46380), .I2(n46379), .I3(byte_transmit_counter[2]), 
            .O(n48819));
    defparam n48816_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1258 (.I0(n43308), .I1(Kp_23__N_1195), .I2(\data_in_frame[9] [1]), 
            .I3(n43465), .O(n10_adj_4613));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33728 (.I0(byte_transmit_counter[1]), 
            .I1(n46427), .I2(n46428), .I3(byte_transmit_counter[2]), .O(n48810));
    defparam byte_transmit_counter_1__bdd_4_lut_33728.LUT_INIT = 16'he4aa;
    SB_LUT4 n48810_bdd_4_lut (.I0(n48810), .I1(n46353), .I2(n46352), .I3(byte_transmit_counter[2]), 
            .O(n48813));
    defparam n48810_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42987));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(Kp_23__N_1195), .I1(n26730), .I2(GND_net), 
            .I3(GND_net), .O(n43468));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_CARRY add_43_15 (.CI(n38216), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n38217));
    SB_LUT4 add_43_14_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n38215), .O(n2_adj_4451)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33723 (.I0(byte_transmit_counter[1]), 
            .I1(n46433), .I2(n46434), .I3(byte_transmit_counter[2]), .O(n48804));
    defparam byte_transmit_counter_1__bdd_4_lut_33723.LUT_INIT = 16'he4aa;
    SB_LUT4 n48804_bdd_4_lut (.I0(n48804), .I1(n46344), .I2(n46343), .I3(byte_transmit_counter[2]), 
            .O(n48807));
    defparam n48804_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_14 (.CI(n38215), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n38216));
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_33718 (.I0(byte_transmit_counter[1]), 
            .I1(n46340), .I2(n46341), .I3(byte_transmit_counter[2]), .O(n48798));
    defparam byte_transmit_counter_1__bdd_4_lut_33718.LUT_INIT = 16'he4aa;
    SB_LUT4 n48798_bdd_4_lut (.I0(n48798), .I1(n46452), .I2(n46451), .I3(byte_transmit_counter[2]), 
            .O(n48801));
    defparam n48798_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_43_13_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n38214), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_4_lut_adj_1261 (.I0(\data_out_frame[5] [3]), .I1(n43318), 
            .I2(n43142), .I3(\data_out_frame[9] [5]), .O(n26656));
    defparam i2_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1262 (.I0(\data_out_frame[9] [4]), .I1(n43314), 
            .I2(n42991), .I3(\data_out_frame[5] [2]), .O(n26863));   // verilog/coms.v(73[16:34])
    defparam i3_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43042));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i15157_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n28668));
    defparam i15157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43502));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1265 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [3]), 
            .I2(n10_adj_4574), .I3(n41137), .O(n43148));
    defparam i5_3_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i15158_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n28669));
    defparam i15158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26504));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1306));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1267 (.I0(\data_out_frame[14] [0]), .I1(n26863), 
            .I2(n26656), .I3(\data_out_frame[11] [6]), .O(n27354));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(n26083), .I1(\data_out_frame[11] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n40238));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n28091));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15159_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n28670));
    defparam i15159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15160_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n28671));
    defparam i15160_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26662));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i15161_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n28672));
    defparam i15161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n28601));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1270 (.I0(n27354), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43183));
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(Kp_23__N_1195), .I1(n43520), .I2(GND_net), 
            .I3(GND_net), .O(n43114));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26599));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(n26730), .I1(n24669), .I2(GND_net), 
            .I3(GND_net), .O(n43126));
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1274 (.I0(n1510), .I1(n25928), .I2(n1513), 
            .I3(n27139), .O(n14_adj_4572));
    defparam i5_3_lut_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i15006_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n28517));
    defparam i15006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15007_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n28518));
    defparam i15007_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15008_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n28519));
    defparam i15008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(CLK_c), 
            .D(n7_adj_4663), .S(n42122));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15009_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n28520));
    defparam i15009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_13 (.CI(n38214), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n38215));
    SB_LUT4 i15010_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n28521));
    defparam i15010_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15011_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n28522));
    defparam i15011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(CLK_c), 
            .D(n7_adj_4664), .S(n42190));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(CLK_c), 
            .D(n42312), .S(n42204));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(CLK_c), 
            .D(n33802), .S(n42206));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(CLK_c), 
            .D(n42310), .S(n42208));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(CLK_c), 
            .D(n42308), .S(n42210));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(CLK_c), 
            .D(n42248), .S(n34417));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(CLK_c), 
            .D(n42306), .S(n42212));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(CLK_c), 
            .D(n7_adj_4665), .S(n8_adj_4666));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(CLK_c), 
            .D(n39601), .S(n42164));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(CLK_c), 
            .D(n42244), .S(n34415));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(CLK_c), 
            .D(n7_adj_4667), .S(n34413));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(CLK_c), 
            .D(n42304), .S(n42214));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(CLK_c), 
            .D(n7_adj_4668), .S(n34411));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(CLK_c), 
            .D(n42302), .S(n42216));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(CLK_c), 
            .D(n42298), .S(n42218));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(CLK_c), 
            .D(n7_adj_4459), .S(n42220));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(CLK_c), 
            .D(n42292), .S(n42222));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(CLK_c), 
            .D(n42286), .S(n42224));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(CLK_c), 
            .D(n42284), .S(n42226));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(CLK_c), 
            .D(n7_adj_4669), .S(n8_adj_4670));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(CLK_c), 
            .D(n42282), .S(n42182));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(CLK_c), 
            .D(n7_c), .S(n42228));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(CLK_c), 
            .D(n42276), .S(n42230));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(CLK_c), 
            .D(n42274), .S(n34409));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(CLK_c), 
            .D(n42272), .S(n42232));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(CLK_c), 
            .D(n42270), .S(n42176));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n42178), .S(n10_adj_4457));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1275 (.I0(n27469), .I1(n42918), .I2(n27296), 
            .I3(n43108), .O(n12_adj_4671));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1276 (.I0(n27262), .I1(n12_adj_4671), .I2(n27425), 
            .I3(\data_out_frame[13] [4]), .O(n26855));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i15012_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n28523));
    defparam i15012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15013_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n28524));
    defparam i15013_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n27804), .D(n44659));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43444));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1278 (.I0(n5_adj_4672), .I1(n43083), .I2(n43126), 
            .I3(n41086), .O(n14_adj_4673));
    defparam i6_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1279 (.I0(n26624), .I1(n14_adj_4673), .I2(n10_adj_4650), 
            .I3(n43114), .O(n25962));
    defparam i7_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1280 (.I0(n42963), .I1(n43296), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(Kp_23__N_1301));
    defparam i2_3_lut_adj_1280.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1281 (.I0(\data_in_frame[10] [3]), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[12] [5]), .I3(n24669), .O(n42949));
    defparam i2_3_lut_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i15144_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n28655));
    defparam i15144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15145_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n28656));
    defparam i15145_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15146_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n28657));
    defparam i15146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15147_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n28658));
    defparam i15147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1282 (.I0(n92[1]), .I1(n63), .I2(n4), .I3(n3813), 
            .O(n42174));   // verilog/coms.v(142[4] 144[7])
    defparam i1_3_lut_4_lut_adj_1282.LUT_INIT = 16'hbbb0;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(\data_out_frame[7] [1]), .I1(n43145), 
            .I2(n43281), .I3(n6_adj_4648), .O(n26083));   // verilog/coms.v(71[16:62])
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1284 (.I0(n41169), .I1(n27149), .I2(n4_adj_4609), 
            .I3(\data_in_frame[16] [2]), .O(n43508));
    defparam i1_2_lut_4_lut_adj_1284.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1285 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[8] [3]), .O(n6_adj_4569));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1286 (.I0(Kp_23__N_1301), .I1(n27377), .I2(n25962), 
            .I3(\data_in_frame[9] [0]), .O(n43222));
    defparam i3_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(n40699), .I1(n27149), .I2(GND_net), 
            .I3(GND_net), .O(n41096));
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1288 (.I0(tx_transmit_N_3513), .I1(n33792), 
            .I2(n26449), .I3(GND_net), .O(n4));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_1288.LUT_INIT = 16'h0e0e;
    SB_LUT4 i2_3_lut_adj_1289 (.I0(n43035), .I1(n43331), .I2(\data_in_frame[1] [3]), 
            .I3(GND_net), .O(n24669));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(n26755), .I1(n43222), .I2(GND_net), 
            .I3(GND_net), .O(n40205));
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i15148_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n28659));
    defparam i15148_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1291 (.I0(n43323), .I1(n43401), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[18] [2]), .O(n43353));
    defparam i1_2_lut_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1292 (.I0(\data_out_frame[16] [2]), .I1(n41182), 
            .I2(n27354), .I3(\data_out_frame[13] [7]), .O(n43484));
    defparam i2_3_lut_4_lut_adj_1292.LUT_INIT = 16'h9669;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n27804), .D(n26801));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n27804), .D(n44637));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n27804), .D(n43088));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n27804), .D(n44713));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15149_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n28660));
    defparam i15149_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n27804), .D(n27241));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n27804), .D(n41104));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n27804), .D(n44272));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n27804), .D(n45206));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n27804), .D(n44687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n27804), .D(n44073));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n27804), .D(n44066));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n27804), .D(n44071));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n27804), .D(n45100));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n27804), .D(n44663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n28600));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_12_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n38213), .O(n2_adj_4436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_12 (.CI(n38213), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n38214));
    SB_LUT4 i15152_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n28663));
    defparam i15152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_11_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n38212), .O(n2_adj_4501)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n38212), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n38213));
    SB_LUT4 i15153_3_lut_4_lut (.I0(n10_adj_4674), .I1(n42810), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n28664));
    defparam i15153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_10_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n38211), .O(n2_adj_4503)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n38211), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n38212));
    SB_LUT4 i2_2_lut_3_lut_adj_1293 (.I0(\data_in_frame[14] [4]), .I1(n43517), 
            .I2(n40922), .I3(GND_net), .O(n8_adj_4589));
    defparam i2_2_lut_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_9_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n38210), .O(n2_adj_4515)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n38210), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n38211));
    SB_LUT4 add_43_8_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n38209), .O(n2_adj_4528)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_8 (.CI(n38209), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n38210));
    SB_LUT4 i2_3_lut_4_lut_adj_1294 (.I0(\data_in_frame[14] [4]), .I1(n43517), 
            .I2(\data_in_frame[12] [3]), .I3(n44882), .O(n26744));
    defparam i2_3_lut_4_lut_adj_1294.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(Kp_23__N_1306), .I1(n43132), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n40336));
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42896));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26843));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1298 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [27]), .O(n42206));
    defparam i1_2_lut_3_lut_4_lut_adj_1298.LUT_INIT = 16'hf800;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [4]), .O(n1247));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1300 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [26]), .O(n42208));
    defparam i1_2_lut_3_lut_4_lut_adj_1300.LUT_INIT = 16'hf800;
    SB_LUT4 i2_3_lut_adj_1301 (.I0(n43311), .I1(n43468), .I2(\data_in_frame[13] [1]), 
            .I3(GND_net), .O(n42932));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1301.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1302 (.I0(n42932), .I1(n43520), .I2(n41086), 
            .I3(n43465), .O(n20_adj_4675));
    defparam i8_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1303 (.I0(n43374), .I1(\data_in_frame[13] [2]), 
            .I2(Kp_23__N_1301), .I3(n43502), .O(n19_adj_4676));
    defparam i7_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1304 (.I0(n4_adj_4609), .I1(n40205), .I2(n24669), 
            .I3(n41096), .O(n21));
    defparam i9_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut_4_lut (.I0(Kp_23__N_1306), .I1(n43132), .I2(n43474), 
            .I3(n42955), .O(n17_adj_4583));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1305 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42912));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1305.LUT_INIT = 16'h6666;
    SB_LUT4 i11_3_lut_adj_1306 (.I0(n21), .I1(n19_adj_4676), .I2(n20_adj_4675), 
            .I3(GND_net), .O(n41143));
    defparam i11_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i14990_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n28501));
    defparam i14990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1307 (.I0(tx_transmit_N_3513), .I1(n33792), 
            .I2(n23534), .I3(n26449), .O(n1));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut_adj_1307.LUT_INIT = 16'h00e0;
    SB_LUT4 i3_4_lut_adj_1308 (.I0(\data_in_frame[17] [5]), .I1(n42867), 
            .I2(\data_in_frame[15] [3]), .I3(n41143), .O(n40393));
    defparam i3_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1093), 
            .I2(GND_net), .I3(GND_net), .O(n27145));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i14991_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n28502));
    defparam i14991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n28090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n28599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n28598));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26717));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_7_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n38208), .O(n2_adj_4530)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n28597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n28596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n28595));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n42938), .I3(GND_net), .O(n27484));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_CARRY add_43_7 (.CI(n38208), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n38209));
    SB_LUT4 add_43_6_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n38207), .O(n2_adj_4531)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1312 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [25]), .O(n42210));
    defparam i1_2_lut_3_lut_4_lut_adj_1312.LUT_INIT = 16'hf800;
    SB_LUT4 i14992_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n28503));
    defparam i14992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1313 (.I0(\data_in_frame[6] [1]), .I1(Kp_23__N_936), 
            .I2(Kp_23__N_1090), .I3(\data_in_frame[6] [2]), .O(Kp_23__N_1186));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i20913_2_lut_3_lut_4_lut (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [24]), .O(n34417));
    defparam i20913_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut_adj_1314 (.I0(\data_out_frame[16] [4]), .I1(n26840), 
            .I2(\data_out_frame[18] [6]), .I3(\data_out_frame[16] [5]), 
            .O(n43209));
    defparam i1_2_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_out_frame[8] [5]), .I1(n1247), 
            .I2(GND_net), .I3(GND_net), .O(n27360));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i14993_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n28504));
    defparam i14993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n28089));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14994_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n28505));
    defparam i14994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14995_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n28506));
    defparam i14995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1316 (.I0(\data_out_frame[20] [6]), .I1(n26676), 
            .I2(n10_adj_4574), .I3(n41137), .O(n41204));
    defparam i1_2_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1317 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [23]), .O(n42212));
    defparam i1_2_lut_3_lut_4_lut_adj_1317.LUT_INIT = 16'hf800;
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n28088));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_1186), 
            .I2(GND_net), .I3(GND_net), .O(n27152));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1319 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [22]), .O(n8_adj_4666));
    defparam i1_2_lut_3_lut_4_lut_adj_1319.LUT_INIT = 16'hf800;
    SB_LUT4 i14996_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n28507));
    defparam i14996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42915));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1321 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n43011));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1321.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27186));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1323 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [21]), .O(n42164));
    defparam i1_2_lut_3_lut_4_lut_adj_1323.LUT_INIT = 16'hf800;
    SB_LUT4 i4_4_lut_adj_1324 (.I0(n27403), .I1(Kp_23__N_936), .I2(n27186), 
            .I3(n6_adj_4661), .O(n26730));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1325 (.I0(\data_in_frame[5] [1]), .I1(n43120), 
            .I2(\data_in_frame[7] [2]), .I3(GND_net), .O(n27149));
    defparam i2_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i20912_2_lut_3_lut_4_lut (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [20]), .O(n34415));
    defparam i20912_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i2_3_lut_adj_1326 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n27500));
    defparam i2_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1327 (.I0(n26449), .I1(\FRAME_MATCHER.i_31__N_2622 ), 
            .I2(tx_active), .I3(r_SM_Main_2__N_3616[0]), .O(n27621));
    defparam i1_3_lut_4_lut_adj_1327.LUT_INIT = 16'hcccd;
    SB_LUT4 i14997_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n28508));
    defparam i14997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1328 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [19]), .O(n34413));
    defparam i1_2_lut_3_lut_4_lut_adj_1328.LUT_INIT = 16'hf800;
    SB_LUT4 i5_3_lut_4_lut_adj_1329 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[6] [0]), .O(n14_adj_4551));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_CARRY add_43_6 (.CI(n38207), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n38208));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1330 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [18]), .O(n42214));
    defparam i1_2_lut_3_lut_4_lut_adj_1330.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[20] [0]), 
            .I2(n40935), .I3(GND_net), .O(n43197));
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_5_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n38206), .O(n2_adj_4532)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n38206), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n38207));
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42902));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1333 (.I0(n43080), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[20] [2]), .I3(\data_out_frame[20] [3]), 
            .O(n27090));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i15136_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n28647));
    defparam i15136_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15137_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n28648));
    defparam i15137_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_4_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n38205), .O(n2_adj_4533)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15138_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n28649));
    defparam i15138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_4 (.CI(n38205), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n38206));
    SB_LUT4 i15139_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n28650));
    defparam i15139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15140_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n28651));
    defparam i15140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15141_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n28652));
    defparam i15141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15142_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n28653));
    defparam i15142_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1334 (.I0(n26855), .I1(n43183), .I2(n4_adj_4656), 
            .I3(n40238), .O(n43401));
    defparam i2_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_3_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n38204), .O(n2_adj_4537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_3 (.CI(n38204), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n38205));
    SB_LUT4 add_43_2_lut (.I0(n3065), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_4487)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1335 (.I0(n43055), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[7] [4]), .I3(n43350), .O(n10_adj_4677));
    defparam i4_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n38204));
    SB_LUT4 i5_3_lut_adj_1336 (.I0(n27253), .I1(n10_adj_4677), .I2(n27500), 
            .I3(GND_net), .O(n26755));
    defparam i5_3_lut_adj_1336.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1337 (.I0(\data_out_frame[20] [0]), .I1(n43080), 
            .I2(n43365), .I3(\data_out_frame[20] [3]), .O(n43154));
    defparam i1_2_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i15143_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n28654));
    defparam i15143_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\data_in_frame[5] [3]), .I1(n26905), 
            .I2(GND_net), .I3(GND_net), .O(n43055));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1339 (.I0(n44105), .I1(\data_in_frame[18] [5]), 
            .I2(n40393), .I3(\data_in_frame[16] [3]), .O(n43008));
    defparam i2_3_lut_4_lut_adj_1339.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [1]), 
            .I2(n25950), .I3(GND_net), .O(n43450));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i20910_2_lut_3_lut_4_lut (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [17]), .O(n34411));
    defparam i20910_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i3_4_lut_adj_1341 (.I0(\data_in_frame[5] [4]), .I1(n43426), 
            .I2(n43347), .I3(n27078), .O(n40225));
    defparam i3_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1342 (.I0(n44105), .I1(\data_in_frame[18] [5]), 
            .I2(n43480), .I3(\data_in_frame[16] [4]), .O(n8_adj_4678));
    defparam i3_3_lut_4_lut_adj_1342.LUT_INIT = 16'h9669;
    SB_LUT4 i14982_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n28493));
    defparam i14982_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14983_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n28494));
    defparam i14983_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_in_frame[4] [7]), .I1(n27500), 
            .I2(GND_net), .I3(GND_net), .O(n42928));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i14984_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n28495));
    defparam i14984_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14985_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n28496));
    defparam i14985_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14986_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n28497));
    defparam i14986_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14987_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n28498));
    defparam i14987_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14988_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n28499));
    defparam i14988_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14989_3_lut_4_lut (.I0(n34442), .I1(n42838), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n28500));
    defparam i14989_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14974_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n28485));
    defparam i14974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14975_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n28486));
    defparam i14975_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14976_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n28487));
    defparam i14976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14977_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n28488));
    defparam i14977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n28594));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14978_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n28489));
    defparam i14978_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14979_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n28490));
    defparam i14979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14980_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n28491));
    defparam i14980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1344 (.I0(n4_adj_4647), .I1(n25928), .I2(n43142), 
            .I3(\data_out_frame[14] [2]), .O(n14_adj_4679));
    defparam i6_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i14981_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42832), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n28492));
    defparam i14981_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1345 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[5] [5]), .O(n43462));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1345.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1346 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[8] [2]), .I3(n43423), .O(n42984));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i14966_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n28477));
    defparam i14966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14967_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n28478));
    defparam i14967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14968_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n28479));
    defparam i14968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15162_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n28673));
    defparam i15162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14969_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n28480));
    defparam i14969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14970_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n28481));
    defparam i14970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1347 (.I0(\data_in_frame[4] [6]), .I1(n27072), 
            .I2(n27062), .I3(\data_in_frame[7] [0]), .O(n43099));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1348 (.I0(\data_in_frame[6] [7]), .I1(n43099), 
            .I2(n26580), .I3(\data_in_frame[6] [6]), .O(n26702));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1349 (.I0(\data_in_frame[7] [3]), .I1(n42952), 
            .I2(n26905), .I3(n27059), .O(n40699));
    defparam i3_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i14971_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n28482));
    defparam i14971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1350 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [12]), .O(n42224));
    defparam i1_2_lut_3_lut_4_lut_adj_1350.LUT_INIT = 16'hf800;
    SB_LUT4 i14972_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n28483));
    defparam i14972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14973_3_lut_4_lut (.I0(n8_adj_4590), .I1(n42832), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n28484));
    defparam i14973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1351 (.I0(\data_out_frame[9] [1]), .I1(n10_adj_4602), 
            .I2(n27139), .I3(\data_out_frame[13] [0]), .O(n43493));
    defparam i1_2_lut_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1352 (.I0(\data_out_frame[9] [1]), .I1(n10_adj_4602), 
            .I2(n27139), .I3(n26855), .O(n43407));
    defparam i1_2_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i14958_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n28469));
    defparam i14958_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n28593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n28592));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n28591));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n28590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n28589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n28587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n28586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n28585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n28584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n28583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n28582));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n28581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n28580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n28579));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n28578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n28546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n28545));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n28544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n28543));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14959_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n28470));
    defparam i14959_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14960_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n28471));
    defparam i14960_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14961_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n28472));
    defparam i14961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n28535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n28534));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14962_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n28473));
    defparam i14962_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n28533));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n28532));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14963_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n28474));
    defparam i14963_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n28531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n28530));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14964_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n28475));
    defparam i14964_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n28528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n28527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n28526));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14965_3_lut_4_lut (.I0(n10_adj_4615), .I1(n42810), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n28476));
    defparam i14965_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n28525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n28524));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [5]), 
            .I2(n27047), .I3(GND_net), .O(n43225));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n28523));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1354 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [5]), 
            .I2(n26504), .I3(n10_adj_4568), .O(n43031));
    defparam i5_3_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n28522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n28521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n28520));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14950_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n28461));
    defparam i14950_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n28519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n28518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n28517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n28516));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1355 (.I0(\data_out_frame[7] [5]), .I1(n14_adj_4679), 
            .I2(n10_adj_4646), .I3(n26863), .O(n26840));
    defparam i7_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n28515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n28514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n28513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n28512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n28511));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14951_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n28462));
    defparam i14951_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n28510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n28509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n28508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n28507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n28506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n28505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n28504));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14952_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n28463));
    defparam i14952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n28503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n28502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n28501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n28500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n28499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n28498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n28497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n28496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n28495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n28494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n28493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n28492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n28491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n28490));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14953_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n28464));
    defparam i14953_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n28489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n28488));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15163_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n28674));
    defparam i15163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n28487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n28486));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n28485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n28484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n28483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n28482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n28481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n28480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n28479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n28478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n28477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n28476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n28475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n28474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n28473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n28472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n28471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n28470));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14954_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n28465));
    defparam i14954_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n28469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n28468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n28467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n28466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n28465));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n28464));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_2186_i5_2_lut (.I0(Kp_23__N_1189), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4672));   // verilog/coms.v(236[9:81])
    defparam equal_2186_i5_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n28463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n28462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n28461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n28460));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n28459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n28458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n28457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n28456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n28455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n28454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n28453));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n28452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n28451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n28450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n28449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n28448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n28447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n28446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n28445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n28438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n28437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n28433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n28432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n28431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n28430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n28429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n28428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n28426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n28425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n28424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n28423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n28422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n28421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n28420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n28416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n28415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n28414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n28413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n28412));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14955_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n28466));
    defparam i14955_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1356 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[1] [7]), 
            .I2(n27062), .I3(n6_adj_4581), .O(Kp_23__N_1099));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i15164_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n28675));
    defparam i15164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14956_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n28467));
    defparam i14956_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1357 (.I0(n26840), .I1(n43401), .I2(n42921), 
            .I3(n27360), .O(n28));
    defparam i10_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1358 (.I0(n26599), .I1(n43275), .I2(n42884), 
            .I3(\data_in_frame[2] [0]), .O(Kp_23__N_1096));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1359 (.I0(Kp_23__N_1099), .I1(n27072), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n42995));
    defparam i2_3_lut_adj_1359.LUT_INIT = 16'h9696;
    SB_LUT4 i15165_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n28676));
    defparam i15165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1360 (.I0(n26593), .I1(n27062), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n27258));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i14957_3_lut_4_lut (.I0(n8_adj_4652), .I1(n42832), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n28468));
    defparam i14957_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1361 (.I0(\data_in_frame[6] [0]), .I1(n42899), 
            .I2(n40197), .I3(n27258), .O(n42955));
    defparam i3_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i15166_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n28677));
    defparam i15166_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43245));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1363 (.I0(\data_in_frame[1] [4]), .I1(n43245), 
            .I2(n42955), .I3(n43028), .O(n41086));
    defparam i3_4_lut_adj_1363.LUT_INIT = 16'h9669;
    SB_LUT4 i15167_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n28678));
    defparam i15167_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14942_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n28453));
    defparam i14942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14943_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n28454));
    defparam i14943_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15168_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n28679));
    defparam i15168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_3_lut (.I0(\data_out_frame[14] [6]), .I1(n28), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n32_adj_4680));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14944_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n28455));
    defparam i14944_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14945_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n28456));
    defparam i14945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n28411));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14946_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n28457));
    defparam i14946_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1364 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [11]), .O(n42226));
    defparam i1_2_lut_3_lut_4_lut_adj_1364.LUT_INIT = 16'hf800;
    SB_LUT4 i3_4_lut_adj_1365 (.I0(\data_in_frame[4] [0]), .I1(n43272), 
            .I2(n42884), .I3(\data_in_frame[1] [4]), .O(Kp_23__N_1090));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i14947_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n28458));
    defparam i14947_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14948_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n28459));
    defparam i14948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14949_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42832), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n28460));
    defparam i14949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1366 (.I0(\data_out_frame[14] [7]), .I1(n43015), 
            .I2(n43493), .I3(n42938), .O(n30));
    defparam i12_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1367 (.I0(n26950), .I1(\data_out_frame[16] [7]), 
            .I2(n27484), .I3(n43441), .O(n8_adj_4538));
    defparam i3_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1368 (.I0(n26604), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [1]), .I3(n6_adj_4582), .O(Kp_23__N_1093));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [10]), .O(n8_adj_4670));
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[8] [4]), .I3(GND_net), .O(n43423));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1371 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(n26456), .I3(\data_out_frame[10] [7]), .O(n8_adj_4594));   // verilog/coms.v(74[16:43])
    defparam i3_3_lut_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1372 (.I0(n42864), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [6]), .I3(n27031), .O(n31_adj_4681));
    defparam i13_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i14636_3_lut_4_lut (.I0(n8_adj_4471), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n28147));
    defparam i14636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(n23743), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n36539), .I3(GND_net), .O(n110));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1374 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43238));
    defparam i1_2_lut_adj_1374.LUT_INIT = 16'h6666;
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n28410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n28409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n28408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n28407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n28406));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15128_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n28639));
    defparam i15128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n28405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n28404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n28403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n28402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n28401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n28400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n28399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n28398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n28397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n28396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n28395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n28394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n28393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n28392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n28391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n28390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n28389));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(\data_out_frame[18] [1]), .I1(n41090), 
            .I2(\data_out_frame[20] [2]), .I3(n45249), .O(n40257));
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'h9669;
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n28388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n28387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n28386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n28385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n28384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n28383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n28382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n28381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n28380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n28379));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n28378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n28377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n28373));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1376 (.I0(\data_out_frame[18] [1]), .I1(n41090), 
            .I2(\data_out_frame[20] [3]), .I3(n43353), .O(n45042));
    defparam i2_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i15129_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n28640));
    defparam i15129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1377 (.I0(\data_in_frame[1] [0]), .I1(n42960), 
            .I2(GND_net), .I3(GND_net), .O(n26637));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1377.LUT_INIT = 16'h6666;
    SB_LUT4 i15130_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n28641));
    defparam i15130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n28361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n28360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n28359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n28358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n28357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n28356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n28355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n28354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n28353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n28352));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15131_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n28642));
    defparam i15131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n28351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n28350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n28349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n28348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n28347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n28346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n28345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n28344));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15132_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n28643));
    defparam i15132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n28343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n28342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n28341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n28340));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15133_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n28644));
    defparam i15133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n28339));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n28338));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15134_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n28645));
    defparam i15134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n28337));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1378 (.I0(n27357), .I1(n27522), .I2(n42984), 
            .I3(n27326), .O(n29));
    defparam i11_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n28336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n28335));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15135_3_lut_4_lut (.I0(n8_adj_4662), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n28646));
    defparam i15135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n28329));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43284));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n28328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n28327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n28326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n28325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n28324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n28323));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_299_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4662));   // verilog/coms.v(154[7:23])
    defparam equal_299_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n28322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n28321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n28320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n28319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n28318));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1380 (.I0(n43284), .I1(n27253), .I2(\data_in_frame[2] [5]), 
            .I3(n42896), .O(n10_adj_4580));   // verilog/coms.v(166[9:87])
    defparam i4_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n28317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n28316));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n28315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n28314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n28313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n28312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n28311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n28310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n28309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n28308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n28307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n28306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n28305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n28304));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n28303));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n28302));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n28301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n28300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n28299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n28298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n28297));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1381 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42816), .I3(\FRAME_MATCHER.i [0]), .O(n42822));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1381.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n28296));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n28295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n28294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n28293));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n28292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n28291));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n28290));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n28289));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n28288));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n28287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n28286));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1382 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42884));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1382.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1383 (.I0(\data_in_frame[1] [4]), .I1(n26667), 
            .I2(n26604), .I3(\data_in_frame[1] [3]), .O(n42960));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1384 (.I0(n42960), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n43347));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1385 (.I0(\data_in_frame[4] [4]), .I1(n26599), 
            .I2(GND_net), .I3(GND_net), .O(n43447));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1385.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n28285));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n28284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n28283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n28282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n28281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n28280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n28279));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n28278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n28277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n28276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n28275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n28274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n28273));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n28272));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n28271));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n28270));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1386 (.I0(\FRAME_MATCHER.state [1]), .I1(n29908), 
            .I2(n21657), .I3(n4452), .O(n2_adj_4682));
    defparam i1_3_lut_4_lut_adj_1386.LUT_INIT = 16'h0080;
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n28269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n28268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n28267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n28266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n28262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n28261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n28260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n28258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n28257));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1387 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42832), .I3(\FRAME_MATCHER.i [0]), .O(n42836));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1387.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n28256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n28255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n28254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n28253));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i17_4_lut_adj_1388 (.I0(n29), .I1(n31_adj_4681), .I2(n30), 
            .I3(n32_adj_4680), .O(n44237));
    defparam i17_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(n3065), .I1(n161), .I2(n10_adj_4615), 
            .I3(GND_net), .O(n42832));
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'hf7f7;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n28252));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n28251));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1390 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42838), .I3(\FRAME_MATCHER.i [0]), .O(n42843));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1390.LUT_INIT = 16'hfbff;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n28250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n28249));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1391 (.I0(n3065), .I1(n161), .I2(n10_adj_4593), 
            .I3(GND_net), .O(n42838));
    defparam i1_2_lut_3_lut_adj_1391.LUT_INIT = 16'hf7f7;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n28248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n28247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n28246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n28245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n28243));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1392 (.I0(\data_in_frame[0] [7]), .I1(n43042), 
            .I2(n42912), .I3(n42902), .O(Kp_23__N_969));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n28242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n28241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n28240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n28239));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1393 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(n10_adj_4536), .I3(n43417), .O(n43441));
    defparam i5_3_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n28087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n28238));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1394 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[4] [0]), .O(n43102));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1395 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(\data_out_frame[15] [0]), 
            .O(n43395));
    defparam i2_3_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1396 (.I0(\data_in_frame[5] [1]), .I1(n43347), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n42952));
    defparam i2_3_lut_adj_1396.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n28237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n28236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n28235));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1397 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26915));
    defparam i2_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1398 (.I0(\data_out_frame[15] [6]), .I1(n40326), 
            .I2(\data_out_frame[16] [1]), .I3(\data_out_frame[16] [0]), 
            .O(n43323));
    defparam i2_3_lut_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1399 (.I0(\data_out_frame[15] [6]), .I1(n40326), 
            .I2(\data_out_frame[17] [7]), .I3(\data_out_frame[18] [0]), 
            .O(n43514));
    defparam i2_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1400 (.I0(n3065), .I1(n161), .I2(\FRAME_MATCHER.i [0]), 
            .I3(n7_adj_4645), .O(n42810));
    defparam i2_3_lut_4_lut_adj_1400.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1401 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [9]), .O(n42182));
    defparam i1_2_lut_3_lut_4_lut_adj_1401.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(n3065), .I1(n161), .I2(n10_adj_4674), 
            .I3(GND_net), .O(n42816));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1403 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [8]), .O(n42228));
    defparam i1_2_lut_3_lut_4_lut_adj_1403.LUT_INIT = 16'hf800;
    SB_LUT4 equal_296_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4593));   // verilog/coms.v(154[7:23])
    defparam equal_296_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26667));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1405 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43028));
    defparam i1_2_lut_adj_1405.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\data_out_frame[9] [1]), .I1(n26915), 
            .I2(GND_net), .I3(GND_net), .O(n42918));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1407 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [7]), .O(n42230));
    defparam i1_2_lut_3_lut_4_lut_adj_1407.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43177));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 equal_304_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4674));   // verilog/coms.v(154[7:23])
    defparam equal_304_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1409 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[3] [6]), .O(n43272));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1410 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43275));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(\data_out_frame[4] [7]), .I1(n43111), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4683));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1412 (.I0(n27072), .I1(n42952), .I2(n43102), 
            .I3(Kp_23__N_969), .O(n24_adj_4684));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1413 (.I0(n43272), .I1(n42957), .I2(n27403), 
            .I3(\data_in_frame[3] [5]), .O(n22_adj_4685));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1414 (.I0(n43120), .I1(n24_adj_4684), .I2(n18_adj_4642), 
            .I3(\data_in_frame[2] [1]), .O(n26_adj_4686));   // verilog/coms.v(74[16:43])
    defparam i12_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1415 (.I0(n26545), .I1(n26_adj_4686), .I2(n22_adj_4685), 
            .I3(\data_in_frame[4] [7]), .O(n40197));   // verilog/coms.v(74[16:43])
    defparam i13_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1416 (.I0(Kp_23__N_1093), .I1(Kp_23__N_1090), .I2(GND_net), 
            .I3(GND_net), .O(n42981));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1416.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1417 (.I0(n2134), .I1(n41177), .I2(\data_out_frame[24] [0]), 
            .I3(\data_out_frame[23] [5]), .O(n6_adj_4441));
    defparam i1_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1418 (.I0(\data_in_frame[6] [7]), .I1(n43523), 
            .I2(\data_in_frame[6] [1]), .I3(n26717), .O(n42899));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1419 (.I0(n2134), .I1(n41177), .I2(\data_out_frame[24] [0]), 
            .I3(n43438), .O(n6_adj_4442));
    defparam i1_2_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1420 (.I0(n42899), .I1(n42981), .I2(n40197), 
            .I3(\data_in_frame[8] [1]), .O(n12_adj_4687));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1421 (.I0(n1168), .I1(\data_out_frame[7] [1]), 
            .I2(n42918), .I3(n6_adj_4683), .O(n27469));   // verilog/coms.v(71[16:69])
    defparam i4_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1422 (.I0(Kp_23__N_936), .I1(n12_adj_4687), .I2(n42995), 
            .I3(Kp_23__N_1096), .O(n44479));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1423 (.I0(n41086), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n41145));
    defparam i1_2_lut_adj_1423.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1424 (.I0(n41145), .I1(n40699), .I2(n26702), 
            .I3(n44479), .O(n16_adj_4688));
    defparam i6_4_lut_adj_1424.LUT_INIT = 16'hfff7;
    SB_LUT4 i7_4_lut_adj_1425 (.I0(n13), .I1(n40225), .I2(n40294), .I3(\data_in_frame[7] [7]), 
            .O(n17_adj_4689));
    defparam i7_4_lut_adj_1425.LUT_INIT = 16'hfeef;
    SB_LUT4 i9_4_lut_adj_1426 (.I0(n17_adj_4689), .I1(n26747), .I2(n16_adj_4688), 
            .I3(n26755), .O(n45310));
    defparam i9_4_lut_adj_1426.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_4_lut_adj_1427 (.I0(n45310), .I1(n4_adj_4609), .I2(n27149), 
            .I3(n26730), .O(n12_adj_4690));
    defparam i5_4_lut_adj_1427.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1428 (.I0(\data_out_frame[5] [4]), .I1(n42921), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n43281));   // verilog/coms.v(71[16:62])
    defparam i2_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1429 (.I0(n27377), .I1(n12_adj_4690), .I2(n27152), 
            .I3(n8_adj_4607), .O(n31));
    defparam i6_4_lut_adj_1429.LUT_INIT = 16'hfffe;
    SB_LUT4 i20909_2_lut_3_lut_4_lut (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [6]), .O(n34409));
    defparam i20909_2_lut_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i3_3_lut_adj_1430 (.I0(n40393), .I1(\data_in_frame[19] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n8_adj_4691));
    defparam i3_3_lut_adj_1430.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1431 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [5]), .O(n42232));
    defparam i1_2_lut_3_lut_4_lut_adj_1431.LUT_INIT = 16'hf800;
    SB_LUT4 i2_4_lut_adj_1432 (.I0(\data_in_frame[19] [3]), .I1(n43386), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[21] [4]), .O(n44982));
    defparam i2_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1433 (.I0(n41184), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[21] [6]), .I3(\data_in_frame[19] [5]), .O(n44432));
    defparam i2_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1434 (.I0(n21657), .I1(n3813), .I2(n42849), 
            .I3(\FRAME_MATCHER.state_c [4]), .O(n42176));
    defparam i1_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'hf800;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(76[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1435 (.I0(n41117), .I1(n43093), .I2(\data_in_frame[19] [7]), 
            .I3(\data_in_frame[20] [1]), .O(n44899));
    defparam i3_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i15098_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n28609));
    defparam i15098_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15099_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n28610));
    defparam i15099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1436 (.I0(\data_in_frame[21] [5]), .I1(n41188), 
            .I2(\data_in_frame[19] [4]), .I3(n6_adj_4640), .O(n45108));
    defparam i4_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i15100_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n28611));
    defparam i15100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1437 (.I0(n43008), .I1(\data_in_frame[19] [0]), 
            .I2(\data_in_frame[16] [4]), .I3(n43241), .O(n10_adj_4692));
    defparam i4_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1438 (.I0(\data_in_frame[20] [3]), .I1(n43174), 
            .I2(n40675), .I3(\data_in_frame[18] [1]), .O(n44441));
    defparam i3_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1439 (.I0(\data_in_frame[21] [1]), .I1(n43487), 
            .I2(n43202), .I3(n41184), .O(n44205));
    defparam i3_4_lut_adj_1439.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1440 (.I0(n40284), .I1(n43487), .I2(n41184), 
            .I3(\data_in_frame[21] [0]), .O(n44203));
    defparam i3_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i15113_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n28624));
    defparam i15113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21117_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n34624), .I2(GND_net), 
            .I3(GND_net), .O(n34626));
    defparam i21117_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15114_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n28625));
    defparam i15114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1441 (.I0(n41169), .I1(n10_adj_4692), .I2(\data_in_frame[20] [7]), 
            .I3(GND_net), .O(n44641));
    defparam i5_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i1_rep_99_2_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n49063));   // verilog/coms.v(85[17:28])
    defparam i1_rep_99_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1442 (.I0(n43093), .I1(n43371), .I2(n41117), 
            .I3(n49063), .O(n12_adj_4693));
    defparam i5_4_lut_adj_1442.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1443 (.I0(\data_out_frame[6] [6]), .I1(n43145), 
            .I2(\data_out_frame[9] [2]), .I3(n1130), .O(n43111));
    defparam i3_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1444 (.I0(\data_in_frame[20] [0]), .I1(n12_adj_4693), 
            .I2(n43432), .I3(n41122), .O(n44064));
    defparam i6_4_lut_adj_1444.LUT_INIT = 16'h9669;
    SB_LUT4 i15115_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n28626));
    defparam i15115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1445 (.I0(\data_in_frame[16] [3]), .I1(n43031), 
            .I2(n43511), .I3(GND_net), .O(n8_adj_4694));
    defparam i3_3_lut_adj_1445.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1446 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[19] [1]), 
            .I2(n26050), .I3(n6_adj_4639), .O(n44594));
    defparam i4_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i15116_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n28627));
    defparam i15116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1447 (.I0(n44982), .I1(\data_in_frame[21] [7]), 
            .I2(n8_adj_4691), .I3(n27174), .O(n20_adj_4695));
    defparam i4_4_lut_adj_1447.LUT_INIT = 16'hbeeb;
    SB_LUT4 i15117_3_lut_4_lut (.I0(n8_adj_4651), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n28628));
    defparam i15117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1448 (.I0(n5_adj_4641), .I1(n44432), .I2(n43432), 
            .I3(n40675), .O(n18_adj_4696));
    defparam i2_4_lut_adj_1448.LUT_INIT = 16'hb77b;
    SB_LUT4 i3_4_lut_adj_1449 (.I0(n44899), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[21] [2]), .I3(n40284), .O(n19_adj_4697));
    defparam i3_4_lut_adj_1449.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_3_lut_adj_1450 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n43314));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1451 (.I0(\data_in_frame[20] [5]), .I1(n44594), 
            .I2(n8_adj_4694), .I3(n43508), .O(n17_adj_4698));
    defparam i1_4_lut_adj_1451.LUT_INIT = 16'hb77b;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(\data_out_frame[5] [1]), .I1(n43314), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4699));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1453 (.I0(\data_in_frame[20] [6]), .I1(n45108), 
            .I2(n8_adj_4678), .I3(n43511), .O(n22_adj_4700));
    defparam i6_4_lut_adj_1453.LUT_INIT = 16'hdeed;
    SB_LUT4 i12_4_lut_adj_1454 (.I0(n44641), .I1(n44203), .I2(n44205), 
            .I3(n44441), .O(n28_adj_4701));
    defparam i12_4_lut_adj_1454.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_4_lut_adj_1455 (.I0(n44064), .I1(n43031), .I2(n43174), 
            .I3(\data_in_frame[20] [4]), .O(n21_adj_4702));
    defparam i5_4_lut_adj_1455.LUT_INIT = 16'hd77d;
    SB_LUT4 i2_3_lut_4_lut_adj_1456 (.I0(\FRAME_MATCHER.state [0]), .I1(n36539), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [3]), 
            .O(n29908));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1456.LUT_INIT = 16'h0002;
    SB_LUT4 i13_4_lut_adj_1457 (.I0(n17_adj_4698), .I1(n19_adj_4697), .I2(n18_adj_4696), 
            .I3(n20_adj_4695), .O(n29_adj_4703));
    defparam i13_4_lut_adj_1457.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1458 (.I0(n29_adj_4703), .I1(n21_adj_4702), .I2(n28_adj_4701), 
            .I3(n22_adj_4700), .O(n3_adj_4439));
    defparam i15_4_lut_adj_1458.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1459 (.I0(\data_out_frame[9] [3]), .I1(n27421), 
            .I2(n43111), .I3(n6_adj_4699), .O(n24464));
    defparam i4_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\FRAME_MATCHER.state [0]), .I1(n36539), 
            .I2(n130), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2624 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h2020;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(\data_out_frame[8] [7]), .I1(n27469), 
            .I2(GND_net), .I3(GND_net), .O(n43180));
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26860));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1463 (.I0(n23743), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n7001));
    defparam i2_3_lut_adj_1463.LUT_INIT = 16'h1010;
    SB_LUT4 i3_4_lut_adj_1464 (.I0(\data_out_frame[13] [5]), .I1(n26860), 
            .I2(n43180), .I3(n24464), .O(n40326));
    defparam i3_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n6_adj_4445));
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43071));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1467 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [4]), .I3(\data_out_frame[15] [2]), 
            .O(n42978));
    defparam i2_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1468 (.I0(\FRAME_MATCHER.state [2]), .I1(n3_adj_4439), 
            .I2(n31), .I3(\FRAME_MATCHER.state [1]), .O(n6_adj_4704));
    defparam i2_4_lut_adj_1468.LUT_INIT = 16'h0a22;
    SB_LUT4 i3_4_lut_adj_1469 (.I0(n34377), .I1(n6_adj_4704), .I2(n23743), 
            .I3(n43606), .O(n27605));
    defparam i3_4_lut_adj_1469.LUT_INIT = 16'h0004;
    SB_LUT4 mux_2022_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7002));
    defparam mux_2022_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31195_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n46275), .I3(n20_adj_4546), .O(n46276));
    defparam i31195_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i5_4_lut_adj_1470 (.I0(\data_out_frame[6] [0]), .I1(n43071), 
            .I2(\data_out_frame[8] [1]), .I3(\data_out_frame[5] [7]), .O(n12_adj_4705));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i31375_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n46455), .I3(n20_adj_4548), .O(n46456));
    defparam i31375_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i31366_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n46446), .I3(n20_adj_4552), .O(n46447));
    defparam i31366_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i15089_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n28600));
    defparam i15089_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15090_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n28601));
    defparam i15090_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1471 (.I0(\data_out_frame[7] [5]), .I1(n12_adj_4705), 
            .I2(n43359), .I3(\data_out_frame[10] [1]), .O(n1513));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i15091_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n28602));
    defparam i15091_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15092_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n28603));
    defparam i15092_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i31222_3_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(n46302), .O(n46303));   // verilog/coms.v(106[34:55])
    defparam i31222_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 i15093_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n28604));
    defparam i15093_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i31164_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n29908), 
            .I2(n21657), .I3(n771), .O(n46187));   // verilog/coms.v(115[11:12])
    defparam i31164_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i7_2_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4706));
    defparam i7_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(Kp_23__N_969), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n24791));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27306));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i31201_3_lut_4_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(n46281), .O(n46282));   // verilog/coms.v(106[34:55])
    defparam i31201_3_lut_4_lut.LUT_INIT = 16'hf202;
    SB_LUT4 i15095_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n28606));
    defparam i15095_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15096_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n28607));
    defparam i15096_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15097_3_lut_4_lut (.I0(n34442), .I1(n42816), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n28608));
    defparam i15097_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1474 (.I0(\data_in_frame[2] [0]), .I1(n23743), 
            .I2(n42941), .I3(n24791), .O(n26_adj_4707));
    defparam i9_4_lut_adj_1474.LUT_INIT = 16'h2100;
    SB_LUT4 i1_3_lut_4_lut_adj_1475 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n26350), .I3(\FRAME_MATCHER.i [1]), .O(n5_c));
    defparam i1_3_lut_4_lut_adj_1475.LUT_INIT = 16'hfefc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46303), .I3(n46301), .O(n7_adj_4547));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1476 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43235));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1476.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_4_lut_adj_1477 (.I0(n42854), .I1(n4_adj_4535), .I2(n53), 
            .I3(n133), .O(n8));   // verilog/coms.v(127[12] 300[6])
    defparam i3_3_lut_4_lut_adj_1477.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(GND_net), .I3(GND_net), .O(n26491));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1479 (.I0(\data_in_frame[1] [7]), .I1(n24_adj_4706), 
            .I2(\data_in_frame[1] [6]), .I3(n42941), .O(n29_adj_4708));
    defparam i12_4_lut_adj_1479.LUT_INIT = 16'h4080;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n43608), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'h0404;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46294), .I3(n46292), .O(n7_adj_4549));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1481 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n34624), .I3(GND_net), .O(n27804));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1481.LUT_INIT = 16'h0404;
    SB_LUT4 i31124_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [7]), 
            .I2(n42902), .I3(\data_in_frame[1] [1]), .O(n46147));
    defparam i31124_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i5_4_lut_adj_1482 (.I0(\data_out_frame[8] [0]), .I1(n43235), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[5] [4]), .O(n12_adj_4709));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1483 (.I0(\data_out_frame[6] [1]), .I1(n12_adj_4709), 
            .I2(n43359), .I3(\data_out_frame[4] [0]), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1484 (.I0(n1516), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [5]), .I3(n26491), .O(n27357));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1485 (.I0(\data_out_frame[23] [1]), .I1(n41137), 
            .I2(\data_out_frame[20] [6]), .I3(n10_adj_4539), .O(n40210));
    defparam i5_3_lut_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\data_out_frame[15] [0]), .I1(n27357), 
            .I2(GND_net), .I3(GND_net), .O(n43206));
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1487 (.I0(n26593), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [2]), .I3(n42907), .O(n28_adj_4710));
    defparam i11_4_lut_adj_1487.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(n44237), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43414));
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(\data_out_frame[15] [1]), .I1(n43414), 
            .I2(n43206), .I3(\data_out_frame[15] [6]), .O(n44005));
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26676));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46288), .I3(n46286), .O(n7_adj_4553));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_3_lut_4_lut_adj_1491 (.I0(\FRAME_MATCHER.state [3]), .I1(n21657), 
            .I2(n3813), .I3(n2_adj_4682), .O(n42178));
    defparam i1_3_lut_4_lut_adj_1491.LUT_INIT = 16'haa80;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46327), .I3(n46325), .O(n7_adj_4601));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_4_lut_adj_1492 (.I0(\data_out_frame[25] [6]), .I1(\data_out_frame[23] [5]), 
            .I2(n43254), .I3(n44012), .O(n44659));
    defparam i2_3_lut_4_lut_adj_1492.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1493 (.I0(n27357), .I1(n43496), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4711));
    defparam i1_2_lut_adj_1493.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_1494 (.I0(\data_out_frame[16] [4]), .I1(n26950), 
            .I2(n10_adj_4455), .I3(n41232), .O(n40271));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1494.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46321), .I3(n46319), .O(n7_adj_4600));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46282), .I3(n46280), .O(n7_adj_4576));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i15_4_lut_adj_1495 (.I0(n29_adj_4708), .I1(n26580), .I2(n26_adj_4707), 
            .I3(n26599), .O(n32_adj_4712));
    defparam i15_4_lut_adj_1495.LUT_INIT = 16'h0020;
    SB_LUT4 i4_4_lut_adj_1496 (.I0(\data_out_frame[17] [7]), .I1(n42978), 
            .I2(n43417), .I3(n6_adj_4711), .O(n44251));
    defparam i4_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1497 (.I0(n2_adj_4470), .I1(n21657), .I2(n42830), 
            .I3(\FRAME_MATCHER.state_c [28]), .O(n42204));
    defparam i1_2_lut_4_lut_adj_1497.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_1498 (.I0(n2_adj_4470), .I1(n21657), .I2(n42830), 
            .I3(\FRAME_MATCHER.state_c [29]), .O(n42190));
    defparam i1_2_lut_4_lut_adj_1498.LUT_INIT = 16'hea00;
    SB_LUT4 i1_2_lut_4_lut_adj_1499 (.I0(n2_adj_4470), .I1(n21657), .I2(n42830), 
            .I3(\FRAME_MATCHER.state_c [31]), .O(n42168));
    defparam i1_2_lut_4_lut_adj_1499.LUT_INIT = 16'hea00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46309), .I3(n46307), .O(n7_adj_4577));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1500 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [4]), 
            .I3(GND_net), .O(n42270));
    defparam i1_2_lut_3_lut_adj_1500.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1501 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [5]), 
            .I3(GND_net), .O(n42272));
    defparam i1_2_lut_3_lut_adj_1501.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n46315), .I3(n46313), .O(n7_adj_4592));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i31126_2_lut (.I0(n27062), .I1(n27500), .I2(GND_net), .I3(GND_net), 
            .O(n46149));
    defparam i31126_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1502 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [6]), 
            .I3(GND_net), .O(n42274));
    defparam i1_2_lut_3_lut_adj_1502.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1503 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [7]), 
            .I3(GND_net), .O(n42276));
    defparam i1_2_lut_3_lut_adj_1503.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1504 (.I0(n44251), .I1(n43180), .I2(n44262), 
            .I3(\data_out_frame[11] [3]), .O(n12_adj_4713));
    defparam i5_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1505 (.I0(n46149), .I1(n32_adj_4712), .I2(n28_adj_4710), 
            .I3(n46147), .O(\FRAME_MATCHER.state_31__N_2724 [3]));
    defparam i16_4_lut_adj_1505.LUT_INIT = 16'h0040;
    SB_LUT4 i1_2_lut_3_lut_adj_1506 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [9]), 
            .I3(GND_net), .O(n42282));
    defparam i1_2_lut_3_lut_adj_1506.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1507 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [10]), 
            .I3(GND_net), .O(n7_adj_4669));
    defparam i1_2_lut_3_lut_adj_1507.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1508 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [11]), 
            .I3(GND_net), .O(n42284));
    defparam i1_2_lut_3_lut_adj_1508.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1509 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [12]), 
            .I3(GND_net), .O(n42286));
    defparam i1_2_lut_3_lut_adj_1509.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_4_lut_adj_1510 (.I0(\FRAME_MATCHER.state_31__N_2724 [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n34626), .I3(n27804), .O(n23568));
    defparam i2_4_lut_adj_1510.LUT_INIT = 16'h8808;
    SB_LUT4 i1_3_lut_4_lut_adj_1511 (.I0(n3813), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n29908), .I3(n771), .O(n42830));
    defparam i1_3_lut_4_lut_adj_1511.LUT_INIT = 16'haaba;
    SB_LUT4 i1_2_lut_3_lut_adj_1512 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [17]), 
            .I3(GND_net), .O(n7_adj_4668));
    defparam i1_2_lut_3_lut_adj_1512.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1513 (.I0(\state[0] ), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(GND_net), .O(n7233));
    defparam i1_2_lut_3_lut_adj_1513.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut_adj_1514 (.I0(\data_out_frame[13] [5]), .I1(n12_adj_4713), 
            .I2(n43398), .I3(\data_out_frame[13] [6]), .O(n41090));
    defparam i6_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(\FRAME_MATCHER.state_c [16]), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4714));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1516 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [18]), 
            .I3(GND_net), .O(n42304));
    defparam i1_2_lut_3_lut_adj_1516.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1517 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [19]), 
            .I3(GND_net), .O(n7_adj_4667));
    defparam i1_2_lut_3_lut_adj_1517.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1518 (.I0(\FRAME_MATCHER.state_c [27]), .I1(\FRAME_MATCHER.state_c [23]), 
            .I2(\FRAME_MATCHER.state_c [15]), .I3(\FRAME_MATCHER.state_c [26]), 
            .O(n12_adj_4715));   // verilog/coms.v(151[5:27])
    defparam i5_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1519 (.I0(\FRAME_MATCHER.state_c [17]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(\FRAME_MATCHER.state_c [18]), .I3(\FRAME_MATCHER.state_c [24]), 
            .O(n48));
    defparam i3_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1520 (.I0(n42891), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[22] [7]), .I3(n43148), .O(n10_adj_4631));
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1521 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [20]), 
            .I3(GND_net), .O(n42244));
    defparam i1_2_lut_3_lut_adj_1521.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_4_lut_adj_1522 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n48), 
            .I2(n12_adj_4715), .I3(n8_adj_4714), .O(n4_adj_4544));   // verilog/coms.v(151[5:27])
    defparam i1_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1523 (.I0(n41208), .I1(n41090), .I2(\data_out_frame[25] [1]), 
            .I3(GND_net), .O(n43199));
    defparam i2_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1524 (.I0(\data_out_frame[21][0] ), .I1(\data_out_frame[23] [3]), 
            .I2(\data_out_frame[25] [4]), .I3(GND_net), .O(n6_adj_4449));
    defparam i1_2_lut_3_lut_adj_1524.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1525 (.I0(\data_out_frame[22] [5]), .I1(n43353), 
            .I2(n41115), .I3(\data_out_frame[18] [3]), .O(n41236));
    defparam i1_2_lut_4_lut_adj_1525.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33763 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48780));
    defparam byte_transmit_counter_0__bdd_4_lut_33763.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_3_lut_adj_1526 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n41175), .I3(GND_net), .O(n10_adj_4446));
    defparam i2_2_lut_3_lut_adj_1526.LUT_INIT = 16'h6969;
    SB_LUT4 i24588_2_lut_3_lut (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [21]), 
            .I3(GND_net), .O(n39601));
    defparam i24588_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1527 (.I0(\data_out_frame[22] [4]), .I1(n43197), 
            .I2(\data_out_frame[24] [5]), .I3(\data_out_frame[24] [4]), 
            .O(n6_adj_4444));
    defparam i1_2_lut_4_lut_adj_1527.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1528 (.I0(\data_out_frame[24] [4]), .I1(\data_out_frame[24] [3]), 
            .I2(n41175), .I3(GND_net), .O(n6_adj_4443));
    defparam i1_2_lut_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1529 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [22]), 
            .I3(GND_net), .O(n7_adj_4665));
    defparam i1_2_lut_3_lut_adj_1529.LUT_INIT = 16'he0e0;
    SB_LUT4 n48780_bdd_4_lut (.I0(n48780), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48783));
    defparam n48780_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1530 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [23]), 
            .I3(GND_net), .O(n42306));
    defparam i1_2_lut_3_lut_adj_1530.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1531 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [24]), 
            .I3(GND_net), .O(n42248));
    defparam i1_2_lut_3_lut_adj_1531.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1532 (.I0(\data_out_frame[25] [6]), .I1(n41177), 
            .I2(n41135), .I3(\data_out_frame[23] [4]), .O(n6));
    defparam i1_2_lut_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1533 (.I0(\FRAME_MATCHER.state_c [25]), .I1(\FRAME_MATCHER.state_c [28]), 
            .I2(\FRAME_MATCHER.state_c [9]), .I3(\FRAME_MATCHER.state_c [12]), 
            .O(n12_adj_4534));   // verilog/coms.v(127[12] 300[6])
    defparam i5_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i33671_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n34624), .I3(GND_net), .O(n34718));
    defparam i33671_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_adj_1534 (.I0(\data_out_frame[16] [2]), .I1(n41182), 
            .I2(GND_net), .I3(GND_net), .O(n43006));
    defparam i1_2_lut_adj_1534.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1535 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n75));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_3_lut_adj_1535.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_adj_1536 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(GND_net), .O(n42308));
    defparam i1_2_lut_3_lut_adj_1536.LUT_INIT = 16'he0e0;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[24] [3]), .I1(n43006), .I2(n43199), 
            .I3(\data_out_frame[24] [1]), .O(n56));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4504));
    defparam select_658_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4502));
    defparam select_658_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19_4_lut_adj_1537 (.I0(n40261), .I1(n43290), .I2(n43090), 
            .I3(n42858), .O(n55));
    defparam i19_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(n44262), .I1(\data_out_frame[23] [1]), .I2(\data_out_frame[17] [1]), 
            .I3(\data_out_frame[24] [0]), .O(n63_adj_4716));
    defparam i27_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1538 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [26]), 
            .I3(GND_net), .O(n42310));
    defparam i1_2_lut_3_lut_adj_1538.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1539 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(GND_net), .O(n33802));
    defparam i1_2_lut_3_lut_adj_1539.LUT_INIT = 16'he0e0;
    SB_LUT4 i21119_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n34624), .I2(GND_net), 
            .I3(GND_net), .O(n34628));
    defparam i21119_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28581_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43600));
    defparam i28581_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i31166_4_lut (.I0(n42854), .I1(n4_adj_4544), .I2(\FRAME_MATCHER.state_c [4]), 
            .I3(n4_adj_4535), .O(n34377));
    defparam i31166_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [28]), 
            .I3(GND_net), .O(n42312));
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1541 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n19789));   // verilog/coms.v(214[11:56])
    defparam i2_3_lut_adj_1541.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1542 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [29]), 
            .I3(GND_net), .O(n7_adj_4664));
    defparam i1_2_lut_3_lut_adj_1542.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1543 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [30]), 
            .I3(GND_net), .O(n7_adj_4663));
    defparam i1_2_lut_3_lut_adj_1543.LUT_INIT = 16'he0e0;
    SB_LUT4 i20930_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n34434));
    defparam i20930_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1544 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n34434), .I3(byte_transmit_counter[2]), .O(n34544));
    defparam i2_4_lut_adj_1544.LUT_INIT = 16'h8880;
    SB_LUT4 i28748_4_lut (.I0(n34377), .I1(\FRAME_MATCHER.state [1]), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n43600), .O(n43770));
    defparam i28748_4_lut.LUT_INIT = 16'hfaea;
    SB_LUT4 i3_4_lut_adj_1545 (.I0(n34544), .I1(n44678), .I2(n33792), 
            .I3(n19789), .O(n44527));
    defparam i3_4_lut_adj_1545.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1546 (.I0(n1), .I1(n2_adj_4682), .I2(\FRAME_MATCHER.state_c [31]), 
            .I3(GND_net), .O(n42268));
    defparam i1_2_lut_3_lut_adj_1546.LUT_INIT = 16'he0e0;
    SB_LUT4 i24_4_lut_adj_1547 (.I0(n43278), .I1(n43196), .I2(n43216), 
            .I3(n43168), .O(n60));
    defparam i24_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n43074), .I1(\data_out_frame[21][2] ), .I2(n42871), 
            .I3(\data_out_frame[24] [2]), .O(n58));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4500));
    defparam select_658_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4498));
    defparam select_658_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4496));
    defparam select_658_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4494));
    defparam select_658_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23_4_lut (.I0(n44005), .I1(n43514), .I2(\data_out_frame[23] [7]), 
            .I3(n43365), .O(n59));
    defparam i23_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut (.I0(\data_out_frame[22] [0]), .I1(n43248), .I2(n43484), 
            .I3(n43187), .O(n57));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4492));
    defparam select_658_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4490));
    defparam select_658_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26_4_lut (.I0(n44237), .I1(n40238), .I2(\data_out_frame[19] [6]), 
            .I3(\data_out_frame[16] [1]), .O(n62));
    defparam i26_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_658_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4488));
    defparam select_658_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4486));
    defparam select_658_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32_3_lut (.I0(n63_adj_4716), .I1(n55), .I2(n56), .I3(GND_net), 
            .O(n68));
    defparam i32_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut_adj_1548 (.I0(n43088), .I1(n42881), .I2(n43068), 
            .I3(n42861), .O(n61));
    defparam i25_4_lut_adj_1548.LUT_INIT = 16'h9669;
    SB_LUT4 select_658_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4484));
    defparam select_658_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    uart_tx tx (.\r_SM_Main_2__N_3613[1] (\r_SM_Main_2__N_3613[1] ), .GND_net(GND_net), 
            .r_SM_Main({r_SM_Main}), .CLK_c(CLK_c), .\r_SM_Main_2__N_3616[0] (r_SM_Main_2__N_3616[0]), 
            .n18940(n18940), .r_Bit_Index({Open_30, Open_31, \r_Bit_Index[0] }), 
            .tx_o(tx_o), .tx_data({tx_data}), .n27763(n27763), .n28054(n28054), 
            .VCC_net(VCC_net), .n48986(n48986), .n28365(n28365), .n28159(n28159), 
            .tx_active(tx_active), .n4(n4_adj_10), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.\r_Bit_Index[0] (\r_Bit_Index[0]_adj_11 ), .GND_net(GND_net), 
            .n27767(n27767), .r_SM_Main({r_SM_Main_adj_18}), .n28056(n28056), 
            .\r_SM_Main_2__N_3542[2] (\r_SM_Main_2__N_3542[2] ), .r_Rx_Data(r_Rx_Data), 
            .n26339(n26339), .n26334(n26334), .n33899(n33899), .CLK_c(CLK_c), 
            .RX_N_10(RX_N_10), .VCC_net(VCC_net), .n28368(n28368), .n42422(n42422), 
            .rx_data_ready(rx_data_ready), .n28142(n28142), .rx_data({rx_data}), 
            .n28141(n28141), .n28140(n28140), .n28139(n28139), .n28138(n28138), 
            .n28128(n28128), .n28127(n28127), .n42722(n42722), .n4(n4_adj_15), 
            .n4_adj_8(n4_adj_16), .n4_adj_9(n4_adj_17), .n28372(n28372)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (\r_SM_Main_2__N_3613[1] , GND_net, r_SM_Main, CLK_c, 
            \r_SM_Main_2__N_3616[0] , n18940, r_Bit_Index, tx_o, tx_data, 
            n27763, n28054, VCC_net, n48986, n28365, n28159, tx_active, 
            n4, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output \r_SM_Main_2__N_3613[1] ;
    input GND_net;
    output [2:0]r_SM_Main;
    input CLK_c;
    input \r_SM_Main_2__N_3616[0] ;
    output n18940;
    output [2:0]r_Bit_Index;
    output tx_o;
    input [7:0]tx_data;
    output n27763;
    output n28054;
    input VCC_net;
    input n48986;
    input n28365;
    input n28159;
    output tx_active;
    output n4;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n44788, n10, n27948, n1;
    wire [8:0]n41;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n46334, n46335, n46338, n46337, n3, n25891, n21053;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index_c;   // verilog/uart_tx.v(33[16:27])
    
    wire n39055, n39054, n39053, n39052, n39051, n39050, n39049, 
        n39048, n34387, n21052, o_Tx_Serial_N_3644, n3_adj_4434, n48792;
    
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n44788));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[8]), .I2(n44788), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3613[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i33015_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n27948));
    defparam i33015_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR r_Clock_Count_2201__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i5560_2_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18940));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5560_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31253_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n46334));
    defparam i31253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31254_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n46335));
    defparam i31254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31257_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n46338));
    defparam i31257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31256_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n46337));
    defparam i31256_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n25891), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n21053), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(CLK_c), .E(n27763), 
            .D(n307[1]), .R(n28054));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(CLK_c), .E(n27763), 
            .D(n307[2]), .R(n28054));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2201__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n27948));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Clock_Count_2201_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n39055), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2201_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n39054), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_9 (.CI(n39054), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n39055));
    SB_LUT4 r_Clock_Count_2201_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n39053), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_8 (.CI(n39053), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n39054));
    SB_LUT4 r_Clock_Count_2201_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n39052), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_7 (.CI(n39052), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n39053));
    SB_LUT4 r_Clock_Count_2201_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n39051), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_6 (.CI(n39051), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n39052));
    SB_LUT4 r_Clock_Count_2201_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n39050), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_5 (.CI(n39050), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n39051));
    SB_LUT4 r_Clock_Count_2201_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n39049), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_4 (.CI(n39049), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n39050));
    SB_LUT4 r_Clock_Count_2201_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n39048), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_3 (.CI(n39048), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n39049));
    SB_LUT4 r_Clock_Count_2201_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n39048));
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n48986));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2363_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2363_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i14543_3_lut (.I0(n27763), .I1(n34387), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28054));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14543_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2356_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2356_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n34387));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7664_4_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(n34387), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3613[1] ), .O(n21052));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7664_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7665_3_lut (.I0(n21052), .I1(\r_SM_Main_2__N_3613[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21053));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7665_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3644), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i9728_2_lut_3_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4434));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i9728_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n28365));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n28159));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4434), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n25891), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n25891), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n25891), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n25891), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n25891), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n25891), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n25891), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index_c[1]), .I1(n46337), 
            .I2(n46338), .I3(r_Bit_Index_c[2]), .O(n48792));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48792_bdd_4_lut (.I0(n48792), .I1(n46335), .I2(n46334), .I3(r_Bit_Index_c[2]), 
            .O(o_Tx_Serial_N_3644));
    defparam n48792_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3613[1] ), .O(n27763));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3616[0] ), 
            .I3(r_SM_Main[1]), .O(n25891));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (\r_Bit_Index[0] , GND_net, n27767, r_SM_Main, n28056, 
            \r_SM_Main_2__N_3542[2] , r_Rx_Data, n26339, n26334, n33899, 
            CLK_c, RX_N_10, VCC_net, n28368, n42422, rx_data_ready, 
            n28142, rx_data, n28141, n28140, n28139, n28138, n28128, 
            n28127, n42722, n4, n4_adj_8, n4_adj_9, n28372) /* synthesis syn_module_defined=1 */ ;
    output \r_Bit_Index[0] ;
    input GND_net;
    output n27767;
    output [2:0]r_SM_Main;
    output n28056;
    output \r_SM_Main_2__N_3542[2] ;
    output r_Rx_Data;
    output n26339;
    output n26334;
    output n33899;
    input CLK_c;
    input RX_N_10;
    input VCC_net;
    input n28368;
    input n42422;
    output rx_data_ready;
    input n28142;
    output [7:0]rx_data;
    input n28141;
    input n28140;
    input n28139;
    input n28138;
    input n28128;
    input n28127;
    input n42722;
    output n4;
    output n4_adj_8;
    output n4_adj_9;
    input n28372;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]n326;
    
    wire n34381;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n6, n46121, n6_adj_4430, n26230, n7, n43772, n27957;
    wire [2:0]r_SM_Main_2__N_3548;
    
    wire n6_adj_4431, n27698, n26259;
    wire [7:0]n37;
    
    wire n3, r_Rx_Data_R, n39047, n39046, n39045, n39044, n39043, 
        n39042, n39041, n47191, n34448, n34516, n1;
    
    SB_LUT4 i2341_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2341_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n34381));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i14545_3_lut (.I0(n27767), .I1(n34381), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28056));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14545_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2334_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2334_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i31098_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n46121));
    defparam i31098_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4430));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20886_4_lut (.I0(r_Clock_Count[0]), .I1(n26230), .I2(n6_adj_4430), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3542[2] ));
    defparam i20886_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n26230));   // verilog/uart_rx.v(68[17:52])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_880 (.I0(r_Rx_Data), .I1(n26230), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_880.LUT_INIT = 16'heeee;
    SB_LUT4 i28750_4_lut (.I0(n46121), .I1(r_SM_Main[0]), .I2(n7), .I3(n6), 
            .O(n43772));
    defparam i28750_4_lut.LUT_INIT = 16'hccc4;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n43772), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[1]), .O(n27957));
    defparam i1_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i2_2_lut_adj_881 (.I0(r_SM_Main_2__N_3548[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4431));
    defparam i2_2_lut_adj_881.LUT_INIT = 16'h4444;
    SB_LUT4 i33003_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4431), 
            .I3(r_Rx_Data), .O(n27698));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33003_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i1_2_lut_adj_882 (.I0(n26259), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26339));
    defparam i1_2_lut_adj_882.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_883 (.I0(n26259), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26334));
    defparam i1_2_lut_adj_883.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20408_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33899));
    defparam i20408_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR r_Clock_Count_2199__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n27698), 
            .D(n37[1]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n27698), 
            .D(n37[2]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n27698), 
            .D(n37[3]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n27698), 
            .D(n37[4]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n27698), 
            .D(n37[5]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n27698), 
            .D(n37[6]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n27698), 
            .D(n37[7]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n27767), 
            .D(n326[1]), .R(n28056));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n27767), 
            .D(n326[2]), .R(n28056));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 r_Clock_Count_2199_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n39047), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2199_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n39046), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_8 (.CI(n39046), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n39047));
    SB_LUT4 r_Clock_Count_2199_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n39045), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_7 (.CI(n39045), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n39046));
    SB_LUT4 r_Clock_Count_2199_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n39044), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_6 (.CI(n39044), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n39045));
    SB_LUT4 r_Clock_Count_2199_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n39043), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_5 (.CI(n39043), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n39044));
    SB_LUT4 r_Clock_Count_2199_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n39042), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_4 (.CI(n39042), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n39043));
    SB_LUT4 r_Clock_Count_2199_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n39041), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_3 (.CI(n39041), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n39042));
    SB_LUT4 r_Clock_Count_2199_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n39041));
    SB_LUT4 i32250_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n47191));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32250_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n47191), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n34448));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFFESR r_Clock_Count_2199__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n27698), 
            .D(n37[0]), .R(n27957));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n34381), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n34516));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n34516), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n26259));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n28368));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n42422));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n28142));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n28141));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n28140));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n28139));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n28138));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n28128));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n28127));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n27767));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n42722));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n34448), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_334_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_334_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_332_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_8));   // verilog/uart_rx.v(97[17:39])
    defparam equal_332_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_331_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_9));   // verilog/uart_rx.v(97[17:39])
    defparam equal_331_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n28372));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4_3_lut_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(n26230), .I3(n6), .O(r_SM_Main_2__N_3548[0]));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'hfff7;
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (reg_B, CLK_c, n45341, GND_net, data_i, 
            VCC_net, n28107, data_o, n28529, n28419);
    output [2:0]reg_B;
    input CLK_c;
    output n45341;
    input GND_net;
    input [2:0]data_i;
    input VCC_net;
    input n28107;
    output [2:0]data_o;
    input n28529;
    input n28419;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n16, n17, n6, cnt_next_9__N_812;
    wire [9:0]n45;
    
    wire n38985, n38984, n38983, n38982, n38981, n38980, n38979, 
        n38978, n38977;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[3]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[9]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[6]), .I2(n16), .I3(cnt_reg[5]), 
            .O(n45341));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(reg_B[1]), .I2(reg_A[0]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n45341), .I1(n6), .I2(reg_B[2]), .I3(reg_A[2]), 
            .O(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdffd;
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2191_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n38985), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2191_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n38984), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_10 (.CI(n38984), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n38985));
    SB_LUT4 cnt_reg_2191_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n38983), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_9 (.CI(n38983), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n38984));
    SB_LUT4 cnt_reg_2191_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n38982), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_8 (.CI(n38982), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n38983));
    SB_LUT4 cnt_reg_2191_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n38981), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_CARRY cnt_reg_2191_add_4_7 (.CI(n38981), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n38982));
    SB_LUT4 cnt_reg_2191_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n38980), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_6 (.CI(n38980), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n38981));
    SB_LUT4 cnt_reg_2191_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n38979), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_5 (.CI(n38979), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n38980));
    SB_LUT4 cnt_reg_2191_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n38978), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_4 (.CI(n38978), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n38979));
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2191_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n38977), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_3 (.CI(n38977), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n38978));
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2191_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n38977));
    SB_DFFSR cnt_reg_2191__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n28107));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n28529));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n28419));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (\state[0] , GND_net, read, \state[1] , \state[3] , 
            \state[0]_adj_6 , CLK_c, \state[2] , n5614, n28155, rw, 
            n42504, data_ready, n122, n10, \state_7__N_4103[3] , n7233, 
            \saved_addr[0] , sda_enable, VCC_net, \state_7__N_4087[0] , 
            scl_enable, scl, sda_out, n28135, data, n28134, n28133, 
            n28132, n28131, n28130, n28129, n4, n4_adj_7, n33869, 
            n28259, n28244, n26367, n26372) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[0] ;
    input GND_net;
    input read;
    output \state[1] ;
    output \state[3] ;
    output \state[0]_adj_6 ;
    input CLK_c;
    output \state[2] ;
    output [0:0]n5614;
    input n28155;
    output rw;
    input n42504;
    output data_ready;
    output n122;
    output n10;
    input \state_7__N_4103[3] ;
    input n7233;
    output \saved_addr[0] ;
    output sda_enable;
    input VCC_net;
    output \state_7__N_4087[0] ;
    output scl_enable;
    output scl;
    output sda_out;
    input n28135;
    output [7:0]data;
    input n28134;
    input n28133;
    input n28132;
    input n28131;
    input n28130;
    input n28129;
    output n4;
    output n4_adj_7;
    output n33869;
    input n28259;
    input n28244;
    output n26367;
    output n26372;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n27697, n27932, n10_c, n9, n144, n7, n26228, n39800;
    wire [15:0]delay_counter_15__N_3989;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire enable, n28, n26, n27, n25, n19, n42378;
    wire [15:0]n4272;
    
    wire n38302, n38301, n38300, n38299, n38298, n38297, n38296, 
        n38295, n38294, n38293, n38292, n38291, n38290, n38289, 
        n38288;
    
    SB_LUT4 i14434_2_lut (.I0(n27697), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27932));   // verilog/eeprom.v(26[8] 58[4])
    defparam i14434_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n27697));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i4_4_lut (.I0(\state[0] ), .I1(n10_c), .I2(\state[1] ), .I3(n9), 
            .O(n144));   // verilog/eeprom.v(51[5:9])
    defparam i4_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i3_4_lut (.I0(n7), .I1(\state[3] ), .I2(\state[0]_adj_6 ), 
            .I3(n26228), .O(n39800));   // verilog/eeprom.v(42[12:28])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[1]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[2]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[3]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[4]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[5]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[6]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[7]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[8]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[9]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[10]), .S(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[11]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[12]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n5614[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[13]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[14]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[15]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n26228));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n27697), 
            .D(delay_counter_15__N_3989[0]), .R(n27932));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n19));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n42378));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n28155));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n42504));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_962_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4272[15]), 
            .I3(n38302), .O(delay_counter_15__N_3989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_962_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4272[15]), 
            .I3(n38301), .O(delay_counter_15__N_3989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_16 (.CI(n38301), .I0(delay_counter[14]), .I1(n4272[15]), 
            .CO(n38302));
    SB_LUT4 add_962_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4272[15]), 
            .I3(n38300), .O(delay_counter_15__N_3989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_15 (.CI(n38300), .I0(delay_counter[13]), .I1(n4272[15]), 
            .CO(n38301));
    SB_LUT4 add_962_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4272[15]), 
            .I3(n38299), .O(delay_counter_15__N_3989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_14 (.CI(n38299), .I0(delay_counter[12]), .I1(n4272[15]), 
            .CO(n38300));
    SB_LUT4 add_962_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4272[15]), 
            .I3(n38298), .O(delay_counter_15__N_3989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_13 (.CI(n38298), .I0(delay_counter[11]), .I1(n4272[15]), 
            .CO(n38299));
    SB_LUT4 add_962_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4272[15]), 
            .I3(n38297), .O(delay_counter_15__N_3989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_12 (.CI(n38297), .I0(delay_counter[10]), .I1(n4272[15]), 
            .CO(n38298));
    SB_LUT4 add_962_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4272[15]), 
            .I3(n38296), .O(delay_counter_15__N_3989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_11 (.CI(n38296), .I0(delay_counter[9]), .I1(n4272[15]), 
            .CO(n38297));
    SB_LUT4 add_962_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4272[15]), 
            .I3(n38295), .O(delay_counter_15__N_3989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_10 (.CI(n38295), .I0(delay_counter[8]), .I1(n4272[15]), 
            .CO(n38296));
    SB_LUT4 add_962_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4272[15]), 
            .I3(n38294), .O(delay_counter_15__N_3989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_9 (.CI(n38294), .I0(delay_counter[7]), .I1(n4272[15]), 
            .CO(n38295));
    SB_LUT4 add_962_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4272[15]), 
            .I3(n38293), .O(delay_counter_15__N_3989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_8 (.CI(n38293), .I0(delay_counter[6]), .I1(n4272[15]), 
            .CO(n38294));
    SB_LUT4 add_962_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4272[15]), 
            .I3(n38292), .O(delay_counter_15__N_3989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_7 (.CI(n38292), .I0(delay_counter[5]), .I1(n4272[15]), 
            .CO(n38293));
    SB_LUT4 add_962_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4272[15]), 
            .I3(n38291), .O(delay_counter_15__N_3989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_6 (.CI(n38291), .I0(delay_counter[4]), .I1(n4272[15]), 
            .CO(n38292));
    SB_LUT4 add_962_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4272[15]), 
            .I3(n38290), .O(delay_counter_15__N_3989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_5 (.CI(n38290), .I0(delay_counter[3]), .I1(n4272[15]), 
            .CO(n38291));
    SB_LUT4 add_962_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4272[15]), 
            .I3(n38289), .O(delay_counter_15__N_3989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_4 (.CI(n38289), .I0(delay_counter[2]), .I1(n4272[15]), 
            .CO(n38290));
    SB_LUT4 add_962_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4272[15]), 
            .I3(n38288), .O(delay_counter_15__N_3989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_3 (.CI(n38288), .I0(delay_counter[1]), .I1(n4272[15]), 
            .CO(n38289));
    SB_LUT4 add_962_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4272[15]), 
            .I3(GND_net), .O(delay_counter_15__N_3989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4272[15]), 
            .CO(n38288));
    i2c_controller i2c (.n39800(n39800), .\state[0] (\state[0] ), .GND_net(GND_net), 
            .\state[1] (\state[1] ), .n144(n144), .n42378(n42378), .n122(n122), 
            .n19(n19), .CLK_c(CLK_c), .n10(n10), .\state[3] (\state[3] ), 
            .\state[2] (\state[2] ), .n10_adj_2(n10_c), .\state_7__N_4103[3] (\state_7__N_4103[3] ), 
            .n7233(n7233), .\saved_addr[0] (\saved_addr[0] ), .\state[1]_adj_3 (state[1]), 
            .\state[0]_adj_4 (\state[0]_adj_6 ), .sda_enable(sda_enable), 
            .VCC_net(VCC_net), .\state_7__N_4087[0] (\state_7__N_4087[0] ), 
            .enable(enable), .scl_enable(scl_enable), .n9(n9), .read(read), 
            .n26228(n26228), .n5614({n5614}), .scl(scl), .sda_out(sda_out), 
            .n28135(n28135), .data({data}), .n28134(n28134), .n28133(n28133), 
            .n28132(n28132), .n28131(n28131), .n28130(n28130), .n28129(n28129), 
            .n4(n4), .n4_adj_5(n4_adj_7), .n33869(n33869), .n28259(n28259), 
            .n28244(n28244), .n26367(n26367), .n26372(n26372), .n4256(n4272[15])) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n39800, \state[0] , GND_net, \state[1] , n144, 
            n42378, n122, n19, CLK_c, n10, \state[3] , \state[2] , 
            n10_adj_2, \state_7__N_4103[3] , n7233, \saved_addr[0] , 
            \state[1]_adj_3 , \state[0]_adj_4 , sda_enable, VCC_net, 
            \state_7__N_4087[0] , enable, scl_enable, n9, read, n26228, 
            n5614, scl, sda_out, n28135, data, n28134, n28133, 
            n28132, n28131, n28130, n28129, n4, n4_adj_5, n33869, 
            n28259, n28244, n26367, n26372, n4256) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input n39800;
    input \state[0] ;
    input GND_net;
    input \state[1] ;
    input n144;
    output n42378;
    output n122;
    output n19;
    input CLK_c;
    output n10;
    output \state[3] ;
    output \state[2] ;
    output n10_adj_2;
    input \state_7__N_4103[3] ;
    input n7233;
    output \saved_addr[0] ;
    output \state[1]_adj_3 ;
    output \state[0]_adj_4 ;
    output sda_enable;
    input VCC_net;
    output \state_7__N_4087[0] ;
    input enable;
    output scl_enable;
    output n9;
    input read;
    input n26228;
    output [0:0]n5614;
    output scl;
    output sda_out;
    input n28135;
    output [7:0]data;
    input n28134;
    input n28133;
    input n28132;
    input n28131;
    input n28130;
    input n28129;
    output n4;
    output n4_adj_5;
    output n33869;
    input n28259;
    input n28244;
    output n26367;
    output n26372;
    output n4256;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n43639, n42852, n44330, n43732;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n27946, n47244, n43675;
    wire [7:0]n119;
    
    wire n27743;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n28001;
    wire [5:0]n29;
    
    wire n12, n6685, n15, n43679, n37, n47190, n47178, n11, 
        n47284, n19209, n7136, n27930, n5, n6692, n34514, n44007, 
        n39091, n39090, n39089, n39088, n39087, enable_slow_N_4189, 
        n27655, n33878, n10_adj_4413, n44900, n34051, n34057, n43702, 
        n11_adj_4414, n44738, i2c_clk_N_4176, scl_enable_N_4177, n27927, 
        sda_out_adj_4415, n9_c, n11_adj_4416, n11_adj_4417, n33772, 
        n27537, n5_adj_4418, n11_adj_4419, n4_c, n33_adj_4420, n6502, 
        n34_adj_4421, n4_adj_4423, n7, n38441, n38440, n38439, n38438, 
        n38437, n38436, n38435, n148;
    
    SB_LUT4 i28619_2_lut (.I0(n39800), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n43639));
    defparam i28619_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n43639), .I1(\state[1] ), .I2(n42852), .I3(n144), 
            .O(n44330));   // verilog/eeprom.v(23[11:16])
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i1_4_lut (.I0(\state[0] ), .I1(n44330), .I2(n144), .I3(n43732), 
            .O(n42378));   // verilog/eeprom.v(23[11:16])
    defparam i1_4_lut.LUT_INIT = 16'hceee;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n27946));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i32363_4_lut (.I0(n122), .I1(n144), .I2(\state[1] ), .I3(n42852), 
            .O(n47244));   // verilog/eeprom.v(23[11:16])
    defparam i32363_4_lut.LUT_INIT = 16'hdc50;
    SB_LUT4 i45_4_lut (.I0(n47244), .I1(n144), .I2(\state[0] ), .I3(n43675), 
            .O(n19));   // verilog/eeprom.v(23[11:16])
    defparam i45_4_lut.LUT_INIT = 16'hc505;
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27743), .D(n119[1]), 
            .S(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27743), .D(n119[2]), 
            .S(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27743), .D(n119[3]), 
            .R(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27743), .D(n119[4]), 
            .R(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27743), .D(n119[5]), 
            .R(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27743), .D(n119[6]), 
            .R(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27743), .D(n119[7]), 
            .R(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2203_2204__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6685));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_2));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28658_2_lut (.I0(\state_7__N_4103[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n43679));
    defparam i28658_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n6685), .I1(n43679), .I2(n7233), .I3(n37), 
            .O(n27743));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i32207_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n47190));   // verilog/i2c_controller.v(198[28:35])
    defparam i32207_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i32197_4_lut (.I0(n47190), .I1(\state[1]_adj_3 ), .I2(counter[0]), 
            .I3(counter[2]), .O(n47178));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i32197_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i32442_4_lut (.I0(n47178), .I1(\state[2] ), .I2(\state[0]_adj_4 ), 
            .I3(n11), .O(n47284));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i32442_4_lut.LUT_INIT = 16'h0322;
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7136), 
            .D(n19209), .S(n27930));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1]_adj_3 ), .C(i2c_clk), .E(n6692), 
            .D(n5), .S(n34514));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i3_4_lut (.I0(n6692), .I1(\state[2] ), .I2(\state[1]_adj_3 ), 
            .I3(\state[3] ), .O(n44007));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 counter2_2203_2204_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n39091), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2203_2204_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n39090), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_6 (.CI(n39090), .I0(GND_net), .I1(counter2[4]), 
            .CO(n39091));
    SB_LUT4 counter2_2203_2204_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n39089), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_5 (.CI(n39089), .I0(GND_net), .I1(counter2[3]), 
            .CO(n39090));
    SB_LUT4 counter2_2203_2204_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n39088), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_4 (.CI(n39088), .I0(GND_net), .I1(counter2[2]), 
            .CO(n39089));
    SB_LUT4 counter2_2203_2204_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n39087), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_3 (.CI(n39087), .I0(GND_net), .I1(counter2[1]), 
            .CO(n39088));
    SB_LUT4 counter2_2203_2204_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n39087));
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4087[0] ), .C(CLK_c), .E(n27655), 
            .D(enable_slow_N_4189));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i2_4_lut_adj_866 (.I0(\state_7__N_4103[3] ), .I1(n33878), .I2(enable), 
            .I3(n10_adj_4413), .O(n44900));
    defparam i2_4_lut_adj_866.LUT_INIT = 16'h008c;
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6692), .D(n34051), 
            .S(n34057));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2_4_lut_adj_867 (.I0(n43702), .I1(\state_7__N_4103[3] ), .I2(n44900), 
            .I3(n11_adj_4414), .O(n44738));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i2_4_lut_adj_867.LUT_INIT = 16'hf5fd;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4176));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4177));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6692), .D(n44738), 
            .S(n44007));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_868 (.I0(i2c_clk), .I1(n27946), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4176));
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4415), .C(i2c_clk), .E(n27927), 
            .D(n47284));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27743), .D(n119[0]), 
            .S(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i33319_2_lut (.I0(\state_7__N_4103[3] ), .I1(n11_adj_4414), 
            .I2(GND_net), .I3(GND_net), .O(n34051));
    defparam i33319_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i20387_2_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(GND_net), .I3(GND_net), .O(n33878));
    defparam i20387_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_869 (.I0(\state[3] ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4413));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(GND_net), .I3(GND_net), .O(n9_c));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20282_2_lut (.I0(n11_adj_4416), .I1(n11_adj_4417), .I2(GND_net), 
            .I3(GND_net), .O(n33772));
    defparam i20282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33010_4_lut (.I0(n27537), .I1(n6685), .I2(n11_adj_4416), 
            .I3(n5_adj_4418), .O(n6692));
    defparam i33010_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i1_4_lut_adj_870 (.I0(n11_adj_4419), .I1(n11_adj_4414), .I2(\state_7__N_4103[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_870.LUT_INIT = 16'h5755;
    SB_LUT4 i1_2_lut_adj_871 (.I0(\state[2] ), .I1(\state[1]_adj_3 ), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(\state[1]_adj_3 ), .I1(n33_adj_4420), .I2(n37), 
            .I3(GND_net), .O(n27930));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i33033_4_lut (.I0(n6502), .I1(n34_adj_4421), .I2(n4_c), .I3(n37), 
            .O(n7136));
    defparam i33033_4_lut.LUT_INIT = 16'haf8c;
    SB_DFFSR counter2_2203_2204__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 equal_265_i9_2_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_265_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16746_4_lut (.I0(read), .I1(n122), .I2(\state[0] ), .I3(n26228), 
            .O(n5614[0]));   // verilog/eeprom.v(23[11:16])
    defparam i16746_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i15_4_lut (.I0(n33772), .I1(\state[0]_adj_4 ), .I2(n6692), 
            .I3(n4_adj_4423), .O(n7));   // verilog/i2c_controller.v(33[12:17])
    defparam i15_4_lut.LUT_INIT = 16'hfc5c;
    SB_LUT4 i20360_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i20360_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2604_2_lut (.I0(sda_out_adj_4415), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n38441), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n28135));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n28134));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n28133));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n28132));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n28131));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n28130));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n28129));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n38440), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter2_2203_2204__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n27946));   // verilog/i2c_controller.v(69[20:35])
    SB_CARRY sub_39_add_2_8 (.CI(n38440), .I0(counter[6]), .I1(VCC_net), 
            .CO(n38441));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n38439), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n38439), .I0(counter[5]), .I1(VCC_net), 
            .CO(n38440));
    SB_LUT4 equal_340_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_340_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_339_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_339_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20378_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33869));
    defparam i20378_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n38438), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n38438), .I0(counter[4]), .I1(VCC_net), 
            .CO(n38439));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n38437), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n38437), .I0(counter[3]), .I1(VCC_net), 
            .CO(n38438));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n38436), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28711_2_lut_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(n122), .I3(n39800), .O(n43732));
    defparam i28711_2_lut_4_lut_4_lut.LUT_INIT = 16'heac8;
    SB_CARRY sub_39_add_2_4 (.CI(n38436), .I0(counter[2]), .I1(VCC_net), 
            .CO(n38437));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n38435), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n38435), .I0(counter[1]), .I1(VCC_net), 
            .CO(n38436));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n38435));
    SB_LUT4 i33615_2_lut_3_lut_4_lut (.I0(\state_7__N_4087[0] ), .I1(\state[0]_adj_4 ), 
            .I2(\state[1]_adj_3 ), .I3(n10_adj_2), .O(enable_slow_N_4189));
    defparam i33615_2_lut_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0]_adj_4 ), 
            .I1(\state[1]_adj_3 ), .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_4419));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_264_i11_2_lut_3_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_264_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_141_i11_2_lut_3_lut_4_lut (.I0(\state[0]_adj_4 ), 
            .I1(\state[1]_adj_3 ), .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4417));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_141_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n122));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33031_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[2] ), 
            .I2(\state[1]_adj_3 ), .I3(\state[3] ), .O(n19209));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i33031_2_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(\state[1]_adj_3 ), .O(n27927));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0136;
    SB_LUT4 i1_2_lut_4_lut_adj_872 (.I0(\state[1]_adj_3 ), .I1(\state[3] ), 
            .I2(\state[2] ), .I3(\state[0]_adj_4 ), .O(n34_adj_4421));
    defparam i1_2_lut_4_lut_adj_872.LUT_INIT = 16'h1104;
    SB_LUT4 i3_2_lut_4_lut (.I0(\state[2] ), .I1(\state[0]_adj_4 ), .I2(\state[1]_adj_3 ), 
            .I3(\state[3] ), .O(n6502));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h0144;
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(GND_net), .O(n11));
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0]_adj_4 ), 
            .I3(\state[1]_adj_3 ), .O(n27537));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'ha888;
    SB_LUT4 i33329_3_lut_4_lut (.I0(n6692), .I1(n11_adj_4416), .I2(n11_adj_4417), 
            .I3(n15), .O(n34514));
    defparam i33329_3_lut_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_4416));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i153_2_lut_3_lut (.I0(\state[3] ), .I1(\state[0]_adj_4 ), .I2(\state[1]_adj_3 ), 
            .I3(GND_net), .O(n148));
    defparam i153_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 state_7__I_0_139_i11_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(n11_adj_4414));   // verilog/i2c_controller.v(117[5:13])
    defparam state_7__I_0_139_i11_2_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_DFFE state_i0_i0 (.Q(\state[0]_adj_4 ), .C(i2c_clk), .E(VCC_net), 
            .D(n7));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_4087[0] ), .I2(n122), 
            .I3(GND_net), .O(n27655));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n28259));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n28244));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2_4_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[3] ), .I3(\state[2] ), .O(scl_enable_N_4177));   // verilog/i2c_controller.v(33[12:17])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i28681_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[1]_adj_3 ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n43702));
    defparam i28681_2_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0]_adj_4 ), 
            .I3(GND_net), .O(n33_adj_4420));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h5252;
    SB_LUT4 i1_3_lut_4_lut_adj_873 (.I0(n9_c), .I1(n10_adj_4413), .I2(n148), 
            .I3(\state[2] ), .O(n5_adj_4418));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_3_lut_4_lut_adj_873.LUT_INIT = 16'h1f11;
    SB_LUT4 i33327_3_lut_4_lut (.I0(n9_c), .I1(n10_adj_4413), .I2(n11_adj_4417), 
            .I3(n6692), .O(n34057));   // verilog/i2c_controller.v(151[5:14])
    defparam i33327_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut_adj_874 (.I0(n9_c), .I1(n10_adj_4413), .I2(counter[0]), 
            .I3(GND_net), .O(n26367));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_874.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_875 (.I0(n9_c), .I1(n10_adj_4413), .I2(counter[0]), 
            .I3(GND_net), .O(n26372));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_875.LUT_INIT = 16'hfefe;
    SB_LUT4 i28621_2_lut_4_lut (.I0(\state[0]_adj_4 ), .I1(\state[3] ), 
            .I2(\state[2] ), .I3(n43679), .O(n28001));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i28621_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_4_lut_adj_876 (.I0(\state[3] ), .I1(\state[1]_adj_3 ), 
            .I2(\state[2] ), .I3(\state[0]_adj_4 ), .O(n37));
    defparam i1_4_lut_4_lut_adj_876.LUT_INIT = 16'h0554;
    SB_LUT4 i1_2_lut_4_lut_adj_877 (.I0(\state[0] ), .I1(\state[1] ), .I2(n122), 
            .I3(read), .O(n42852));
    defparam i1_2_lut_4_lut_adj_877.LUT_INIT = 16'hc8ff;
    SB_LUT4 i28654_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n122), 
            .I3(n39800), .O(n43675));
    defparam i28654_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i1_3_lut_4_lut_adj_878 (.I0(\state[2] ), .I1(n148), .I2(n5_adj_4418), 
            .I3(\state_7__N_4087[0] ), .O(n4_adj_4423));
    defparam i1_3_lut_4_lut_adj_878.LUT_INIT = 16'hf1f0;
    SB_LUT4 i1_2_lut_3_lut_adj_879 (.I0(\state[2] ), .I1(n148), .I2(n26228), 
            .I3(GND_net), .O(n4256));
    defparam i1_2_lut_3_lut_adj_879.LUT_INIT = 16'h1010;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (b_prev, GND_net, a_new, direction_N_3907, 
            ENCODER1_B_N_keep, n1668, ENCODER1_A_N_keep, encoder1_position, 
            VCC_net, n28417, n1673) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3907;
    input ENCODER1_B_N_keep;
    input n1668;
    input ENCODER1_A_N_keep;
    output [31:0]encoder1_position;
    input VCC_net;
    input n28417;
    output n1673;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3910, debounce_cnt, a_prev, direction_N_3906;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_N_3913;
    wire [31:0]n133;
    
    wire n39023, n39022, n39021, n39020, n39019, n39018, n39017, 
        n39016, n39015, n39014, n39013, n39012, n39011, n39010, 
        n39009, n39008, n39007, n39006, n39005, n39004, n39003, 
        n39002, n39001, n39000, n38999, n38998, n38997, n38996, 
        n38995, n38994, n38993, n28418, n28334;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33024_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i33024_4_lut.LUT_INIT = 16'h8421;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2193_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[31]), .I3(n39023), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2193_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[30]), .I3(n39022), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_32 (.CI(n39022), .I0(direction_N_3906), 
            .I1(encoder1_position[30]), .CO(n39023));
    SB_LUT4 position_2193_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[29]), .I3(n39021), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_31 (.CI(n39021), .I0(direction_N_3906), 
            .I1(encoder1_position[29]), .CO(n39022));
    SB_LUT4 position_2193_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[28]), .I3(n39020), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_30 (.CI(n39020), .I0(direction_N_3906), 
            .I1(encoder1_position[28]), .CO(n39021));
    SB_LUT4 position_2193_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[27]), .I3(n39019), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_29 (.CI(n39019), .I0(direction_N_3906), 
            .I1(encoder1_position[27]), .CO(n39020));
    SB_LUT4 position_2193_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[26]), .I3(n39018), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_28 (.CI(n39018), .I0(direction_N_3906), 
            .I1(encoder1_position[26]), .CO(n39019));
    SB_LUT4 position_2193_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[25]), .I3(n39017), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_27 (.CI(n39017), .I0(direction_N_3906), 
            .I1(encoder1_position[25]), .CO(n39018));
    SB_LUT4 position_2193_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[24]), .I3(n39016), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_26 (.CI(n39016), .I0(direction_N_3906), 
            .I1(encoder1_position[24]), .CO(n39017));
    SB_LUT4 position_2193_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[23]), .I3(n39015), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_25 (.CI(n39015), .I0(direction_N_3906), 
            .I1(encoder1_position[23]), .CO(n39016));
    SB_LUT4 position_2193_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[22]), .I3(n39014), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_24 (.CI(n39014), .I0(direction_N_3906), 
            .I1(encoder1_position[22]), .CO(n39015));
    SB_LUT4 position_2193_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[21]), .I3(n39013), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_23 (.CI(n39013), .I0(direction_N_3906), 
            .I1(encoder1_position[21]), .CO(n39014));
    SB_LUT4 position_2193_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[20]), .I3(n39012), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_22 (.CI(n39012), .I0(direction_N_3906), 
            .I1(encoder1_position[20]), .CO(n39013));
    SB_LUT4 position_2193_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[19]), .I3(n39011), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_21 (.CI(n39011), .I0(direction_N_3906), 
            .I1(encoder1_position[19]), .CO(n39012));
    SB_LUT4 position_2193_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[18]), .I3(n39010), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_20 (.CI(n39010), .I0(direction_N_3906), 
            .I1(encoder1_position[18]), .CO(n39011));
    SB_LUT4 position_2193_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[17]), .I3(n39009), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_19 (.CI(n39009), .I0(direction_N_3906), 
            .I1(encoder1_position[17]), .CO(n39010));
    SB_LUT4 position_2193_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[16]), .I3(n39008), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_18 (.CI(n39008), .I0(direction_N_3906), 
            .I1(encoder1_position[16]), .CO(n39009));
    SB_LUT4 position_2193_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[15]), .I3(n39007), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_17 (.CI(n39007), .I0(direction_N_3906), 
            .I1(encoder1_position[15]), .CO(n39008));
    SB_LUT4 position_2193_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[14]), .I3(n39006), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_16 (.CI(n39006), .I0(direction_N_3906), 
            .I1(encoder1_position[14]), .CO(n39007));
    SB_LUT4 position_2193_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[13]), .I3(n39005), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_15 (.CI(n39005), .I0(direction_N_3906), 
            .I1(encoder1_position[13]), .CO(n39006));
    SB_LUT4 position_2193_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[12]), .I3(n39004), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_14 (.CI(n39004), .I0(direction_N_3906), 
            .I1(encoder1_position[12]), .CO(n39005));
    SB_LUT4 position_2193_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[11]), .I3(n39003), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_13 (.CI(n39003), .I0(direction_N_3906), 
            .I1(encoder1_position[11]), .CO(n39004));
    SB_LUT4 position_2193_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[10]), .I3(n39002), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_12 (.CI(n39002), .I0(direction_N_3906), 
            .I1(encoder1_position[10]), .CO(n39003));
    SB_LUT4 position_2193_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[9]), .I3(n39001), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_11 (.CI(n39001), .I0(direction_N_3906), 
            .I1(encoder1_position[9]), .CO(n39002));
    SB_LUT4 position_2193_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[8]), .I3(n39000), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_10 (.CI(n39000), .I0(direction_N_3906), 
            .I1(encoder1_position[8]), .CO(n39001));
    SB_LUT4 position_2193_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[7]), .I3(n38999), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_9 (.CI(n38999), .I0(direction_N_3906), 
            .I1(encoder1_position[7]), .CO(n39000));
    SB_LUT4 position_2193_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[6]), .I3(n38998), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_8 (.CI(n38998), .I0(direction_N_3906), 
            .I1(encoder1_position[6]), .CO(n38999));
    SB_LUT4 position_2193_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[5]), .I3(n38997), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_7 (.CI(n38997), .I0(direction_N_3906), 
            .I1(encoder1_position[5]), .CO(n38998));
    SB_LUT4 position_2193_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[4]), .I3(n38996), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_6 (.CI(n38996), .I0(direction_N_3906), 
            .I1(encoder1_position[4]), .CO(n38997));
    SB_LUT4 position_2193_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[3]), .I3(n38995), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_5 (.CI(n38995), .I0(direction_N_3906), 
            .I1(encoder1_position[3]), .CO(n38996));
    SB_LUT4 position_2193_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[2]), .I3(n38994), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_4 (.CI(n38994), .I0(direction_N_3906), 
            .I1(encoder1_position[2]), .CO(n38995));
    SB_LUT4 position_2193_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[1]), .I3(n38993), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_3 (.CI(n38993), .I0(direction_N_3906), 
            .I1(encoder1_position[1]), .CO(n38994));
    SB_LUT4 position_2193_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n38993));
    SB_DFFE position_2193__i31 (.Q(encoder1_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i30 (.Q(encoder1_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i29 (.Q(encoder1_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i28 (.Q(encoder1_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i27 (.Q(encoder1_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i26 (.Q(encoder1_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i25 (.Q(encoder1_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i24 (.Q(encoder1_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i23 (.Q(encoder1_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i22 (.Q(encoder1_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i21 (.Q(encoder1_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i20 (.Q(encoder1_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i19 (.Q(encoder1_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i18 (.Q(encoder1_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i17 (.Q(encoder1_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i16 (.Q(encoder1_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i15 (.Q(encoder1_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i14 (.Q(encoder1_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i13 (.Q(encoder1_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i12 (.Q(encoder1_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i11 (.Q(encoder1_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i10 (.Q(encoder1_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i9 (.Q(encoder1_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i8 (.Q(encoder1_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i7 (.Q(encoder1_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i6 (.Q(encoder1_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i5 (.Q(encoder1_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i4 (.Q(encoder1_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i3 (.Q(encoder1_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i2 (.Q(encoder1_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i1 (.Q(encoder1_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i0 (.Q(encoder1_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n28418));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1673), .C(n1668), .D(n28417));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n28334));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i14907_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n28418));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14823_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n28334));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14823_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (CS_c, CS_CLK_c, GND_net, state_7__N_4293, \data[15] , 
            n44589, n9, CLK_c, n11, VCC_net, n5, n5_adj_1, n33894, 
            n28153, current, n28623, n28622, n28621, n28620, n28619, 
            n28618, n28617, n28616, n28615, n28614, n28613, n28612, 
            n28125, n28124, \data[12] , n28123, \data[11] , n28122, 
            \data[10] , n28121, \data[9] , n28120, \data[8] , n28119, 
            \data[7] , n28118, \data[6] , n28117, \data[5] , n28116, 
            \data[4] , n28115, \data[3] , n28114, \data[2] , n28113, 
            \data[1] , n26390, n26377, n26385, n26380, n28427, \data[0] ) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output CS_c;
    output CS_CLK_c;
    input GND_net;
    output state_7__N_4293;
    output \data[15] ;
    output n44589;
    output n9;
    input CLK_c;
    output n11;
    input VCC_net;
    output n5;
    output n5_adj_1;
    output n33894;
    input n28153;
    output [12:0]current;
    input n28623;
    input n28622;
    input n28621;
    input n28620;
    input n28619;
    input n28618;
    input n28617;
    input n28616;
    input n28615;
    input n28614;
    input n28613;
    input n28612;
    input n28125;
    input n28124;
    output \data[12] ;
    input n28123;
    output \data[11] ;
    input n28122;
    output \data[10] ;
    input n28121;
    output \data[9] ;
    input n28120;
    output \data[8] ;
    input n28119;
    output \data[7] ;
    input n28118;
    output \data[6] ;
    input n28117;
    output \data[5] ;
    input n28116;
    output \data[4] ;
    input n28115;
    output \data[3] ;
    input n28114;
    output \data[2] ;
    input n28113;
    output \data[1] ;
    output n26390;
    output n26377;
    output n26385;
    output n26380;
    input n28427;
    output \data[0] ;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire clk_out;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n47179, n23309, n47180, n23307, n47181, n23305, n15, 
        n33987, n1, n27700, n10077, n27791, n27914;
    wire [7:0]n37;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n27966, n6, clk_slow_N_4206;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n6_adj_4404, n44197, n44224, n44580, delay_counter_15__N_4288;
    wire [4:0]n25;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n39040, n39039, n39038, n39037;
    wire [13:0]n61;
    
    wire n39036, n39035, n39034, n39033, n39032, n39031, n39030, 
        n39029, n39028, n39027, n39026, n39025, n39024, n38992, 
        n38991, n38990, n38989, n38988, n38987, n38986, n47225, 
        n6_adj_4406, clk_slow_N_4207, n23320, n9_adj_4407, n28157;
    
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i9833_3_lut (.I0(state[0]), .I1(n47179), .I2(state[1]), .I3(GND_net), 
            .O(n23309));   // verilog/tli4970.v(53[24:39])
    defparam i9833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9831_3_lut (.I0(state[0]), .I1(n47180), .I2(state[1]), .I3(GND_net), 
            .O(n23307));   // verilog/tli4970.v(53[24:39])
    defparam i9831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9829_3_lut (.I0(state[0]), .I1(n47181), .I2(state[1]), .I3(GND_net), 
            .O(n23305));   // verilog/tli4970.v(53[24:39])
    defparam i9829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33309_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n33987));
    defparam i33309_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4796_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));   // verilog/tli4970.v(41[5] 65[12])
    defparam i4796_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_7__I_0_76_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4293));   // verilog/tli4970.v(51[7:17])
    defparam state_7__I_0_76_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14318_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27700));
    defparam i14318_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n27791), .D(n10077), 
            .R(n27914));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNESR bit_counter_2192__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27700), 
            .D(n37[4]), .R(n27966));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27700), 
            .D(n37[5]), .R(n27966));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27700), 
            .D(n37[6]), .R(n27966));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27700), 
            .D(n37[7]), .R(n27966));   // verilog/tli4970.v(53[24:39])
    SB_LUT4 i2_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), .I3(GND_net), 
            .O(n44589));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_257_i9_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/tli4970.v(54[12:26])
    defparam equal_257_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_DFF clk_slow_62 (.Q(clk_slow), .C(CLK_c), .D(clk_slow_N_4206));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6), .O(n15));   // verilog/tli4970.v(54[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(delay_counter[5]), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4404));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(delay_counter[0]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[2]), .O(n44197));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_861 (.I0(n44197), .I1(n6_adj_4404), .I2(delay_counter[7]), 
            .I3(delay_counter[4]), .O(n44224));
    defparam i3_4_lut_adj_861.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_862 (.I0(n44224), .I1(delay_counter[8]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n44580));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'h8000;
    SB_LUT4 i2303_4_lut (.I0(n44580), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(delay_counter_15__N_4288));
    defparam i2303_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 mux_2295_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n10077));
    defparam mux_2295_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 counter_2196_2197_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n39040), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2196_2197_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n39039), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_5 (.CI(n39039), .I0(GND_net), .I1(counter[3]), 
            .CO(n39040));
    SB_LUT4 counter_2196_2197_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n39038), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_4 (.CI(n39038), .I0(GND_net), .I1(counter[2]), 
            .CO(n39039));
    SB_LUT4 counter_2196_2197_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n39037), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_3 (.CI(n39037), .I0(GND_net), .I1(counter[1]), 
            .CO(n39038));
    SB_LUT4 counter_2196_2197_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n39037));
    SB_LUT4 delay_counter_2194_2195_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n39036), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2194_2195_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n39035), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_14 (.CI(n39035), .I0(GND_net), 
            .I1(delay_counter[12]), .CO(n39036));
    SB_LUT4 delay_counter_2194_2195_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n39034), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_13 (.CI(n39034), .I0(GND_net), 
            .I1(delay_counter[11]), .CO(n39035));
    SB_LUT4 delay_counter_2194_2195_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n39033), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_12 (.CI(n39033), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n39034));
    SB_LUT4 delay_counter_2194_2195_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n39032), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_11 (.CI(n39032), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n39033));
    SB_LUT4 delay_counter_2194_2195_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n39031), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_10 (.CI(n39031), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n39032));
    SB_LUT4 delay_counter_2194_2195_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n39030), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_9 (.CI(n39030), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n39031));
    SB_LUT4 delay_counter_2194_2195_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n39029), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_8 (.CI(n39029), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n39030));
    SB_LUT4 delay_counter_2194_2195_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n39028), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_7 (.CI(n39028), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n39029));
    SB_LUT4 delay_counter_2194_2195_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n39027), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_6 (.CI(n39027), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n39028));
    SB_LUT4 delay_counter_2194_2195_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n39026), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_5 (.CI(n39026), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n39027));
    SB_LUT4 delay_counter_2194_2195_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n39025), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_4 (.CI(n39025), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n39026));
    SB_LUT4 delay_counter_2194_2195_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n39024), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_3 (.CI(n39024), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n39025));
    SB_LUT4 delay_counter_2194_2195_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n39024));
    SB_LUT4 bit_counter_2192_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n38992), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2192_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n38991), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_8 (.CI(n38991), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n38992));
    SB_LUT4 bit_counter_2192_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n38990), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_7 (.CI(n38990), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n38991));
    SB_LUT4 equal_314_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(52[9:26])
    defparam equal_314_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_313_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_1));   // verilog/tli4970.v(52[9:26])
    defparam equal_313_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 bit_counter_2192_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n38989), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_6 (.CI(n38989), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n38990));
    SB_LUT4 bit_counter_2192_add_4_5_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n38988), .O(n47181)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_5 (.CI(n38988), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n38989));
    SB_LUT4 bit_counter_2192_add_4_4_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n38987), .O(n47180)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_4 (.CI(n38987), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n38988));
    SB_LUT4 bit_counter_2192_add_4_3_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n38986), .O(n47179)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_3 (.CI(n38986), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n38987));
    SB_LUT4 bit_counter_2192_add_4_2_lut (.I0(n1), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n47225)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n38986));
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n27791), .D(n33987), 
            .S(n27914));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i2_2_lut_adj_863 (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4406));
    defparam i2_2_lut_adj_863.LUT_INIT = 16'heeee;
    SB_DFFSR counter_2196_2197__i5 (.Q(counter[4]), .C(CLK_c), .D(n25[4]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i2298_4_lut (.I0(counter[0]), .I1(counter[4]), .I2(n6_adj_4406), 
            .I3(counter[3]), .O(clk_slow_N_4207));
    defparam i2298_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 clk_slow_I_0_71_2_lut (.I0(clk_slow), .I1(clk_slow_N_4207), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4206));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_71_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR counter_2196_2197__i4 (.Q(counter[3]), .C(CLK_c), .D(n25[3]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2196_2197__i3 (.Q(counter[2]), .C(CLK_c), .D(n25[2]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2196_2197__i2 (.Q(counter[1]), .C(CLK_c), .D(n25[1]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2194_2195__i14 (.Q(delay_counter[13]), .C(clk_slow), 
            .D(n61[13]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i13 (.Q(delay_counter[12]), .C(clk_slow), 
            .D(n61[12]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n61[11]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n61[10]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n61[9]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n61[8]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n61[7]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n61[6]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n61[5]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n61[4]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n61[3]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n61[2]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n61[1]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNE bit_counter_2192__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27700), 
            .D(n23305));   // verilog/tli4970.v(53[24:39])
    SB_DFFNE bit_counter_2192__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27700), 
            .D(n23307));   // verilog/tli4970.v(53[24:39])
    SB_DFFNE bit_counter_2192__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27700), 
            .D(n23309));   // verilog/tli4970.v(53[24:39])
    SB_LUT4 i20403_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n33894));
    defparam i20403_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9841_3_lut (.I0(state[0]), .I1(n47225), .I2(state[1]), .I3(GND_net), 
            .O(n23320));   // verilog/tli4970.v(53[24:39])
    defparam i9841_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFN clk_out_66 (.Q(clk_out), .C(clk_slow), .D(n9_adj_4407));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN slave_select_65 (.Q(CS_c), .C(clk_slow), .D(n28157));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i0 (.Q(current[0]), .C(clk_slow), .D(n28153));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i1 (.Q(current[1]), .C(clk_slow), .D(n28623));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i2 (.Q(current[2]), .C(clk_slow), .D(n28622));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i3 (.Q(current[3]), .C(clk_slow), .D(n28621));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i4 (.Q(current[4]), .C(clk_slow), .D(n28620));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i5 (.Q(current[5]), .C(clk_slow), .D(n28619));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i6 (.Q(current[6]), .C(clk_slow), .D(n28618));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i7 (.Q(current[7]), .C(clk_slow), .D(n28617));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNE bit_counter_2192__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27700), 
            .D(n23320));   // verilog/tli4970.v(53[24:39])
    SB_DFFN current_i0_i8 (.Q(current[8]), .C(clk_slow), .D(n28616));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i9 (.Q(current[9]), .C(clk_slow), .D(n28615));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNSR delay_counter_2194_2195__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n61[0]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFN current_i0_i10 (.Q(current[10]), .C(clk_slow), .D(n28614));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFSR counter_2196_2197__i1 (.Q(counter[0]), .C(CLK_c), .D(n25[0]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFN current_i0_i11 (.Q(current[11]), .C(clk_slow), .D(n28613));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i12 (.Q(current[12]), .C(clk_slow), .D(n28612));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n28125));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n28124));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n28123));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n28122));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n28121));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n28120));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n28119));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n28118));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n28117));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n28116));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n28115));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n28114));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n28113));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n26390));   // verilog/tli4970.v(54[12:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_257_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[12:26])
    defparam equal_257_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_864 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n26377));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut_adj_864.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_865 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n26385));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut_adj_865.LUT_INIT = 16'hffbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n26380));   // verilog/tli4970.v(41[5] 65[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n28427));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i14646_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n28157));   // verilog/tli4970.v(41[5] 65[12])
    defparam i14646_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i33686_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9_adj_4407));   // verilog/tli4970.v(41[5] 65[12])
    defparam i33686_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i14456_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27966));   // verilog/tli4970.v(53[24:39])
    defparam i14456_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), .I3(delay_counter_15__N_4288), 
            .O(n27791));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i14403_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(delay_counter_15__N_4288), .O(n27914));
    defparam i14403_2_lut_4_lut.LUT_INIT = 16'h0b00;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, pwm_setpoint, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input [23:0]pwm_setpoint;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire pwm_out_N_797;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n45150, n22, n15, n20, n24, n19, pwm_counter_23__N_795;
    wire [23:0]n101;
    
    wire n38976, n38975, n38974, n38973, n38972, n38971, n38970, 
        n38969, n38968, n38967, n38966, n38965, n38964, n38963, 
        n41, n39, n45, n43, n38962, n38961, n38960, n38959, 
        n38958, n38957, n38956, n38955, n38954, n23, n25, n35, 
        n37, n29, n33, n11, n13, n15_adj_4401, n27, n9, n17, 
        n19_adj_4402, n21, n47267, n47261, n12, n30, n47317, n47562, 
        n47547, n47945, n31, n47771, n47999, n6, n47951, n47952, 
        n16, n24_adj_4403, n47519, n8, n47517, n47799, n47894, 
        n4, n47947, n47948, n47256, n10, n47528, n48001, n28, 
        n48043, n48044, n48022, n47521, n47955, n47589, n48009;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_797));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n45150));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[15]), .I1(pwm_counter[16]), .I2(pwm_counter[20]), 
            .I3(pwm_counter[19]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n45150), .I1(pwm_counter[22]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[13]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(pwm_counter[12]), .I3(pwm_counter[18]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[14]), .I1(pwm_counter[17]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33693_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(pwm_counter_23__N_795));   // verilog/pwm.v(18[8:40])
    defparam i33693_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 pwm_counter_2190_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n38976), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2190_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n38975), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_24 (.CI(n38975), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n38976));
    SB_LUT4 pwm_counter_2190_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n38974), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_23 (.CI(n38974), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n38975));
    SB_LUT4 pwm_counter_2190_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n38973), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_22 (.CI(n38973), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n38974));
    SB_LUT4 pwm_counter_2190_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n38972), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_21 (.CI(n38972), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n38973));
    SB_LUT4 pwm_counter_2190_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n38971), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_20 (.CI(n38971), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n38972));
    SB_LUT4 pwm_counter_2190_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n38970), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_19 (.CI(n38970), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n38971));
    SB_LUT4 pwm_counter_2190_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n38969), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_18 (.CI(n38969), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n38970));
    SB_LUT4 pwm_counter_2190_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n38968), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_17 (.CI(n38968), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n38969));
    SB_LUT4 pwm_counter_2190_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n38967), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_16 (.CI(n38967), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n38968));
    SB_LUT4 pwm_counter_2190_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n38966), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_15 (.CI(n38966), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n38967));
    SB_LUT4 pwm_counter_2190_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n38965), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_14 (.CI(n38965), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n38966));
    SB_DFFSR pwm_counter_2190__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2190_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n38964), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_counter_2190__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_CARRY pwm_counter_2190_add_4_13 (.CI(n38964), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n38965));
    SB_LUT4 pwm_counter_2190_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n38963), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY pwm_counter_2190_add_4_12 (.CI(n38963), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n38964));
    SB_LUT4 pwm_counter_2190_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n38962), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_11 (.CI(n38962), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n38963));
    SB_LUT4 pwm_counter_2190_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n38961), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_10 (.CI(n38961), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n38962));
    SB_LUT4 pwm_counter_2190_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n38960), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_9 (.CI(n38960), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n38961));
    SB_LUT4 pwm_counter_2190_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n38959), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_8 (.CI(n38959), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n38960));
    SB_LUT4 pwm_counter_2190_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n38958), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_7 (.CI(n38958), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n38959));
    SB_LUT4 pwm_counter_2190_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n38957), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_6 (.CI(n38957), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n38958));
    SB_LUT4 pwm_counter_2190_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n38956), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_5 (.CI(n38956), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n38957));
    SB_LUT4 pwm_counter_2190_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n38955), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_4 (.CI(n38955), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n38956));
    SB_LUT4 pwm_counter_2190_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n38954), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_3 (.CI(n38954), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n38955));
    SB_LUT4 pwm_counter_2190_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n38954));
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4401));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4402));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32186_4_lut (.I0(n21), .I1(n19_adj_4402), .I2(n17), .I3(n9), 
            .O(n47267));
    defparam i32186_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32180_4_lut (.I0(n27), .I1(n15_adj_4401), .I2(n13), .I3(n11), 
            .O(n47261));
    defparam i32180_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32481_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n47317), 
            .O(n47562));
    defparam i32481_4_lut.LUT_INIT = 16'heeef;
    SB_DFFSR pwm_counter_2190__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i32466_4_lut (.I0(n19_adj_4402), .I1(n17), .I2(n15_adj_4401), 
            .I3(n47562), .O(n47547));
    defparam i32466_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32864_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n47547), 
            .O(n47945));
    defparam i32864_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32690_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n47945), 
            .O(n47771));
    defparam i32690_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32918_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n47771), 
            .O(n47999));
    defparam i32918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32870_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n47951));   // verilog/pwm.v(21[8:24])
    defparam i32870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32871_3_lut (.I0(n47951), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n47952));   // verilog/pwm.v(21[8:24])
    defparam i32871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4403));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32438_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n47267), 
            .O(n47519));
    defparam i32438_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32718_4_lut (.I0(n24_adj_4403), .I1(n8), .I2(n45), .I3(n47517), 
            .O(n47799));   // verilog/pwm.v(21[8:24])
    defparam i32718_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32813_3_lut (.I0(n47952), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n47894));   // verilog/pwm.v(21[8:24])
    defparam i32813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i32866_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n47947));   // verilog/pwm.v(21[8:24])
    defparam i32866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32436_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n47517));
    defparam i32436_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32867_3_lut (.I0(n47947), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n47948));   // verilog/pwm.v(21[8:24])
    defparam i32867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32175_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n47261), 
            .O(n47256));
    defparam i32175_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32447_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n47528));
    defparam i32447_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32920_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n47528), 
            .O(n48001));   // verilog/pwm.v(21[8:24])
    defparam i32920_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32815_3_lut (.I0(n47948), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n28));   // verilog/pwm.v(21[8:24])
    defparam i32815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32962_4_lut (.I0(n28), .I1(n48001), .I2(n35), .I3(n47256), 
            .O(n48043));   // verilog/pwm.v(21[8:24])
    defparam i32962_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32963_3_lut (.I0(n48043), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n48044));   // verilog/pwm.v(21[8:24])
    defparam i32963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32941_3_lut (.I0(n48044), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n48022));   // verilog/pwm.v(21[8:24])
    defparam i32941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32440_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n47999), 
            .O(n47521));
    defparam i32440_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32874_4_lut (.I0(n47894), .I1(n47799), .I2(n45), .I3(n47519), 
            .O(n47955));   // verilog/pwm.v(21[8:24])
    defparam i32874_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32508_3_lut (.I0(n48022), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n47589));   // verilog/pwm.v(21[8:24])
    defparam i32508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32928_4_lut (.I0(n47589), .I1(n47955), .I2(n45), .I3(n47521), 
            .O(n48009));   // verilog/pwm.v(21[8:24])
    defparam i32928_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32929_3_lut (.I0(n48009), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_797));   // verilog/pwm.v(21[8:24])
    defparam i32929_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32236_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n47317));   // verilog/pwm.v(21[8:24])
    defparam i32236_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    
endmodule
