// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Dec  7 13:46:38 2021
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    
    wire n1759;
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(352[11:24])
    
    wire n60538;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(360[15:20])
    
    wire pwm_setpoint_23__N_207, n11648, n11650, n11652, n11654, n11656, 
        n11658, n11660, n11662, n11664, n11666, n11668, n11670, 
        n11672, n11674, n11676, n11678, n60537, n260, n11686, 
        n11684, n294, n298, n299, n300, n301, n302, n303, n304, 
        n305, n306, n307, n308, n309;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n22465, n60626;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216, n1761, n1763, n1765;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, n29619, RX_N_2, n1757, n1755, n1753, n1751, 
        n72122, n1749, n1747;
    wire [31:0]motor_state_23__N_91;
    wire [36:0]encoder1_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        read_N_409, n6, n34686, n1323, n62, n26, n1797;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1829, n1831, n39034;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    
    wire n72119, n60650, n25, n24, n23, n22, n21, n20, n19, 
        n60536, n29616, n29613, n19_adj_5708, n17, n16, n15, n13, 
        n11, n9, n18, n17_adj_5709, n2828, n16_adj_5710;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n15_adj_5711, n14, n13_adj_5712, n2, n14_adj_5713, n15_adj_5714, 
        n16_adj_5715, n17_adj_5716, n18_adj_5717, n19_adj_5718, n20_adj_5719, 
        n21_adj_5720, n22_adj_5721, n23_adj_5722, n24_adj_5723, n25_adj_5724, 
        n24_adj_5725, n39467, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n20682;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n4937, n4936, n4935, n4915, 
        n4914, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
        n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
        n4931, n4932, n4933, n4934, n60630, n3483, n2881, n15430, 
        n161, n39188, n34584, n48532, n56696, n1, n53594, n53746, 
        n53745, n53744, n53743, n53742, n53741, n53740, n53739, 
        n53738, n53737, n53736, n29097, n53577, n8, n59068, n24_adj_5726, 
        n63208, n17_adj_5727, n15_adj_5728, n8_adj_5729, n53735, n34395, 
        n34394, n53734, n53733, n53436, \FRAME_MATCHER.i_31__N_2509 , 
        n39530, n29520, n29513, n59922, n53732, n29501, n29498, 
        n29495, n29492, n29489, n29486, n29483, n29480, n29477, 
        n29473, n29466, n29463, n29460, n29459, n29456, n29451, 
        n29448, n29445, n29442, n29439, n29436, n60419, n29377, 
        n29347, n29346, n29345, n29344, n29343, n29342, n29341, 
        n29340, n29339, n29338, n29328, n29327, n29326, n29325, 
        n29324, n29323, n29322, n29321, n29320, n29319, n29318, 
        n29317, n29316, n29315, n29314, n29313, n29312, n29311, 
        n29310, n29239, n29238, n29237, n29236, n29235, n29214, 
        n29211, n29208, n29205, n29199, n29196, n29193, n29190, 
        n29187, n29184, n29181, n7, n6_adj_5730, n5, n4, n24_adj_5731, 
        n19_adj_5732, n17_adj_5733, n16_adj_5734, n15_adj_5735, n13_adj_5736, 
        n11_adj_5737, n9_adj_5738, n8_adj_5739, n7_adj_5740, n6_adj_5741, 
        n5_adj_5742, n4_adj_5743, n72092, n30, n70525, n23_adj_5744, 
        n21_adj_5745, n19_adj_5746, n17_adj_5747, n16_adj_5748, n15_adj_5749, 
        n13_adj_5750, n11_adj_5751, n10, n9_adj_5752, n8_adj_5753, 
        n7_adj_5754, n6_adj_5755, n4_adj_5756, n60632, n60631, n60535, 
        n60534, n60533, n60624, n28930, n60532, n60475, n60531, 
        n60530, n60529, n60544, n60528, n4_adj_5757, n4_adj_5758, 
        n4_adj_5759, n25158, n10_adj_5760, n6_adj_5761, n29178, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n53731, n63449, n53730, n25302, n11646, n60527, n238, 
        n258, n284, n290, n336, n337, n338, n339, n341, n342, 
        n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n53729, 
        n53728, n5227, n5224, n29175, n29172, n3172, n53727, n6_adj_5762, 
        n5_adj_5763, n15_adj_5764, n11_adj_5765, n60302;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, n39420, position_31__N_3836, 
        n45, n43, n41, n39, n33, n22661, n15_adj_5766;
    wire [1:0]a_new_adj_5908;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5909;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5769, b_prev_adj_5770, debounce_cnt_N_3833_adj_5771, 
        position_31__N_3836_adj_5772, n31, n72086, n65545, n12, n11_adj_5773, 
        n10_adj_5774, n4_adj_5775, n3, n2_adj_5776;
    wire [7:0]data_adj_5921;   // verilog/eeprom.v(23[12:16])
    wire [7:0]state_7__N_3918;
    
    wire n15440, n53726, n60627, n6910, n7_adj_5777, n71513, n53725, 
        n25345, n13228, clk_out;
    wire [15:0]data_adj_5928;   // verilog/tli4970.v(27[14:18])
    
    wire n22_adj_5786;
    wire [7:0]state_adj_5930;   // verilog/tli4970.v(29[13:18])
    
    wire n71401, n65211, n17_adj_5789, n35689, n15_adj_5790, n5_adj_5791, 
        n62322, n53724, n11680, n11682, state_7__N_4319, n9_adj_5792, 
        n8_adj_5793, n7_adj_5794, n6_adj_5795, n5_adj_5796, n29948, 
        n29945, n29942, n29939, n53593, n29936, n29933, n29930, 
        n25153, n60474, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n29927, n69921;
    wire [24:0]o_Rx_DV_N_3488;
    wire [2:0]r_SM_Main_2__N_3446;
    wire [2:0]r_SM_Main_adj_5944;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5945;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5946;   // verilog/uart_tx.v(34[16:27])
    
    wire n60951, n71483;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n39431, n29880, n29879, n29878, n29877, n29875, n29874, 
        n29872, n29871, n29869, n29868;
    wire [7:0]state_adj_5954;   // verilog/i2c_controller.v(33[12:17])
    
    wire enable_slow_N_4213, n8_adj_5810, n29866, n29865, n29864, 
        n29863, n29862, n29861, n29860, n29859, n29858;
    wire [7:0]state_7__N_4110;
    
    wire n29857, n29856, n29855, n29854, n29853, n29852, n29851, 
        n29850, n29849, n25348, n6714, n29848, n29847, n29846, 
        n29845, n29844, n29843, n29840, n29839;
    wire [7:0]state_7__N_4126;
    
    wire n29142, n29139, n29136, n60620, n60526, n60525, n60524, 
        n60640, n27664, n60477, n60523, n60639, n60522, n60521, 
        n60520, n60519, n60518, n27645, n60641, n60517, n60637, 
        n60545, n60516, n60515, n60619, n4_adj_5811, n8_adj_5812, 
        n10_adj_5813, n12_adj_5814, n20_adj_5815, n31_adj_5816, n37, 
        n60636, n60514, n39_adj_5817, n60513, n60512, n60511, n60510, 
        n60509, n60508, n60507, n60506, n60648, n60505, n60539, 
        n60649, n60541, n60504, n60503, n60647, n60502, n60501, 
        n60646, n60500, n13229, n15443, n71512, n13220, n15433, 
        n15434, n70762, n204, n13221, n10003, n71396, n54439, 
        n54438, n54437, n54436, n15425, n13222, n54435, n15435, 
        n54434, n54433, n131, n53692, n53691, n53690, n53689, 
        n53688, n53576, n72056, n71302, n53687, n53686, n53685, 
        n53592, n15426, n15436, n53964, n53963, n13223, n71942, 
        n53962, n53961, n53960, n53959, n53958, n53957, n53956, 
        n53575, n53684, n53955, n53954, n53683, n53682, n53591, 
        n53590, n53681, n53953, n53952, n53951, n53680, n53950, 
        n53679, n13224, n24820, n53949, n53948, n53947, n53946, 
        n53945, n53678, n53677, n53944, n15427, n53676, n53589, 
        n53675, n53574, n53674, n15437, n71247, n53673, n53672, 
        n15_adj_5818, n69867, n14_adj_5819, n13225, n71939, n60499, 
        n71218, n53671, n53588, n13226, n53587, n53670, n53934, 
        n15428, n15438, n60498, n53933, n53932, n25289, n53931, 
        n25_adj_5820, n60621, n53930, n60644, n60497, n39146, n13227, 
        n15429, n15439, n53929, n26311, n55945, n26215, n25298, 
        n71168, n60496, n60495, n60494, n60415, n60622, n60643, 
        n4_adj_5821, n6_adj_5822, n8_adj_5823, n9_adj_5824, n11_adj_5825, 
        n13_adj_5826, n15_adj_5827, n60642, n4_adj_5828, n6_adj_5829, 
        n8_adj_5830, n9_adj_5831, n27514, n27511, n27507, n60645, 
        n38, n39_adj_5832, n40, n41_adj_5833, n42, n43_adj_5834, 
        n44, n45_adj_5835, n29133, n29130, n15_adj_5836, n27489, 
        n60493, n27482, n15431, n60492, n27465, n60491, n60490, 
        n60543, n60489, n60638, n27441, n60488, n60635, n60487, 
        n60486, n60485, n60540, n60542, n60634, n60484, n14_adj_5837, 
        n56545, n56501, n56624, n60658, n60657, n60656, n60655, 
        n60654, n60653, n60652, n60651, n60483, n60618, n60482, 
        n60617, n60481, n60616, n60480, n60615, n60479, n60614, 
        n60613, n60478, n60612, n60611, n60610, n60609, n60608, 
        n60607, n60606, n60605, n29002, n60604, n60603, n60602, 
        n60601, n60600, n60599, n60598, n60597, n60596, n60595, 
        n60594, n60593, n60592, n60591, n60590, n60589, n60588, 
        n60587, n60586, n60585, n60584, n56640, n60583, n60582, 
        n60581, n60580, n60579, n60578, n60577, n60576, n60575, 
        n60574, n60573, n60572, n60571, n28828, n60570, n60569, 
        n60568, n60567, n60566, n60565, n60564, n60563, n60562, 
        n60561, n60560, n60559, n60558, n60557, n29020, n60556, 
        n60555, n60554, n53928, n60476, n60553, n60552, n60551, 
        n60550, n60549, n60548, n60547, n60546, n28127, n28117, 
        n28113, n28102, n60766, n28096, n60413, n60771, n28543, 
        n28534, n14_adj_5838, n13_adj_5839, n25156, n60633, n20628, 
        n15441, n9940, n9938, n27417, n72442, n71906, n71903, 
        n59876, n59930, n7_adj_5840, n53586, n11644, n65632, n29739, 
        n29738, n29736, n29734, n29733, n29732, n29731, n29730, 
        n29729, n29728, n29727, n29726, n29725, n29724, n29723, 
        n29722, n13211, n13210, n70965, n70964, n68899, n13212, 
        n29127, n29126, n29125, n29124, n29721, n29720, n29719, 
        n29718, n13213, n69733, n60700, n29123, n62711, n13214, 
        n20719, n29683, n13215, n29119, n53927, n29114, n29679, 
        n29674, n25712, n13217, n13216, n53926, n13218, n29671, 
        n29668, n29663, n29661, n29660, n29659, n29658, n29654, 
        n29652, n29646, n29645, n29644, n29642, n15442, n29110, 
        n29641, n29640, n29639, n29635, n71307, n29632, n29629, 
        n53925, n53924, n3_adj_5841, n31_adj_5842, n28, n1_adj_5843, 
        n70807, n53923, n53922, n53921, n53920, n60628, n21407, 
        n53919, n70435, n53918, n53917, n53916, n72053, n10_adj_5844, 
        n39001, n25994, n60625, n68794, n61210, n22_adj_5845, n60623, 
        n65193, n63296, n68790, n56754, n63448, n68775, n72606, 
        n6_adj_5846, n72329, n25732, n72323, n72317, n72311, n37935, 
        n37938, n25647, n37941, n72305, n60, n37953, n112, n37967, 
        n72299, n71550, n115, n72293, n72287, n37982, n94, n70806, 
        n72281, n65629, n55578, n72275, n72269, n110, n72263, 
        n72257, n13219, n25328, n34791, n25316, n25296, n38983, 
        n72251, n53585, n60629, n72245, n15432, n70524, n70523, 
        n56565, n72239, n69899, n69775, n39133, n39100, n53884, 
        n53573, n53883, n53882, n53881, n53880, n53584, n53879, 
        n53878, n6_adj_5847, n53877, n53876, n53875, n53874, n53873, 
        n4_adj_5848, n53872, n53871, n53870, n53869, n53868, n53867, 
        n53583, n53572, n72233, n53828, n53827, n53826, n53582, 
        n53825, n53824, n53823, n53822, n53821, n53820, n53581, 
        n53819, n53818, n53817, n53816, n53571, n69757, n53600, 
        n53599, n69754, n53580, n53579, n53598, n53597, n53578, 
        n53596, n72227, n53595, n53570, n70814, n72221, n70473, 
        n70960, n8_adj_5849, n69628, n69626, n70487, n72215, n69608, 
        n14_adj_5850, n69600, n10_adj_5851, n65191, n70493, n64235, 
        n62686, n64217, n64211, n72203, n64205, n61501, n72026, 
        n65059, n64199, n61483, n64193, n61481, n64187, n64181, 
        n29, n27, n64175, n23_adj_5852, n64169, n72023, n70961, 
        n64167, n17_adj_5853, n31_adj_5854, n16_adj_5855, n64163, 
        n64157, n64151, n65055, n64145, n69345, n64139, n64133, 
        n69315, n69299, n4_adj_5856, n64131, n64127, n69265, n59166, 
        n63545, n69259, n64121, n69251, n64115, n64109, n64103, 
        n64097, n64091, n64085, n64079, n63193, n61213, n61288, 
        n60896, n68468, n61134, n71402, n4_adj_5857, n68441, n68438, 
        n68433, n68429, n61442, n63212, n71233, n4_adj_5858, n68422, 
        n68421, n61461, n6_adj_5859, n5_adj_5860, n71482, n63843, 
        n63837, n63831, n72152, n63825, n68344, n63821, n63819, 
        n59920, n14_adj_5861, n10_adj_5862, n6_adj_5863, n9_adj_5864, 
        n70707, n71393, n6_adj_5865, n65633, n65630, n65063, n6_adj_5866, 
        n68285, n23_adj_5867, n12_adj_5868, n63691, n61245, n63635, 
        n8_adj_5869, n7_adj_5870, n65551, n65549, n65548, n6_adj_5871, 
        n68243;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27417), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i48542_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65632));
    defparam i48542_3_lut.LUT_INIT = 16'hcaca;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .GND_net(GND_net), 
            .state({state}), .timer({timer}), .VCC_net(VCC_net), .n29377(n29377), 
            .bit_ctr({Open_0, Open_1, Open_2, bit_ctr[1], Open_3}), 
            .n5(n5_adj_5860), .n29347(n29347), .t0({t0}), .n29346(n29346), 
            .n29345(n29345), .n27645(n27645), .n29344(n29344), .n29343(n29343), 
            .n29342(n29342), .n29341(n29341), .n29340(n29340), .n29339(n29339), 
            .n29338(n29338), .n35689(n35689), .\bit_ctr[0] (bit_ctr[0]), 
            .NEOPXL_c(NEOPXL_c), .n29126(n29126), .neopxl_color({neopxl_color}), 
            .LED_c(LED_c), .n39530(n39530), .n3172(n3172), .n23(n23_adj_5867)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_LUT4 LessThan_1178_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5829));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51685_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n68775));   // verilog/uart_rx.v(119[17:57])
    defparam i51685_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48543_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65633));
    defparam i48543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13344_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n28102), .I3(GND_net), .O(n29205));   // verilog/coms.v(130[12] 305[6])
    defparam i13344_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15_4_lut (.I0(\data_in_frame[18] [5]), .I1(n60419), .I2(n28117), 
            .I3(rx_data[5]), .O(n59922));   // verilog/coms.v(130[12] 305[6])
    defparam i15_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i13264_3_lut (.I0(b_prev_adj_5770), .I1(b_new_adj_5909[1]), 
            .I2(debounce_cnt_N_3833_adj_5771), .I3(GND_net), .O(n29125));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48540_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65630));
    defparam i48540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48539_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65629));
    defparam i48539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(n94), .I1(\FRAME_MATCHER.i [5]), .I2(n8_adj_5849), 
            .I3(n161), .O(n60419));
    defparam i5_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i15_4_lut_adj_1763 (.I0(\data_in_frame[18] [6]), .I1(n60419), 
            .I2(n28117), .I3(rx_data[6]), .O(n59920));   // verilog/coms.v(130[12] 305[6])
    defparam i15_4_lut_adj_1763.LUT_INIT = 16'hca0a;
    SB_LUT4 i51704_3_lut_4_lut (.I0(r_Clock_Count_adj_5945[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5945[2]), .O(n68794));   // verilog/uart_tx.v(117[17:57])
    defparam i51704_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i22170_4_lut (.I0(n68422), .I1(n68421), .I2(rx_data[7]), .I3(\data_in_frame[18] [7]), 
            .O(n37953));   // verilog/coms.v(94[13:20])
    defparam i22170_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22171_3_lut (.I0(n37953), .I1(\data_in_frame[18] [7]), .I2(reset), 
            .I3(GND_net), .O(n29513));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5724));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1181_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5945[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5822));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_91[7]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i18578_3_lut (.I0(n28102), .I1(rx_data[3]), .I2(\data_in_frame[11] [3]), 
            .I3(GND_net), .O(n29520));   // verilog/coms.v(94[13:20])
    defparam i18578_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 n9940_bdd_4_lut (.I0(n9940), .I1(current[15]), .I2(duty[22]), 
            .I3(n9938), .O(n72329));
    defparam n9940_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5723));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n72329_bdd_4_lut (.I0(n72329), .I1(duty[19]), .I2(n4918), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[19]));
    defparam n72329_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5722));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5721));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9940_bdd_4_lut_55150 (.I0(n9940), .I1(current[15]), .I2(duty[21]), 
            .I3(n9938), .O(n72323));
    defparam n9940_bdd_4_lut_55150.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5720));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n72323_bdd_4_lut (.I0(n72323), .I1(duty[18]), .I2(n4919), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[18]));
    defparam n72323_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5719));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9940_bdd_4_lut_55145 (.I0(n9940), .I1(current[15]), .I2(duty[20]), 
            .I3(n9938), .O(n72317));
    defparam n9940_bdd_4_lut_55145.LUT_INIT = 16'he4aa;
    SB_LUT4 n72317_bdd_4_lut (.I0(n72317), .I1(duty[17]), .I2(n4920), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[17]));
    defparam n72317_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13978_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n27465), .I3(GND_net), .O(n29839));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13979_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[1]), .I2(n5_adj_5763), 
            .I3(n25298), .O(n29840));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13979_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13281_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n28096), 
            .I3(GND_net), .O(n29142));   // verilog/coms.v(130[12] 305[6])
    defparam i13281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13278_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n28096), 
            .I3(GND_net), .O(n29139));   // verilog/coms.v(130[12] 305[6])
    defparam i13278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5718));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13982_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n27465), .I3(GND_net), .O(n29843));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13983_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n338), 
            .I2(n27465), .I3(GND_net), .O(n29844));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13984_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n27465), .I3(GND_net), .O(n29845));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18562_3_lut (.I0(n238), .I1(n290), .I2(n284), .I3(GND_net), 
            .O(n34394));
    defparam i18562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18563_3_lut (.I0(n34394), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n34395));
    defparam i18563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13338_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n28102), .I3(GND_net), .O(n29199));   // verilog/coms.v(130[12] 305[6])
    defparam i13338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n34395), .I2(n27465), 
            .I3(GND_net), .O(n29846));
    defparam i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13986_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n341), 
            .I2(n27465), .I3(GND_net), .O(n29847));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13987_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n27465), .I3(GND_net), .O(n29848));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5717));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13988_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n27465), .I3(GND_net), .O(n29849));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13989_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n27465), .I3(GND_net), .O(n29850));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9940_bdd_4_lut_55140 (.I0(n9940), .I1(current[15]), .I2(duty[19]), 
            .I3(n9938), .O(n72311));
    defparam n9940_bdd_4_lut_55140.LUT_INIT = 16'he4aa;
    SB_LUT4 i13990_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n27465), .I3(GND_net), .O(n29851));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13991_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n27465), .I3(GND_net), .O(n29852));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13992_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n27465), .I3(GND_net), .O(n29853));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13993_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n27465), .I3(GND_net), .O(n29854));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13994_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n27465), .I3(GND_net), .O(n29855));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54936 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[20] [0]), .I2(\data_out_frame[21] [0]), 
            .I3(byte_transmit_counter[2]), .O(n72053));
    defparam byte_transmit_counter_0__bdd_4_lut_54936.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n53828), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n72053_bdd_4_lut (.I0(n72053), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[2]), 
            .O(n72056));
    defparam n72053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13995_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n27465), .I3(GND_net), .O(n29856));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n72311_bdd_4_lut (.I0(n72311), .I1(duty[16]), .I2(n4921), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[16]));
    defparam n72311_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13996_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n27465), .I3(GND_net), .O(n29857));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13996_3_lut.LUT_INIT = 16'hcaca;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13997_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n27465), .I3(GND_net), .O(n29858));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13998_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n27465), .I3(GND_net), .O(n29859));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9940_bdd_4_lut_55135 (.I0(n9940), .I1(current[15]), .I2(duty[18]), 
            .I3(n9938), .O(n72305));
    defparam n9940_bdd_4_lut_55135.LUT_INIT = 16'he4aa;
    SB_LUT4 i13999_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n27465), .I3(GND_net), .O(n29860));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13999_3_lut.LUT_INIT = 16'hcaca;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n59166));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14000_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n27465), .I3(GND_net), .O(n29861));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_243_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_91[8]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14001_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n27465), .I3(GND_net), .O(n29862));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5716));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n53827), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n53827), .I0(GND_net), .I1(n2), 
            .CO(n53828));
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i14002_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n27465), .I3(GND_net), .O(n29863));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14003_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n27465), .I3(GND_net), .O(n29864));   // verilog/motorControl.v(42[14] 73[8])
    defparam i14003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14004_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[2]), .I2(n5_adj_5791), 
            .I3(n25298), .O(n29865));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14004_4_lut.LUT_INIT = 16'hccca;
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n53572), .O(n1240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14005_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[3]), .I2(n39133), 
            .I3(n25298), .O(n29866));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14005_4_lut.LUT_INIT = 16'hccac;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5715));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5713), 
            .I3(n53826), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(n23_adj_5852), .I1(o_Rx_DV_N_3488[12]), .I2(n5227), 
            .I3(r_SM_Main_adj_5944[0]), .O(n64235));
    defparam i1_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n64235), .O(n62322));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i13275_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n28096), 
            .I3(GND_net), .O(n29136));   // verilog/coms.v(130[12] 305[6])
    defparam i13275_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n53826), .I0(GND_net), .I1(n14_adj_5713), 
            .CO(n53827));
    SB_LUT4 n72305_bdd_4_lut (.I0(n72305), .I1(duty[15]), .I2(n4922), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[15]));
    defparam n72305_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14007_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[4]), .I2(n6_adj_5762), 
            .I3(n25289), .O(n29868));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14007_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13265_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3172), .I3(GND_net), 
            .O(n29126));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14008_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[5]), .I2(n6_adj_5762), 
            .I3(n25316), .O(n29869));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14008_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13272_3_lut (.I0(\data_in_frame[8] [4]), .I1(rx_data[4]), .I2(n28096), 
            .I3(GND_net), .O(n29133));   // verilog/coms.v(130[12] 305[6])
    defparam i13272_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i14010_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[6]), .I2(n6_adj_5762), 
            .I3(n25345), .O(n29871));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14010_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14011_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[7]), .I2(n6_adj_5762), 
            .I3(n25328), .O(n29872));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14011_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13269_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n28096), 
            .I3(GND_net), .O(n29130));   // verilog/coms.v(130[12] 305[6])
    defparam i13269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5714), 
            .I3(n53825), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i14013_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[8]), .I2(n6_adj_5761), 
            .I3(n25289), .O(n29874));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14013_4_lut.LUT_INIT = 16'hccca;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 i14014_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[9]), .I2(n6_adj_5761), 
            .I3(n25316), .O(n29875));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14014_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13266_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n28096), 
            .I3(GND_net), .O(n29127));   // verilog/coms.v(130[12] 305[6])
    defparam i13266_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n53825), .I0(GND_net), .I1(n15_adj_5714), 
            .CO(n53826));
    SB_LUT4 i14016_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[10]), .I2(n6_adj_5761), 
            .I3(n25345), .O(n29877));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14016_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14017_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[11]), .I2(n6_adj_5761), 
            .I3(n25328), .O(n29878));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14017_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14018_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[12]), .I2(n39146), 
            .I3(n25289), .O(n29879));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14018_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14019_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[15]), .I2(n39146), 
            .I3(n25328), .O(n29880));   // verilog/tli4970.v(35[10] 68[6])
    defparam i14019_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5715), 
            .I3(n53824), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9940_bdd_4_lut_55130 (.I0(n9940), .I1(current[15]), .I2(duty[17]), 
            .I3(n9938), .O(n72299));
    defparam n9940_bdd_4_lut_55130.LUT_INIT = 16'he4aa;
    SB_LUT4 n72299_bdd_4_lut (.I0(n72299), .I1(duty[14]), .I2(n4923), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[14]));
    defparam n72299_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55125 (.I0(n9940), .I1(current[15]), .I2(duty[16]), 
            .I3(n9938), .O(n72293));
    defparam n9940_bdd_4_lut_55125.LUT_INIT = 16'he4aa;
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 n72293_bdd_4_lut (.I0(n72293), .I1(duty[13]), .I2(n4924), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[13]));
    defparam n72293_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n53824), .I0(GND_net), .I1(n16_adj_5715), 
            .CO(n53825));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5716), 
            .I3(n53823), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14066_3_lut (.I0(\data_in_frame[2] [0]), .I1(rx_data[0]), .I2(n60766), 
            .I3(GND_net), .O(n29927));   // verilog/coms.v(130[12] 305[6])
    defparam i14066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14069_3_lut (.I0(\data_in_frame[2] [1]), .I1(rx_data[1]), .I2(n60766), 
            .I3(GND_net), .O(n29930));   // verilog/coms.v(130[12] 305[6])
    defparam i14069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14072_3_lut (.I0(\data_in_frame[2] [2]), .I1(rx_data[2]), .I2(n60766), 
            .I3(GND_net), .O(n29933));   // verilog/coms.v(130[12] 305[6])
    defparam i14072_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14075_3_lut (.I0(\data_in_frame[2] [3]), .I1(rx_data[3]), .I2(n60766), 
            .I3(GND_net), .O(n29936));   // verilog/coms.v(130[12] 305[6])
    defparam i14075_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n53823), .I0(GND_net), .I1(n17_adj_5716), 
            .CO(n53824));
    SB_LUT4 n9940_bdd_4_lut_55120 (.I0(n9940), .I1(current[15]), .I2(duty[15]), 
            .I3(n9938), .O(n72287));
    defparam n9940_bdd_4_lut_55120.LUT_INIT = 16'he4aa;
    SB_LUT4 i14078_3_lut (.I0(\data_in_frame[2] [4]), .I1(rx_data[4]), .I2(n60766), 
            .I3(GND_net), .O(n29939));   // verilog/coms.v(130[12] 305[6])
    defparam i14078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5714));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n72287_bdd_4_lut (.I0(n72287), .I1(duty[12]), .I2(n4925), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[12]));
    defparam n72287_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5713));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i11_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14081_3_lut (.I0(\data_in_frame[2] [5]), .I1(rx_data[5]), .I2(n60766), 
            .I3(GND_net), .O(n29942));   // verilog/coms.v(130[12] 305[6])
    defparam i14081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14084_3_lut (.I0(\data_in_frame[2] [6]), .I1(rx_data[6]), .I2(n60766), 
            .I3(GND_net), .O(n29945));   // verilog/coms.v(130[12] 305[6])
    defparam i14084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14087_3_lut (.I0(\data_in_frame[2] [7]), .I1(rx_data[7]), .I2(n60766), 
            .I3(GND_net), .O(n29948));   // verilog/coms.v(130[12] 305[6])
    defparam i14087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5717), 
            .I3(n53822), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n53822), .I0(GND_net), .I1(n18_adj_5717), 
            .CO(n53823));
    SB_CARRY add_151_14 (.CI(n53581), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n53582));
    SB_LUT4 n9940_bdd_4_lut_55115 (.I0(n9940), .I1(current[11]), .I2(duty[14]), 
            .I3(n9938), .O(n72281));
    defparam n9940_bdd_4_lut_55115.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5718), 
            .I3(n53821), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n72281_bdd_4_lut (.I0(n72281), .I1(duty[11]), .I2(n4926), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[11]));
    defparam n72281_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n53821), .I0(GND_net), .I1(n19_adj_5718), 
            .CO(n53822));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5719), 
            .I3(n53820), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9940_bdd_4_lut_55110 (.I0(n9940), .I1(current[10]), .I2(duty[13]), 
            .I3(n9938), .O(n72275));
    defparam n9940_bdd_4_lut_55110.LUT_INIT = 16'he4aa;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n53820), .I0(GND_net), .I1(n20_adj_5719), 
            .CO(n53821));
    SB_LUT4 n72275_bdd_4_lut (.I0(n72275), .I1(duty[10]), .I2(n4927), 
            .I3(n9938), .O(pwm_setpoint_23__N_3[10]));
    defparam n72275_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55105 (.I0(n9940), .I1(current[9]), .I2(duty[12]), 
            .I3(n9938), .O(n72269));
    defparam n9940_bdd_4_lut_55105.LUT_INIT = 16'he4aa;
    SB_LUT4 n72269_bdd_4_lut (.I0(n72269), .I1(duty[9]), .I2(n4928), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n72269_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55100 (.I0(n9940), .I1(current[8]), .I2(duty[11]), 
            .I3(n9938), .O(n72263));
    defparam n9940_bdd_4_lut_55100.LUT_INIT = 16'he4aa;
    SB_LUT4 n72263_bdd_4_lut (.I0(n72263), .I1(duty[8]), .I2(n4929), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n72263_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55095 (.I0(n9940), .I1(current[7]), .I2(duty[10]), 
            .I3(n9938), .O(n72257));
    defparam n9940_bdd_4_lut_55095.LUT_INIT = 16'he4aa;
    SB_LUT4 n72257_bdd_4_lut (.I0(n72257), .I1(duty[7]), .I2(n4930), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n72257_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55090 (.I0(n9940), .I1(current[6]), .I2(duty[9]), 
            .I3(n9938), .O(n72251));
    defparam n9940_bdd_4_lut_55090.LUT_INIT = 16'he4aa;
    SB_LUT4 n72251_bdd_4_lut (.I0(n72251), .I1(duty[6]), .I2(n4931), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n72251_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55085 (.I0(n9940), .I1(current[5]), .I2(duty[8]), 
            .I3(n9938), .O(n72245));
    defparam n9940_bdd_4_lut_55085.LUT_INIT = 16'he4aa;
    SB_LUT4 n72245_bdd_4_lut (.I0(n72245), .I1(duty[5]), .I2(n4932), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n72245_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55080 (.I0(n9940), .I1(current[4]), .I2(duty[7]), 
            .I3(n9938), .O(n72239));
    defparam n9940_bdd_4_lut_55080.LUT_INIT = 16'he4aa;
    SB_LUT4 n72239_bdd_4_lut (.I0(n72239), .I1(duty[4]), .I2(n4933), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n72239_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9940_bdd_4_lut_55075 (.I0(n9940), .I1(current[3]), .I2(duty[6]), 
            .I3(n9938), .O(n72233));
    defparam n9940_bdd_4_lut_55075.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_5838));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1765 (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5839));   // verilog/TinyFPGA_B.v(378[12:17])
    defparam i5_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i23238_4_lut (.I0(n13_adj_5839), .I1(baudrate[0]), .I2(n14_adj_5838), 
            .I3(n25296), .O(n39001));
    defparam i23238_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 i1_3_lut (.I0(n23_adj_5852), .I1(o_Rx_DV_N_3488[12]), .I2(n5227), 
            .I3(GND_net), .O(n63635));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63635), .O(r_SM_Main_2__N_3536[1]));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_1181_i9_2_lut (.I0(r_Clock_Count_adj_5945[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5824));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_243_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_91[9]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_1181_i13_2_lut (.I0(r_Clock_Count_adj_5945[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5826));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i11_2_lut (.I0(r_Clock_Count_adj_5945[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5825));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i15_2_lut (.I0(r_Clock_Count_adj_5945[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5827));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i4_4_lut (.I0(r_Clock_Count_adj_5945[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5945[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5821));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53716_3_lut (.I0(n4_adj_5821), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5825), 
            .I3(GND_net), .O(n70806));   // verilog/uart_tx.v(117[17:57])
    defparam i53716_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53717_3_lut (.I0(n70806), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5826), 
            .I3(GND_net), .O(n70807));   // verilog/uart_tx.v(117[17:57])
    defparam i53717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52667_4_lut (.I0(n13_adj_5826), .I1(n11_adj_5825), .I2(n9_adj_5824), 
            .I3(n68794), .O(n69757));
    defparam i52667_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1181_i8_3_lut (.I0(n6_adj_5822), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5824), .I3(GND_net), .O(n8_adj_5823));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52664_3_lut (.I0(n70807), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5827), 
            .I3(GND_net), .O(n69754));   // verilog/uart_tx.v(117[17:57])
    defparam i52664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53345_4_lut (.I0(n69754), .I1(n8_adj_5823), .I2(n15_adj_5827), 
            .I3(n69757), .O(n70435));   // verilog/uart_tx.v(117[17:57])
    defparam i53345_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53346_3_lut (.I0(n70435), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5945[8]), 
            .I3(GND_net), .O(n5227));   // verilog/uart_tx.v(117[17:57])
    defparam i53346_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1767 (.I0(o_Rx_DV_N_3488[12]), .I1(n5227), .I2(n60413), 
            .I3(GND_net), .O(n63825));
    defparam i1_3_lut_adj_1767.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n63825), .O(n63831));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5720), 
            .I3(n53819), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n53819), .I0(GND_net), .I1(n21_adj_5720), 
            .CO(n53820));
    SB_LUT4 n72233_bdd_4_lut (.I0(n72233), .I1(duty[3]), .I2(n4934), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n72233_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5721), 
            .I3(n53818), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n53818), .I0(GND_net), .I1(n22_adj_5721), 
            .CO(n53819));
    SB_LUT4 n9940_bdd_4_lut_55070 (.I0(n9940), .I1(current[2]), .I2(duty[5]), 
            .I3(n9938), .O(n72227));
    defparam n9940_bdd_4_lut_55070.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5722), 
            .I3(n53817), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n53817), .I0(GND_net), .I1(n23_adj_5722), 
            .CO(n53818));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5723), 
            .I3(n53816), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n53816), .I0(GND_net), .I1(n24_adj_5723), 
            .CO(n53817));
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n23_adj_5852), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5224), .I3(o_Rx_DV_N_3488[8]), .O(n63691));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n63691), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 i13640_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n28117), .I3(GND_net), .O(n29501));   // verilog/coms.v(130[12] 305[6])
    defparam i13640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n72227_bdd_4_lut (.I0(n72227), .I1(duty[2]), .I2(n4935), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n72227_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_1178_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5831));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1178_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5828));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1178_i8_3_lut (.I0(n6_adj_5829), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5831), .I3(GND_net), .O(n8_adj_5830));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54311_4_lut (.I0(n8_adj_5830), .I1(n4_adj_5828), .I2(n9_adj_5831), 
            .I3(n68775), .O(n71401));   // verilog/uart_rx.v(119[17:57])
    defparam i54311_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54312_3_lut (.I0(n71401), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n71402));   // verilog/uart_rx.v(119[17:57])
    defparam i54312_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54212_3_lut (.I0(n71402), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n71302));   // verilog/uart_rx.v(119[17:57])
    defparam i54212_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54037_3_lut (.I0(n71302), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5224));   // verilog/uart_rx.v(119[17:57])
    defparam i54037_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n60415), .O(n63837));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n39420), .I1(GND_net), .I2(n25_adj_5724), 
            .I3(VCC_net), .O(n68285)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n63837), .O(n63843));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5724), 
            .CO(n53816));
    SB_LUT4 n9940_bdd_4_lut_55065 (.I0(n9940), .I1(current[1]), .I2(duty[4]), 
            .I3(n9938), .O(n72221));
    defparam n9940_bdd_4_lut_55065.LUT_INIT = 16'he4aa;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n65629), .I2(n65630), .I3(byte_transmit_counter[1]), .O(n72023));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n72221_bdd_4_lut (.I0(n72221), .I1(duty[1]), .I2(n4936), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n72221_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n72023_bdd_4_lut (.I0(n72023), .I1(n65633), .I2(n65632), .I3(byte_transmit_counter[1]), 
            .O(n72026));
    defparam n72023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 dti_counter_2038_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n54439), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 dti_counter_2038_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n54438), .O(n39_adj_5832)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY dti_counter_2038_add_4_8 (.CI(n54438), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n54439));
    SB_LUT4 dti_counter_2038_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n54437), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY dti_counter_2038_add_4_7 (.CI(n54437), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n54438));
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_LUT4 dti_counter_2038_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n54436), .O(n41_adj_5833)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_6 (.CI(n54436), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n54437));
    SB_LUT4 dti_counter_2038_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n54435), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(321[10] 325[6])
    SB_CARRY dti_counter_2038_add_4_5 (.CI(n54435), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n54436));
    SB_DFFESR dti_counter_2038__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n27664), 
            .D(n45_adj_5835), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 n9940_bdd_4_lut_55060 (.I0(n9940), .I1(current[0]), .I2(duty[3]), 
            .I3(n9938), .O(n72215));
    defparam n9940_bdd_4_lut_55060.LUT_INIT = 16'he4aa;
    SB_LUT4 dti_counter_2038_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n54434), .O(n43_adj_5834)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_4 (.CI(n54434), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n54435));
    SB_LUT4 dti_counter_2038_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n54433), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n72215_bdd_4_lut (.I0(n72215), .I1(duty[0]), .I2(n4937), .I3(n9938), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n72215_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY dti_counter_2038_add_4_3 (.CI(n54433), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n54434));
    SB_LUT4 dti_counter_2038_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45_adj_5835)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n54433));
    SB_LUT4 i51585_4_lut (.I0(data_ready), .I1(n6910), .I2(n24_adj_5726), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n68438));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i51585_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i52196_2_lut (.I0(n24_adj_5726), .I1(n6910), .I2(GND_net), 
            .I3(GND_net), .O(n68441));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i52196_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n68441), .I1(n68438), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5863), .O(n59068));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55051 (.I0(byte_transmit_counter[3]), 
            .I1(n70707), .I2(n68433), .I3(byte_transmit_counter[4]), .O(n72203));
    defparam byte_transmit_counter_3__bdd_4_lut_55051.LUT_INIT = 16'he4aa;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/administrator/lscc/iCEcube2.2020.12/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n72203_bdd_4_lut (.I0(n72203), .I1(n72152), .I2(n7_adj_5840), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n72203_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5727));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i13813_4_lut (.I0(n63821), .I1(r_Bit_Index[0]), .I2(n61483), 
            .I3(n27511), .O(n29674));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13813_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i13810_4_lut (.I0(n63819), .I1(r_Bit_Index_adj_5946[0]), .I2(n61481), 
            .I3(n27514), .O(n29671));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13810_4_lut.LUT_INIT = 16'h32c8;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [4]), .I1(n60700), .I2(n28127), 
            .I3(rx_data[4]), .O(n59930));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_DFFESR dti_counter_2038__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27664), 
            .D(n38), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27664), 
            .D(n39_adj_5832), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27664), 
            .D(n40), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27664), 
            .D(n41_adj_5833), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27664), 
            .D(n42), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27664), 
            .D(n43_adj_5834), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_2038__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27664), 
            .D(n44), .R(n28828));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n63545));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n61501));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_91[4]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14_3_lut (.I0(hall2), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n6_adj_5871));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1773 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_1773.LUT_INIT = 16'h1414;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n53580), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27482), 
            .D(n1242), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i18867_4_lut_4_lut (.I0(PWMLimit[1]), .I1(setpoint[1]), .I2(setpoint[0]), 
            .I3(PWMLimit[0]), .O(n4_adj_5811));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i18867_4_lut_4_lut.LUT_INIT = 16'h44d4;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27482), 
            .D(n1241), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27482), 
            .D(n1240), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27482), 
            .D(n1239), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27482), 
            .D(n1238), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27482), 
            .D(n1237), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27482), 
            .D(n1236), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27482), 
            .D(n1235), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27482), 
            .D(n1234), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27482), 
            .D(n1233), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27482), 
            .D(n1232), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27482), 
            .D(n1231), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27482), 
            .D(n1230), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27482), 
            .D(n1229), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27482), 
            .D(n1228), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27482), 
            .D(n1243), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i12667_2_lut (.I0(n27441), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i12667_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27482), 
            .D(n1227), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i54470_4_lut (.I0(commutation_state[1]), .I1(n22661), .I2(dti), 
            .I3(commutation_state[2]), .O(n27441));
    defparam i54470_4_lut.LUT_INIT = 16'hc5cf;
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27482), 
            .D(n1226), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27482), 
            .D(n1225), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27482), 
            .D(n1224), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27482), 
            .D(n1223), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27482), 
            .D(n1222), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i9_2_lut (.I0(n290), .I1(n238), .I2(GND_net), .I3(GND_net), 
            .O(n39_adj_5817));
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27482), 
            .D(n1221), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27482), 
            .D(n1220), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27482), 
            .D(n1219), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27482), 
            .D(n1218), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27482), 
            .D(n1217), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27482), 
            .D(n1216), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27482), 
            .D(n1215), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27482), 
            .D(n1214), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27482), 
            .D(n1213), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27482), 
            .D(n1212), .R(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27441), .D(GHC_N_391), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27441), .D(GHB_N_377), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27441), .D(GHA_N_355), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n6_adj_5871), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27441), .D(GLA_N_372), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27441), .D(GLB_N_386), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27441), .D(GLC_N_400), 
            .R(n28534));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    GND i1 (.Y(GND_net));
    SB_CARRY add_151_13 (.CI(n53580), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n53581));
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5851));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1774 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5850));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5850), .I2(n10_adj_5851), 
            .I3(dti_counter[3]), .O(n22661));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5856));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'h7bde;
    SB_LUT4 i54713_2_lut (.I0(n22661), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i54713_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[16] [6]), .I3(GND_net), .O(n61134));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
           .D(n60302));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n59068));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    SB_LUT4 i12726_4_lut (.I0(n27482), .I1(n1323), .I2(n68344), .I3(n39100), 
            .O(n28543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i12726_4_lut.LUT_INIT = 16'ha088;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i2_2_lut_3_lut (.I0(hall1), .I1(hall3), .I2(hall2), .I3(GND_net), 
            .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n63545));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n53579), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_23_lut (.I0(GND_net), .I1(n13210), .I2(encoder1_position[25]), 
            .I3(n53964), .O(encoder1_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_22_lut (.I0(GND_net), .I1(n13211), .I2(encoder1_position[24]), 
            .I3(n53963), .O(encoder1_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_22 (.CI(n53963), .I0(n13211), .I1(encoder1_position[24]), 
            .CO(n53964));
    SB_LUT4 add_4773_21_lut (.I0(GND_net), .I1(n13212), .I2(encoder1_position[23]), 
            .I3(n53962), .O(encoder1_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_21 (.CI(n53962), .I0(n13212), .I1(encoder1_position[23]), 
            .CO(n53963));
    SB_LUT4 add_4773_20_lut (.I0(GND_net), .I1(n13213), .I2(encoder1_position[22]), 
            .I3(n53961), .O(encoder1_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_20 (.CI(n53961), .I0(n13213), .I1(encoder1_position[22]), 
            .CO(n53962));
    SB_LUT4 add_4773_19_lut (.I0(GND_net), .I1(n13214), .I2(encoder1_position[21]), 
            .I3(n53960), .O(encoder1_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_19 (.CI(n53960), .I0(n13214), .I1(encoder1_position[21]), 
            .CO(n53961));
    SB_LUT4 add_4773_18_lut (.I0(GND_net), .I1(n13215), .I2(encoder1_position[20]), 
            .I3(n53959), .O(encoder1_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_18 (.CI(n53959), .I0(n13215), .I1(encoder1_position[20]), 
            .CO(n53960));
    SB_LUT4 add_4773_17_lut (.I0(GND_net), .I1(n13216), .I2(encoder1_position[19]), 
            .I3(n53958), .O(encoder1_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_17 (.CI(n53958), .I0(n13216), .I1(encoder1_position[19]), 
            .CO(n53959));
    SB_LUT4 add_4773_16_lut (.I0(GND_net), .I1(n13217), .I2(encoder1_position[18]), 
            .I3(n53957), .O(encoder1_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_16 (.CI(n53957), .I0(n13217), .I1(encoder1_position[18]), 
            .CO(n53958));
    SB_LUT4 add_4773_15_lut (.I0(GND_net), .I1(n13218), .I2(encoder1_position[17]), 
            .I3(n53956), .O(encoder1_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_15 (.CI(n53956), .I0(n13218), .I1(encoder1_position[17]), 
            .CO(n53957));
    SB_LUT4 add_4773_14_lut (.I0(GND_net), .I1(n13219), .I2(encoder1_position[16]), 
            .I3(n53955), .O(encoder1_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_14 (.CI(n53955), .I0(n13219), .I1(encoder1_position[16]), 
            .CO(n53956));
    SB_LUT4 add_4773_13_lut (.I0(GND_net), .I1(n13220), .I2(encoder1_position[15]), 
            .I3(n53954), .O(encoder1_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_13 (.CI(n53954), .I0(n13220), .I1(encoder1_position[15]), 
            .CO(n53955));
    SB_LUT4 add_4773_12_lut (.I0(GND_net), .I1(n13221), .I2(encoder1_position[14]), 
            .I3(n53953), .O(encoder1_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_12 (.CI(n53953), .I0(n13221), .I1(encoder1_position[14]), 
            .CO(n53954));
    SB_LUT4 add_4773_11_lut (.I0(GND_net), .I1(n13222), .I2(encoder1_position[13]), 
            .I3(n53952), .O(encoder1_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13374_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29235));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13374_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4773_11 (.CI(n53952), .I0(n13222), .I1(encoder1_position[13]), 
            .CO(n53953));
    SB_LUT4 add_4773_10_lut (.I0(GND_net), .I1(n13223), .I2(encoder1_position[12]), 
            .I3(n53951), .O(encoder1_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n10003));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n11686));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i2_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4773_10 (.CI(n53951), .I0(n13223), .I1(encoder1_position[12]), 
            .CO(n53952));
    SB_LUT4 add_4773_9_lut (.I0(GND_net), .I1(n13224), .I2(encoder1_position[11]), 
            .I3(n53950), .O(encoder1_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_9 (.CI(n53950), .I0(n13224), .I1(encoder1_position[11]), 
            .CO(n53951));
    SB_LUT4 add_4773_8_lut (.I0(GND_net), .I1(n13225), .I2(encoder1_position[10]), 
            .I3(n53949), .O(encoder1_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n11684));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n11682));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i4_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4773_8 (.CI(n53949), .I0(n13225), .I1(encoder1_position[10]), 
            .CO(n53950));
    SB_CARRY add_151_5 (.CI(n53572), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n53573));
    SB_LUT4 i13376_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29237));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n11680));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n11678));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n11676));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n11674));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n11672));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n11670));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n11668));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n11666));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i12_3_lut.LUT_INIT = 16'h3535;
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1792(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .\a_new[1] (a_new[1]), 
            .\b_new[1] (b_new[1]), .n29238(n29238), .n1747(n1747), .n29237(n29237), 
            .a_prev(a_prev), .n29235(n29235), .b_prev(b_prev), .position_31__N_3836(position_31__N_3836), 
            .\encoder0_position[0] (encoder0_position[0]), .\encoder0_position[1] (encoder0_position[1]), 
            .\encoder0_position[2] (encoder0_position[2]), .\encoder0_position[3] (encoder0_position[3]), 
            .\encoder0_position[4] (encoder0_position[4]), .\encoder0_position[5] (encoder0_position[5]), 
            .\encoder0_position[6] (encoder0_position[6]), .\encoder0_position[7] (encoder0_position[7]), 
            .\encoder0_position[8] (encoder0_position[8]), .\encoder0_position[9] (encoder0_position[9]), 
            .\encoder0_position[10] (encoder0_position[10]), .\encoder0_position[11] (encoder0_position[11]), 
            .\encoder0_position[12] (encoder0_position[12]), .\encoder0_position[13] (encoder0_position[13]), 
            .\encoder0_position[14] (encoder0_position[14]), .\encoder0_position[15] (encoder0_position[15]), 
            .\encoder0_position[16] (encoder0_position[16]), .\encoder0_position[17] (encoder0_position[17]), 
            .\encoder0_position[18] (encoder0_position[18]), .\encoder0_position[19] (encoder0_position[19]), 
            .\encoder0_position[20] (encoder0_position[20]), .\encoder0_position[21] (encoder0_position[21]), 
            .\encoder0_position[22] (encoder0_position[22]), .n1765(n1765), 
            .n1763(n1763), .n1761(n1761), .n1759(n1759), .n1757(n1757), 
            .n1755(n1755), .n1753(n1753), .n1751(n1751), .n1749(n1749), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(305[27] 311[6])
    SB_LUT4 i13378_3_lut (.I0(a_prev_adj_5769), .I1(a_new_adj_5908[1]), 
            .I2(debounce_cnt_N_3833_adj_5771), .I3(GND_net), .O(n29239));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13378_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_12 (.CI(n53579), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n53580));
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n53578), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_7_lut (.I0(GND_net), .I1(n13226), .I2(encoder1_position[9]), 
            .I3(n53948), .O(encoder1_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n11664));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i13_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4773_7 (.CI(n53948), .I0(n13226), .I1(encoder1_position[9]), 
            .CO(n53949));
    SB_LUT4 add_4773_6_lut (.I0(GND_net), .I1(n13227), .I2(encoder1_position[8]), 
            .I3(n53947), .O(encoder1_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_6 (.CI(n53947), .I0(n13227), .I1(encoder1_position[8]), 
            .CO(n53948));
    SB_LUT4 add_4773_5_lut (.I0(GND_net), .I1(n13228), .I2(encoder1_position[7]), 
            .I3(n53946), .O(encoder1_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_5 (.CI(n53946), .I0(n13228), .I1(encoder1_position[7]), 
            .CO(n53947));
    SB_LUT4 add_4773_4_lut (.I0(GND_net), .I1(n13229), .I2(encoder1_position[6]), 
            .I3(n53945), .O(encoder1_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n11662));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n53571), .O(n1241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_11 (.CI(n53578), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n53579));
    SB_CARRY add_4773_4 (.CI(n53945), .I0(n13229), .I1(encoder1_position[6]), 
            .CO(n53946));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n53600), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4773_3_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[5]), 
            .I3(n53944), .O(encoder1_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_3 (.CI(n53944), .I0(encoder1_position[3]), .I1(encoder1_position[5]), 
            .CO(n53945));
    SB_LUT4 add_4773_2_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[4]), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4773_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4773_2 (.CI(GND_net), .I0(encoder1_position[2]), .I1(encoder1_position[4]), 
            .CO(n53944));
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n53599), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_32 (.CI(n53599), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n53600));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n53598), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n53598), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n53599));
    SB_LUT4 mux_1677_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n11660));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n53577), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n11658));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i16_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_151_4 (.CI(n53571), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n53572));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n53597), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4875_21_lut (.I0(GND_net), .I1(n15425), .I2(encoder1_position[23]), 
            .I3(n53934), .O(n13210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4875_20_lut (.I0(GND_net), .I1(n15426), .I2(encoder1_position[22]), 
            .I3(n53933), .O(n13211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_20 (.CI(n53933), .I0(n15426), .I1(encoder1_position[22]), 
            .CO(n53934));
    SB_LUT4 add_4875_19_lut (.I0(GND_net), .I1(n15427), .I2(encoder1_position[21]), 
            .I3(n53932), .O(n13212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_19 (.CI(n53932), .I0(n15427), .I1(encoder1_position[21]), 
            .CO(n53933));
    SB_LUT4 add_4875_18_lut (.I0(GND_net), .I1(n15428), .I2(encoder1_position[20]), 
            .I3(n53931), .O(n13213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n11656));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i17_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_151_30 (.CI(n53597), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n53598));
    SB_CARRY add_4875_18 (.CI(n53931), .I0(n15428), .I1(encoder1_position[20]), 
            .CO(n53932));
    SB_LUT4 add_4875_17_lut (.I0(GND_net), .I1(n15429), .I2(encoder1_position[19]), 
            .I3(n53930), .O(n13214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_17 (.CI(n53930), .I0(n15429), .I1(encoder1_position[19]), 
            .CO(n53931));
    SB_LUT4 add_4875_16_lut (.I0(GND_net), .I1(n15430), .I2(encoder1_position[18]), 
            .I3(n53929), .O(n13215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n11654));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i18_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4875_16 (.CI(n53929), .I0(n15430), .I1(encoder1_position[18]), 
            .CO(n53930));
    SB_LUT4 add_4875_15_lut (.I0(GND_net), .I1(n15431), .I2(encoder1_position[17]), 
            .I3(n53928), .O(n13216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_15 (.CI(n53928), .I0(n15431), .I1(encoder1_position[17]), 
            .CO(n53929));
    SB_LUT4 add_4875_14_lut (.I0(GND_net), .I1(n15432), .I2(encoder1_position[16]), 
            .I3(n53927), .O(n13217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_14 (.CI(n53927), .I0(n15432), .I1(encoder1_position[16]), 
            .CO(n53928));
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n53596), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4875_13_lut (.I0(GND_net), .I1(n15433), .I2(encoder1_position[15]), 
            .I3(n53926), .O(n13218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_13 (.CI(n53926), .I0(n15433), .I1(encoder1_position[15]), 
            .CO(n53927));
    SB_LUT4 add_4875_12_lut (.I0(GND_net), .I1(n15434), .I2(encoder1_position[14]), 
            .I3(n53925), .O(n13219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_12 (.CI(n53925), .I0(n15434), .I1(encoder1_position[14]), 
            .CO(n53926));
    SB_LUT4 add_4875_11_lut (.I0(GND_net), .I1(n15435), .I2(encoder1_position[13]), 
            .I3(n53924), .O(n13220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_11 (.CI(n53924), .I0(n15435), .I1(encoder1_position[13]), 
            .CO(n53925));
    SB_LUT4 add_4875_10_lut (.I0(GND_net), .I1(n15436), .I2(encoder1_position[12]), 
            .I3(n53923), .O(n13221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n11652));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i19_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4875_10 (.CI(n53923), .I0(n15436), .I1(encoder1_position[12]), 
            .CO(n53924));
    SB_LUT4 add_4875_9_lut (.I0(GND_net), .I1(n15437), .I2(encoder1_position[11]), 
            .I3(n53922), .O(n13222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n11650));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i20_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4875_9 (.CI(n53922), .I0(n15437), .I1(encoder1_position[11]), 
            .CO(n53923));
    SB_LUT4 add_4875_8_lut (.I0(GND_net), .I1(n15438), .I2(encoder1_position[10]), 
            .I3(n53921), .O(n13223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_8 (.CI(n53921), .I0(n15438), .I1(encoder1_position[10]), 
            .CO(n53922));
    SB_LUT4 add_4875_7_lut (.I0(GND_net), .I1(n15439), .I2(encoder1_position[9]), 
            .I3(n53920), .O(n13224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_7 (.CI(n53920), .I0(n15439), .I1(encoder1_position[9]), 
            .CO(n53921));
    SB_LUT4 add_4875_6_lut (.I0(GND_net), .I1(n15440), .I2(encoder1_position[8]), 
            .I3(n53919), .O(n13225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_6 (.CI(n53919), .I0(n15440), .I1(encoder1_position[8]), 
            .CO(n53920));
    SB_LUT4 add_4875_5_lut (.I0(GND_net), .I1(n15441), .I2(encoder1_position[7]), 
            .I3(n53918), .O(n13226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n11648));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5776), .I3(n53746), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_5 (.CI(n53918), .I0(n15441), .I1(encoder1_position[7]), 
            .CO(n53919));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3), .I3(n53745), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4875_4_lut (.I0(GND_net), .I1(n15442), .I2(encoder1_position[6]), 
            .I3(n53917), .O(n13227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n11646));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i22_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n53745), .I0(encoder0_position_scaled[22]), 
            .I1(n3), .CO(n53746));
    SB_CARRY add_4875_4 (.CI(n53917), .I0(n15442), .I1(encoder1_position[6]), 
            .CO(n53918));
    SB_LUT4 add_4875_3_lut (.I0(GND_net), .I1(n15443), .I2(encoder1_position[5]), 
            .I3(n53916), .O(n13228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4875_3 (.CI(n53916), .I0(n15443), .I1(encoder1_position[5]), 
            .CO(n53917));
    SB_LUT4 add_4875_2_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[4]), 
            .I3(GND_net), .O(n13229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4875_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n11644));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1677_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5775), .I3(n53744), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n53744), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5775), .CO(n53745));
    SB_CARRY add_4875_2 (.CI(GND_net), .I0(encoder1_position[2]), .I1(encoder1_position[4]), 
            .CO(n53916));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5796), .I3(n53743), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n53743), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5796), .CO(n53744));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5795), .I3(n53742), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n53742), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5795), .CO(n53743));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5794), .I3(n53741), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n53741), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5794), .CO(n53742));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5793), .I3(n53740), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n53740), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5793), .CO(n53741));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5792), .I3(n53739), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n53739), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5792), .CO(n53740));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5774), .I3(n53738), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n53738), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5774), .CO(n53739));
    SB_CARRY add_151_29 (.CI(n53596), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n53597));
    SB_CARRY add_151_10 (.CI(n53577), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n53578));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5773), .I3(n53737), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n53737), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5773), .CO(n53738));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n53595), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n53570), .O(n1242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12), .I3(n53736), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n53736), .I0(encoder0_position_scaled[13]), 
            .I1(n12), .CO(n53737));
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n53576), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5712), .I3(n53735), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n53735), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5712), .CO(n53736));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n53734), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n53734), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n53735));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5711), .I3(n53733), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n53733), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5711), .CO(n53734));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5710), .I3(n53732), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n53732), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5710), .CO(n53733));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5709), .I3(n53731), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_28 (.CI(n53595), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n53596));
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n53594), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n53731), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5709), .CO(n53732));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18), .I3(n53730), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n53730), .I0(encoder0_position_scaled[7]), 
            .I1(n18), .CO(n53731));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n53729), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n53729), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n53730));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n53728), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n53728), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n53729));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n53727), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n53727), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n53728));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n53726), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n53726), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n53727));
    SB_CARRY add_151_27 (.CI(n53594), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n53595));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n53725), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n53725), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n53726));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n53593), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n53724), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n53724), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n53725));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25), .CO(n53724));
    SB_CARRY add_151_26 (.CI(n53593), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n53594));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n53592), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_9 (.CI(n53576), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n53577));
    SB_CARRY add_151_25 (.CI(n53592), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n53593));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n53591), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_24 (.CI(n53591), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n53592));
    SB_CARRY add_151_3 (.CI(n53570), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n53571));
    SB_LUT4 add_4873_20_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(encoder1_position[21]), 
            .I3(n53884), .O(n15425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_19_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(encoder1_position[20]), 
            .I3(n53883), .O(n15426)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_19 (.CI(n53883), .I0(encoder1_position[19]), .I1(encoder1_position[20]), 
            .CO(n53884));
    SB_LUT4 add_4873_18_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(encoder1_position[19]), 
            .I3(n53882), .O(n15427)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_18 (.CI(n53882), .I0(encoder1_position[18]), .I1(encoder1_position[19]), 
            .CO(n53883));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n53575), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_17_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(encoder1_position[18]), 
            .I3(n53881), .O(n15428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_17 (.CI(n53881), .I0(encoder1_position[17]), .I1(encoder1_position[18]), 
            .CO(n53882));
    SB_LUT4 add_4873_16_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(encoder1_position[17]), 
            .I3(n53880), .O(n15429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_16 (.CI(n53880), .I0(encoder1_position[16]), .I1(encoder1_position[17]), 
            .CO(n53881));
    SB_LUT4 add_4873_15_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(encoder1_position[16]), 
            .I3(n53879), .O(n15430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_15 (.CI(n53879), .I0(encoder1_position[15]), .I1(encoder1_position[16]), 
            .CO(n53880));
    SB_LUT4 add_4873_14_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(encoder1_position[15]), 
            .I3(n53878), .O(n15431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_14 (.CI(n53878), .I0(encoder1_position[14]), .I1(encoder1_position[15]), 
            .CO(n53879));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n53590), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_13_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(encoder1_position[14]), 
            .I3(n53877), .O(n15432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n53590), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n53591));
    SB_CARRY add_4873_13 (.CI(n53877), .I0(encoder1_position[13]), .I1(encoder1_position[14]), 
            .CO(n53878));
    SB_LUT4 add_4873_12_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(encoder1_position[13]), 
            .I3(n53876), .O(n15433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_12 (.CI(n53876), .I0(encoder1_position[12]), .I1(encoder1_position[13]), 
            .CO(n53877));
    SB_LUT4 add_4873_11_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(encoder1_position[12]), 
            .I3(n53875), .O(n15434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_11 (.CI(n53875), .I0(encoder1_position[11]), .I1(encoder1_position[12]), 
            .CO(n53876));
    SB_LUT4 add_4873_10_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(encoder1_position[11]), 
            .I3(n53874), .O(n15435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_10 (.CI(n53874), .I0(encoder1_position[10]), .I1(encoder1_position[11]), 
            .CO(n53875));
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n53589), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_9_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(encoder1_position[10]), 
            .I3(n53873), .O(n15436)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_8 (.CI(n53575), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n53576));
    SB_CARRY add_151_22 (.CI(n53589), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n53590));
    SB_CARRY add_4873_9 (.CI(n53873), .I0(encoder1_position[9]), .I1(encoder1_position[10]), 
            .CO(n53874));
    SB_LUT4 add_4873_8_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(encoder1_position[9]), 
            .I3(n53872), .O(n15437)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_8 (.CI(n53872), .I0(encoder1_position[8]), .I1(encoder1_position[9]), 
            .CO(n53873));
    SB_LUT4 add_4873_7_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(encoder1_position[8]), 
            .I3(n53871), .O(n15438)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_7 (.CI(n53871), .I0(encoder1_position[7]), .I1(encoder1_position[8]), 
            .CO(n53872));
    SB_LUT4 add_4873_6_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(encoder1_position[7]), 
            .I3(n53870), .O(n15439)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_6 (.CI(n53870), .I0(encoder1_position[6]), .I1(encoder1_position[7]), 
            .CO(n53871));
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n53588), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n53574), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_5_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(encoder1_position[6]), 
            .I3(n53869), .O(n15440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_21 (.CI(n53588), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n53589));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n53587), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_20 (.CI(n53587), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n53588));
    SB_CARRY add_4873_5 (.CI(n53869), .I0(encoder1_position[5]), .I1(encoder1_position[6]), 
            .CO(n53870));
    SB_LUT4 add_4873_4_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(encoder1_position[5]), 
            .I3(n53868), .O(n15441)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_4 (.CI(n53868), .I0(encoder1_position[4]), .I1(encoder1_position[5]), 
            .CO(n53869));
    SB_LUT4 add_4873_3_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[4]), 
            .I3(n53867), .O(n15442)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_3 (.CI(n53867), .I0(encoder1_position[3]), .I1(encoder1_position[4]), 
            .CO(n53868));
    SB_LUT4 add_1190_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n53692), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4873_2_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[3]), 
            .I3(GND_net), .O(n15443)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4873_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_24_lut (.I0(GND_net), .I1(GND_net), .I2(n11644), 
            .I3(n53691), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4873_2 (.CI(GND_net), .I0(encoder1_position[2]), .I1(encoder1_position[3]), 
            .CO(n53867));
    SB_CARRY add_1190_24 (.CI(n53691), .I0(GND_net), .I1(n11644), .CO(n53692));
    SB_LUT4 add_1190_23_lut (.I0(GND_net), .I1(GND_net), .I2(n11646), 
            .I3(n53690), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_23 (.CI(n53690), .I0(GND_net), .I1(n11646), .CO(n53691));
    SB_LUT4 add_1190_22_lut (.I0(GND_net), .I1(GND_net), .I2(n11648), 
            .I3(n53689), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_22 (.CI(n53689), .I0(GND_net), .I1(n11648), .CO(n53690));
    SB_LUT4 add_1190_21_lut (.I0(GND_net), .I1(GND_net), .I2(n11650), 
            .I3(n53688), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_21 (.CI(n53688), .I0(GND_net), .I1(n11650), .CO(n53689));
    SB_LUT4 add_1190_20_lut (.I0(GND_net), .I1(GND_net), .I2(n11652), 
            .I3(n53687), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_20 (.CI(n53687), .I0(GND_net), .I1(n11652), .CO(n53688));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n53586), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_19_lut (.I0(GND_net), .I1(GND_net), .I2(n11654), 
            .I3(n53686), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_19 (.CI(n53686), .I0(GND_net), .I1(n11654), .CO(n53687));
    SB_CARRY add_151_19 (.CI(n53586), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n53587));
    SB_LUT4 add_1190_18_lut (.I0(GND_net), .I1(GND_net), .I2(n11656), 
            .I3(n53685), .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_18 (.CI(n53685), .I0(GND_net), .I1(n11656), .CO(n53686));
    SB_LUT4 add_1190_17_lut (.I0(GND_net), .I1(GND_net), .I2(n11658), 
            .I3(n53684), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_17 (.CI(n53684), .I0(GND_net), .I1(n11658), .CO(n53685));
    SB_LUT4 add_1190_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11660), 
            .I3(n53683), .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_16 (.CI(n53683), .I0(GND_net), .I1(n11660), .CO(n53684));
    SB_LUT4 add_1190_15_lut (.I0(GND_net), .I1(GND_net), .I2(n11662), 
            .I3(n53682), .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_15 (.CI(n53682), .I0(GND_net), .I1(n11662), .CO(n53683));
    SB_LUT4 add_1190_14_lut (.I0(GND_net), .I1(GND_net), .I2(n11664), 
            .I3(n53681), .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13263_3_lut_4_lut (.I0(n1797), .I1(b_prev_adj_5770), .I2(a_new_adj_5908[1]), 
            .I3(position_31__N_3836_adj_5772), .O(n29124));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13263_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_CARRY add_1190_14 (.CI(n53681), .I0(GND_net), .I1(n11664), .CO(n53682));
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n53585), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1190_13_lut (.I0(GND_net), .I1(GND_net), .I2(n11666), 
            .I3(n53680), .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_13 (.CI(n53680), .I0(GND_net), .I1(n11666), .CO(n53681));
    SB_CARRY add_151_18 (.CI(n53585), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n53586));
    SB_LUT4 add_1190_12_lut (.I0(GND_net), .I1(GND_net), .I2(n11668), 
            .I3(n53679), .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_12 (.CI(n53679), .I0(GND_net), .I1(n11668), .CO(n53680));
    SB_LUT4 add_1190_11_lut (.I0(GND_net), .I1(GND_net), .I2(n11670), 
            .I3(n53678), .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_11 (.CI(n53678), .I0(GND_net), .I1(n11670), .CO(n53679));
    SB_LUT4 add_1190_10_lut (.I0(GND_net), .I1(GND_net), .I2(n11672), 
            .I3(n53677), .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_10 (.CI(n53677), .I0(GND_net), .I1(n11672), .CO(n53678));
    SB_LUT4 add_1190_9_lut (.I0(GND_net), .I1(GND_net), .I2(n11674), .I3(n53676), 
            .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_9 (.CI(n53676), .I0(GND_net), .I1(n11674), .CO(n53677));
    SB_LUT4 add_1190_8_lut (.I0(GND_net), .I1(GND_net), .I2(n11676), .I3(n53675), 
            .O(n4931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_7 (.CI(n53574), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n53575));
    SB_CARRY add_1190_8 (.CI(n53675), .I0(GND_net), .I1(n11676), .CO(n53676));
    SB_LUT4 add_1190_7_lut (.I0(GND_net), .I1(GND_net), .I2(n11678), .I3(n53674), 
            .O(n4932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n53584), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n53570));
    SB_CARRY add_1190_7 (.CI(n53674), .I0(GND_net), .I1(n11678), .CO(n53675));
    SB_LUT4 add_1190_6_lut (.I0(GND_net), .I1(GND_net), .I2(n11680), .I3(n53673), 
            .O(n4933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n53573), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_6 (.CI(n53673), .I0(GND_net), .I1(n11680), .CO(n53674));
    SB_LUT4 add_1190_5_lut (.I0(GND_net), .I1(GND_net), .I2(n11682), .I3(n53672), 
            .O(n4934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n53584), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n53585));
    SB_CARRY add_1190_5 (.CI(n53672), .I0(GND_net), .I1(n11682), .CO(n53673));
    SB_LUT4 add_1190_4_lut (.I0(GND_net), .I1(GND_net), .I2(n11684), .I3(n53671), 
            .O(n4935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_4 (.CI(n53671), .I0(GND_net), .I1(n11684), .CO(n53672));
    SB_LUT4 add_1190_3_lut (.I0(GND_net), .I1(GND_net), .I2(n11686), .I3(n53670), 
            .O(n4936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_3 (.CI(n53670), .I0(GND_net), .I1(n11686), .CO(n53671));
    SB_LUT4 add_1190_2_lut (.I0(GND_net), .I1(GND_net), .I2(n10003), .I3(VCC_net), 
            .O(n4937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n53583), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_2 (.CI(VCC_net), .I0(GND_net), .I1(n10003), .CO(n53670));
    SB_CARRY add_151_6 (.CI(n53573), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n53574));
    SB_CARRY add_151_16 (.CI(n53583), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n53584));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n53582), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n53582), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n53583));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n53581), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13262_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5944[1]), 
            .I2(r_SM_Main_adj_5944[2]), .I3(n6_adj_5846), .O(n29123));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13262_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_LUT4 i1_2_lut_3_lut (.I0(n37935), .I1(reset), .I2(n39431), .I3(GND_net), 
            .O(n37938));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i23665_2_lut_3_lut (.I0(n3483), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n39431));
    defparam i23665_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i13752_3_lut_4_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(n37938), .I3(n39467), .O(n29613));   // verilog/coms.v(130[12] 305[6])
    defparam i13752_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut (.I0(n34395), .I1(Ki[2]), .I2(GND_net), .I3(GND_net), 
            .O(n204));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1776 (.I0(n34395), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n131));
    defparam i1_2_lut_adj_1776.LUT_INIT = 16'h8888;
    SB_LUT4 i5240_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5240_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i5238_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i5238_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i5242_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i5242_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5244_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i5244_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2828), .O(n25_adj_5820));   // verilog/TinyFPGA_B.v(377[7:11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5709));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5710));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5711));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5712));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5773));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_91[10]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n39431), .I3(n110), .O(n60));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5774));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5792));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22689_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(n1_adj_5843));
    defparam i22689_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22690_3_lut (.I0(encoder0_position_scaled[11]), .I1(n1_adj_5843), 
            .I2(n15_adj_5766), .I3(GND_net), .O(n3_adj_5841));
    defparam i22690_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5793));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_91[12]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5794));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51799_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n39431), .I3(n37941), .O(n68421));
    defparam i51799_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5795));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_91[13]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5796));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_91[14]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5775));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5776));   // verilog/TinyFPGA_B.v(324[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_91[15]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_91[16]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5755));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_91[17]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_243_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_91[18]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_91[19]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5753));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_4_lut_adj_1777 (.I0(n260), .I1(n65191), .I2(duty[23]), 
            .I3(n22_adj_5845), .O(n9938));
    defparam i1_4_lut_4_lut_adj_1777.LUT_INIT = 16'h1505;
    SB_LUT4 i52209_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n69299));
    defparam i52209_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_91[20]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_91[21]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i37054_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[22]));
    defparam i37054_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5741));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_243_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_91[22]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i52161_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n69251));
    defparam i52161_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i17_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(n16_adj_5855));
    defparam i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i18_3_lut (.I0(encoder0_position_scaled[23]), .I1(n16_adj_5855), 
            .I2(n15_adj_5766), .I3(GND_net), .O(n17_adj_5853));
    defparam i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5739));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52411_2_lut (.I0(displacement[0]), .I1(n15_adj_5790), .I2(GND_net), 
            .I3(GND_net), .O(n68243));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam i52411_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_91[1]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_91[2]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_91[3]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13619_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29480));
    defparam i13619_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13602_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29463));
    defparam i13602_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13616_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29477));
    defparam i13616_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13599_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29460));
    defparam i13599_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13612_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29473));
    defparam i13612_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13449_3_lut (.I0(current[11]), .I1(data_adj_5928[11]), .I2(n27489), 
            .I3(GND_net), .O(n29310));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1778 (.I0(\data_out_frame[10] [6]), .I1(n56545), 
            .I2(n26215), .I3(GND_net), .O(n61245));
    defparam i1_2_lut_3_lut_adj_1778.LUT_INIT = 16'h6969;
    SB_LUT4 i13625_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29486));
    defparam i13625_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13450_3_lut (.I0(current[10]), .I1(data_adj_5928[10]), .I2(n27489), 
            .I3(GND_net), .O(n29311));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54981 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n72119));
    defparam byte_transmit_counter_0__bdd_4_lut_54981.LUT_INIT = 16'he4aa;
    SB_LUT4 i13622_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29483));
    defparam i13622_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13605_3_lut_4_lut (.I0(n37938), .I1(n8_adj_5810), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29466));
    defparam i13605_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i52048_3_lut_4_lut (.I0(state_7__N_4110[0]), .I1(n10_adj_5760), 
            .I2(state_adj_5954[0]), .I3(enable_slow_N_4213), .O(n68468));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i52048_3_lut_4_lut.LUT_INIT = 16'h54fc;
    SB_LUT4 i13451_3_lut (.I0(current[9]), .I1(data_adj_5928[9]), .I2(n27489), 
            .I3(GND_net), .O(n29312));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n72119_bdd_4_lut (.I0(n72119), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n72122));
    defparam n72119_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13516_4_lut_4_lut (.I0(n27645), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n29377));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13516_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i13452_3_lut (.I0(current[8]), .I1(data_adj_5928[8]), .I2(n27489), 
            .I3(GND_net), .O(n29313));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(n56501), .I1(\data_out_frame[16] [4]), .I2(n60951), 
            .I3(n6_adj_5859), .O(n24820));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13453_3_lut (.I0(current[7]), .I1(data_adj_5928[7]), .I2(n27489), 
            .I3(GND_net), .O(n29314));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1956_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1323), .I3(n39001), .O(n6910));   // verilog/TinyFPGA_B.v(362[5] 388[12])
    defparam i1956_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i13454_3_lut (.I0(current[6]), .I1(data_adj_5928[6]), .I2(n27489), 
            .I3(GND_net), .O(n29315));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13455_3_lut (.I0(current[5]), .I1(data_adj_5928[5]), .I2(n27489), 
            .I3(GND_net), .O(n29316));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13456_3_lut (.I0(current[4]), .I1(data_adj_5928[4]), .I2(n27489), 
            .I3(GND_net), .O(n29317));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13457_3_lut (.I0(current[3]), .I1(data_adj_5928[3]), .I2(n27489), 
            .I3(GND_net), .O(n29318));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13458_3_lut (.I0(current[2]), .I1(data_adj_5928[2]), .I2(n27489), 
            .I3(GND_net), .O(n29319));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13459_3_lut (.I0(current[1]), .I1(data_adj_5928[1]), .I2(n27489), 
            .I3(GND_net), .O(n29320));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13460_3_lut (.I0(baudrate[31]), .I1(data_adj_5921[7]), .I2(n63193), 
            .I3(GND_net), .O(n29321));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13460_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main[0]), .O(n64167));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i13461_3_lut (.I0(baudrate[30]), .I1(data_adj_5921[6]), .I2(n63193), 
            .I3(GND_net), .O(n29322));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_4_lut_adj_1779 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_Bit_Index[0]), .O(n64131));
    defparam i1_3_lut_4_lut_adj_1779.LUT_INIT = 16'hffef;
    SB_LUT4 i3_4_lut_adj_1780 (.I0(n61134), .I1(n56696), .I2(\data_in_frame[17] [0]), 
            .I3(n56640), .O(n56565));
    defparam i3_4_lut_adj_1780.LUT_INIT = 16'h6996;
    SB_LUT4 i13462_3_lut (.I0(baudrate[29]), .I1(data_adj_5921[5]), .I2(n63193), 
            .I3(GND_net), .O(n29323));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13463_3_lut (.I0(baudrate[28]), .I1(data_adj_5921[4]), .I2(n63193), 
            .I3(GND_net), .O(n29324));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13464_3_lut (.I0(baudrate[27]), .I1(data_adj_5921[3]), .I2(n63193), 
            .I3(GND_net), .O(n29325));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13465_3_lut (.I0(baudrate[26]), .I1(data_adj_5921[2]), .I2(n63193), 
            .I3(GND_net), .O(n29326));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13466_3_lut (.I0(baudrate[25]), .I1(data_adj_5921[1]), .I2(n63193), 
            .I3(GND_net), .O(n29327));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13467_3_lut (.I0(baudrate[24]), .I1(data_adj_5921[0]), .I2(n63193), 
            .I3(GND_net), .O(n29328));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1781 (.I0(\data_out_frame[5] [2]), .I1(n31_adj_5842), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5862));
    defparam i2_2_lut_adj_1781.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1782 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[5] [4]), 
            .I2(n61210), .I3(n55578), .O(n14_adj_5861));
    defparam i6_4_lut_adj_1782.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1783 (.I0(\data_out_frame[14] [1]), .I1(n14_adj_5861), 
            .I2(n10_adj_5862), .I3(n61288), .O(n62686));
    defparam i7_4_lut_adj_1783.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n60534));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1784 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n60533));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1784.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1785 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n60532));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1785.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1786 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n60531));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1786.LUT_INIT = 16'h2300;
    SB_LUT4 i13477_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3172), .I3(GND_net), 
            .O(n29338));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1787 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n28930));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1787.LUT_INIT = 16'h2300;
    SB_LUT4 i13478_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3172), .I3(GND_net), 
            .O(n29339));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1788 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n60530));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1788.LUT_INIT = 16'h2300;
    SB_LUT4 i13479_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3172), .I3(GND_net), 
            .O(n29340));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1789 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n60474));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1789.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1790 (.I0(n55945), .I1(n61213), .I2(GND_net), 
            .I3(GND_net), .O(n56624));
    defparam i1_2_lut_adj_1790.LUT_INIT = 16'h6666;
    SB_LUT4 i13480_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3172), .I3(GND_net), 
            .O(n29341));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1791 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n60529));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1791.LUT_INIT = 16'h2300;
    SB_LUT4 i13481_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3172), .I3(GND_net), 
            .O(n29342));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13482_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3172), .I3(GND_net), 
            .O(n29343));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1792 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n60528));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1792.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n60527));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1793.LUT_INIT = 16'h2300;
    SB_LUT4 i13483_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3172), .I3(GND_net), 
            .O(n29344));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1794 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n60526));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1794.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1795 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n60525));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1795.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1796 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n60524));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1796.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1797 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n60523));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1797.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1798 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n60522));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1798.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1799 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n60476));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1799.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1800 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n60521));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1800.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1801 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n60520));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1801.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1802 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n60519));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1802.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1803 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n60646));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1803.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1804 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n60645));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1804.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1805 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n60644));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1805.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1806 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n60643));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1806.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1807 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n60642));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1807.LUT_INIT = 16'h2300;
    SB_LUT4 i13332_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n28102), .I3(GND_net), .O(n29193));   // verilog/coms.v(130[12] 305[6])
    defparam i13332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1808 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n60658));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1808.LUT_INIT = 16'h2300;
    SB_LUT4 i13484_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3172), .I3(GND_net), 
            .O(n29345));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_91[5]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n60641));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n60518));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1811 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n60517));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1811.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1812 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n60516));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1812.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n60515));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 i48461_3_lut (.I0(n4917), .I1(duty[20]), .I2(n9940), .I3(GND_net), 
            .O(n65551));
    defparam i48461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48463_3_lut (.I0(n65551), .I1(n65549), .I2(n9938), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i48463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48458_3_lut (.I0(n4916), .I1(duty[21]), .I2(n9940), .I3(GND_net), 
            .O(n65548));
    defparam i48458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48460_3_lut (.I0(n65548), .I1(n65549), .I2(n9938), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i48460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48459_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n9940), 
            .I3(GND_net), .O(n65549));
    defparam i48459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48455_3_lut (.I0(n4915), .I1(duty[22]), .I2(n9940), .I3(GND_net), 
            .O(n65545));
    defparam i48455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n60514));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 i48457_3_lut (.I0(n65545), .I1(n65549), .I2(n9938), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i48457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n60513));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 i5892_3_lut (.I0(n4914), .I1(current[15]), .I2(n9938), .I3(GND_net), 
            .O(n21407));
    defparam i5892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1816 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n60512));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1816.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1817 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n60511));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1817.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1818 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n60510));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1818.LUT_INIT = 16'h2300;
    SB_LUT4 i5893_3_lut (.I0(n21407), .I1(duty[23]), .I2(n9940), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i5893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13485_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3172), .I3(GND_net), 
            .O(n29346));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13486_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3172), .I3(GND_net), 
            .O(n29347));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1819 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n60509));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1819.LUT_INIT = 16'h2300;
    SB_LUT4 i17_2_lut (.I0(n31_adj_5842), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26311));   // verilog/coms.v(100[12:26])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1820 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n61210));
    defparam i1_2_lut_adj_1820.LUT_INIT = 16'h6666;
    SB_LUT4 i13236_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n27465), .I3(GND_net), .O(n29097));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n60508));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1822 (.I0(r_SM_Main[1]), .I1(n6_adj_5866), .I2(r_Bit_Index[0]), 
            .I3(n4_adj_5759), .O(n64187));
    defparam i1_4_lut_adj_1822.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n60507));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1824 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64187), .O(n64193));
    defparam i1_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64193), .O(n64199));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i13778_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n64199), 
            .I3(n27), .O(n29639));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13778_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1826 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n60506));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1826.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64133), .O(n64139));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1828 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n60505));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1828.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1829 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64139), .O(n64145));
    defparam i1_4_lut_adj_1829.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n60504));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_LUT4 i13779_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n64145), 
            .I3(n27), .O(n29640));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13779_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n60503));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64097), .O(n64103));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64103), .O(n64109));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i13780_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n64109), 
            .I3(n27), .O(n29641));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13780_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n60502));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n60501));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1836 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n60500));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1836.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1837 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n60499));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1837.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_1838 (.I0(n56501), .I1(n61461), .I2(\data_out_frame[18] [6]), 
            .I3(n25712), .O(n55945));
    defparam i3_4_lut_adj_1838.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1839 (.I0(\data_out_frame[18] [7]), .I1(n25994), 
            .I2(GND_net), .I3(GND_net), .O(n61442));
    defparam i1_2_lut_adj_1839.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n60640));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n60639));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1842 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1842.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n60638));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1844 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64151), .O(n64157));
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1845 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64157), .O(n64163));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i13781_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n64163), 
            .I3(n27), .O(n29642));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13781_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n60498));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n60497));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n60496));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n60495));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64169), .O(n64175));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1851 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64175), .O(n64181));
    defparam i1_4_lut_adj_1851.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1852 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n60494));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1852.LUT_INIT = 16'h2300;
    SB_LUT4 i13783_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n64181), 
            .I3(n27), .O(n29644));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13783_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1853 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n60493));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1853.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1854 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n60492));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1854.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n60637));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n60491));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64079), .O(n64085));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n60490));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64085), .O(n64091));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'hfffe;
    SB_LUT4 i13784_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n64091), 
            .I3(n27), .O(n29645));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13784_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13377_3_lut_4_lut (.I0(n1747), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n29238));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13377_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_4_lut_adj_1860 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64205), .O(n64211));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1861 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n60489));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1861.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1862 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n60636));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1862.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64211), .O(n64217));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'hfffe;
    SB_LUT4 i13785_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n64217), 
            .I3(n27), .O(n29646));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13785_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4290_4_lut (.I0(n25156), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5725));
    defparam i4290_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5725), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n63449));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i13326_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n60771), .I3(GND_net), .O(n29187));   // verilog/coms.v(130[12] 305[6])
    defparam i13326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1864 (.I0(n63449), .I1(delay_counter[18]), .I2(n25153), 
            .I3(GND_net), .O(n63296));
    defparam i2_3_lut_adj_1864.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1865 (.I0(delay_counter[23]), .I1(n63296), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5777));
    defparam i2_4_lut_adj_1865.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n60635));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_LUT4 i4_4_lut_adj_1867 (.I0(n7_adj_5777), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n25158), .O(n62));
    defparam i4_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main_adj_5944[0]), .I1(o_Rx_DV_N_3488[24]), 
            .I2(n27), .I3(GND_net), .O(n14_adj_5837));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i23336_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(366[12:35])
    defparam i23336_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_adj_1868 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_5819));
    defparam i5_3_lut_adj_1868.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1869 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5818));
    defparam i6_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1870 (.I0(n29), .I1(o_Rx_DV_N_3488[12]), .I2(n23_adj_5852), 
            .I3(n5227), .O(n15_adj_5836));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i6_4_lut_adj_1870.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5818), .I1(delay_counter[2]), .I2(n14_adj_5819), 
            .I3(delay_counter[6]), .O(n25156));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1871 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5868));
    defparam i5_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1872 (.I0(delay_counter[28]), .I1(n12_adj_5868), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25158));
    defparam i6_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1873 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25153));
    defparam i2_3_lut_adj_1873.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_4_lut_adj_1874 (.I0(n15_adj_5836), .I1(n1), .I2(n14_adj_5837), 
            .I3(r_SM_Main_adj_5944[1]), .O(n72442));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i8_4_lut_adj_1874.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1875 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5858));
    defparam i1_2_lut_adj_1875.LUT_INIT = 16'heeee;
    SB_LUT4 i13375_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29236));   // verilog/coms.v(130[12] 305[6])
    defparam i13375_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1876 (.I0(delay_counter[9]), .I1(n4_adj_5858), 
            .I2(delay_counter[10]), .I3(n25156), .O(n63448));
    defparam i2_4_lut_adj_1876.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1877 (.I0(n63448), .I1(n25153), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n62711));
    defparam i2_4_lut_adj_1877.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5869));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1878 (.I0(delay_counter[22]), .I1(n62711), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5870));
    defparam i2_4_lut_adj_1878.LUT_INIT = 16'ha8a0;
    SB_LUT4 i23268_4_lut (.I0(n7_adj_5870), .I1(delay_counter[31]), .I2(n25158), 
            .I3(n8_adj_5869), .O(n1323));   // verilog/TinyFPGA_B.v(380[14:38])
    defparam i23268_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i589_2_lut (.I0(n1323), .I1(n39001), .I2(GND_net), .I3(GND_net), 
            .O(n2828));   // verilog/TinyFPGA_B.v(384[18] 386[12])
    defparam i589_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13791_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[1]), 
            .I2(n10_adj_5844), .I3(n25302), .O(n29652));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13791_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48130_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n65211));
    defparam i48130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13323_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n60771), .I3(GND_net), .O(n29184));   // verilog/coms.v(130[12] 305[6])
    defparam i13323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54722_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6910), .I2(n65211), 
            .I3(n25_adj_5820), .O(n17_adj_5727));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i54722_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n60634));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n60633));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1881 (.I0(state[0]), .I1(n23_adj_5867), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5857));
    defparam i1_2_lut_adj_1881.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut (.I0(n35689), .I1(n39530), .I2(state[1]), .I3(n4_adj_5857), 
            .O(n5_adj_5860));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i13793_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[2]), 
            .I2(n4_adj_5757), .I3(n25348), .O(n29654));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13793_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n60632));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1883 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n60631));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1883.LUT_INIT = 16'h2300;
    SB_LUT4 i13320_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n60771), .I3(GND_net), .O(n29181));   // verilog/coms.v(130[12] 305[6])
    defparam i13320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n60630));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 i13317_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n60771), .I3(GND_net), .O(n29178));   // verilog/coms.v(130[12] 305[6])
    defparam i13317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n60629));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 i13314_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n60771), .I3(GND_net), .O(n29175));   // verilog/coms.v(130[12] 305[6])
    defparam i13314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n60628));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n60488));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n60627));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n60626));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n60625));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_adj_1891 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n61213));
    defparam i1_2_lut_3_lut_adj_1891.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n60542));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n60487));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 i13797_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[3]), 
            .I2(n4_adj_5757), .I3(n25302), .O(n29658));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13797_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13798_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[4]), 
            .I2(n4_adj_5758), .I3(n25348), .O(n29659));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13798_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n60486));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_LUT4 i13799_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[5]), 
            .I2(n4_adj_5758), .I3(n25302), .O(n29660));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13799_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n60485));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n60484));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 i44471_4_lut_4_lut (.I0(hall3), .I1(hall2), .I2(hall1), .I3(commutation_state[2]), 
            .O(n61501));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i44471_4_lut_4_lut.LUT_INIT = 16'h8b0a;
    SB_LUT4 i13800_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[6]), 
            .I2(n39188), .I3(n25348), .O(n29661));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13800_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n60483));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1898 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n60482));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1898.LUT_INIT = 16'h2300;
    SB_LUT4 i13311_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n60771), .I3(GND_net), .O(n29172));   // verilog/coms.v(130[12] 305[6])
    defparam i13311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n60481));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1900 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n60480));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1900.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n60479));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i13802_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[7]), 
            .I2(n39188), .I3(n25302), .O(n29663));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13802_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n60478));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n60477));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n60624));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n60623));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 i14_4_lut (.I0(n68468), .I1(state_adj_5954[0]), .I2(n6714), 
            .I3(n39034), .O(n6_adj_5865));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14_4_lut.LUT_INIT = 16'h5cfc;
    SB_LUT4 i13807_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5921[0]), 
            .I2(n10_adj_5844), .I3(n25348), .O(n29668));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13807_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n60543));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i23223_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i23223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23222_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i23222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23343_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i23343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n31_adj_5854));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n60622));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n60621));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n60620));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n29020));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54832 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[2]), .O(n71939));
    defparam byte_transmit_counter_0__bdd_4_lut_54832.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n60619));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n60618));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n60617));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n60616));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n60615));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1917 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n60657));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1917.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n60656));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1919 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n60655));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1919.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n60654));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n60653));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n60652));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n60651));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 i13249_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n22465), .I3(GND_net), .O(n29110));   // verilog/coms.v(130[12] 305[6])
    defparam i13249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n60650));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 n71939_bdd_4_lut (.I0(n71939), .I1(\data_out_frame[19] [0]), 
            .I2(\data_out_frame[18] [0]), .I3(byte_transmit_counter[2]), 
            .O(n71942));
    defparam n71939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n60649));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n60648));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n60647));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n60614));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n60613));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n60612));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1931 (.I0(n4_adj_5759), .I1(r_SM_Main[1]), .I2(n6_adj_5866), 
            .I3(r_Bit_Index[0]), .O(n64115));
    defparam i1_4_lut_adj_1931.LUT_INIT = 16'hfffb;
    SB_LUT4 i51766_2_lut (.I0(n72092), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68433));
    defparam i51766_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n60611));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n60610));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n60609));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n60608));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 i13335_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n28102), .I3(GND_net), .O(n29196));   // verilog/coms.v(130[12] 305[6])
    defparam i13335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n60607));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n60606));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 i54530_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n39001), .I3(GND_net), .O(n27482));
    defparam i54530_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i51775_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n68344));
    defparam i51775_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n60605));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1939 (.I0(o_Rx_DV_N_3488[12]), .I1(n5224), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n64115), .O(n64121));
    defparam i1_4_lut_adj_1939.LUT_INIT = 16'hfffe;
    SB_LUT4 i23337_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n39001), .I3(GND_net), .O(n39100));
    defparam i23337_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n60604));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i53617_3_lut (.I0(n72056), .I1(n71942), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n70707));
    defparam i53617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1941 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5852), 
            .I3(n64121), .O(n64127));
    defparam i1_4_lut_adj_1941.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1942 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n60603));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1942.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n29002));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n60602));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n60601));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n60600));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n60599));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_LUT4 i13818_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n64127), 
            .I3(n27), .O(n29679));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13818_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13822_4_lut (.I0(CS_MISO_c), .I1(data_adj_5928[0]), .I2(n11_adj_5765), 
            .I3(state_7__N_4319), .O(n29683));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13822_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n60598));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n60597));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n60596));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n60595));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5744));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5754));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5752));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5747));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n60594));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n60593));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5746));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5745));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5735));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5736));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5732));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5733));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5740));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n60592));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5738));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5737));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5742));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52175_4_lut (.I0(n11_adj_5737), .I1(n9_adj_5738), .I2(n7_adj_5740), 
            .I3(n5_adj_5742), .O(n69265));
    defparam i52175_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5739), .I1(current_limit[9]), 
            .I2(n19_adj_5732), .I3(GND_net), .O(n16_adj_5734));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5743));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i53870_3_lut (.I0(n4_adj_5743), .I1(current_limit[5]), .I2(n11_adj_5737), 
            .I3(GND_net), .O(n70960));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53871_3_lut (.I0(n70960), .I1(current_limit[6]), .I2(n13_adj_5736), 
            .I3(GND_net), .O(n70961));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i53871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52169_4_lut (.I0(n17_adj_5733), .I1(n15_adj_5735), .I2(n13_adj_5736), 
            .I3(n69265), .O(n69259));
    defparam i52169_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54217_4_lut (.I0(n16_adj_5734), .I1(n6_adj_5741), .I2(n19_adj_5732), 
            .I3(n69251), .O(n71307));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54217_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52518_3_lut (.I0(n70961), .I1(current_limit[7]), .I2(n15_adj_5735), 
            .I3(GND_net), .O(n69608));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54422_4_lut (.I0(n69608), .I1(n71307), .I2(n19_adj_5732), 
            .I3(n69259), .O(n71512));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54422_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54423_3_lut (.I0(n71512), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n71513));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54423_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54331_3_lut (.I0(n71513), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5731));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i54331_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1955 (.I0(current_limit[13]), .I1(n24_adj_5731), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n63208));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1955.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n60591));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1957 (.I0(current_limit[13]), .I1(n24_adj_5731), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n63212));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1957.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n60590));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1959 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n63212), .I3(n63208), .O(n260));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i1_4_lut_adj_1959.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n60589));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5751));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n60588));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5750));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5749));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5708));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n60587));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n60586));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n60585));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n60584));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n60583));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37681_2_lut_3_lut_4_lut (.I0(n34395), .I1(Ki[0]), .I2(n341), 
            .I3(Ki[1]), .O(n20628));
    defparam i37681_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n68285), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53874_3_lut (.I0(n4), .I1(n305), .I2(n11), .I3(GND_net), 
            .O(n70964));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53875_3_lut (.I0(n70964), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n70965));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i53875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37683_2_lut_3_lut_4_lut (.I0(n34395), .I1(Ki[0]), .I2(n341), 
            .I3(Ki[1]), .O(n53436));
    defparam i37683_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8_adj_5729));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n60582));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7), .I3(GND_net), 
            .O(n6_adj_5730));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5729), .I1(n301), .I2(n19_adj_5708), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n60581));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 i52255_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n69345));
    defparam i52255_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37627_3_lut_4_lut (.I0(n34395), .I1(Ki[3]), .I2(n4_adj_5848), 
            .I3(n20719), .O(n6_adj_5847));
    defparam i37627_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n60580));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i52225_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n69345), 
            .O(n69315));
    defparam i52225_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54157_4_lut (.I0(n16), .I1(n6_adj_5730), .I2(n19_adj_5708), 
            .I3(n69299), .O(n71247));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54157_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n60579));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n60578));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_4_lut_adj_1972 (.I0(n34395), .I1(Ki[3]), .I2(n4_adj_5848), 
            .I3(n20719), .O(n20682));
    defparam i1_3_lut_4_lut_adj_1972.LUT_INIT = 16'h8778;
    SB_LUT4 i52510_3_lut (.I0(n70965), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n69600));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54392_4_lut (.I0(n69600), .I1(n71247), .I2(n19_adj_5708), 
            .I3(n69315), .O(n71482));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54392_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54393_3_lut (.I0(n71482), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n71483));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54393_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n60577));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 i54303_3_lut (.I0(n71483), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n71393));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i54303_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n60576));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 i47982_3_lut (.I0(duty[22]), .I1(duty[17]), .I2(n294), .I3(GND_net), 
            .O(n65059));
    defparam i47982_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i26_3_lut (.I0(n71393), .I1(n298), .I2(duty[12]), 
            .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47986_3_lut (.I0(duty[13]), .I1(duty[21]), .I2(n294), .I3(GND_net), 
            .O(n65063));
    defparam i47986_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i48112_4_lut (.I0(duty[15]), .I1(n65059), .I2(duty[20]), .I3(n294), 
            .O(n65193));
    defparam i48112_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i47978_3_lut (.I0(duty[14]), .I1(duty[18]), .I2(n294), .I3(GND_net), 
            .O(n65055));
    defparam i47978_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i10_4_lut (.I0(n294), .I1(n65193), .I2(n65063), .I3(n26), 
            .O(n22_adj_5845));
    defparam i10_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n60575));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i48110_4_lut (.I0(duty[19]), .I1(n65055), .I2(duty[16]), .I3(n294), 
            .O(n65191));
    defparam i48110_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1976 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n60574));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1976.LUT_INIT = 16'h2300;
    SB_LUT4 i52809_3_lut (.I0(n15_adj_5749), .I1(n13_adj_5750), .I2(n11_adj_5751), 
            .I3(GND_net), .O(n69899));
    defparam i52809_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i52685_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n69899), .O(n69775));
    defparam i52685_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n60573));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n60572));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 i51809_4_lut (.I0(n21_adj_5745), .I1(n19_adj_5746), .I2(n17_adj_5747), 
            .I3(n9_adj_5752), .O(n68899));
    defparam i51809_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52831_4_lut (.I0(n9_adj_5752), .I1(n7_adj_5754), .I2(current[2]), 
            .I3(duty[2]), .O(n69921));
    defparam i52831_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53403_4_lut (.I0(n15_adj_5749), .I1(n13_adj_5750), .I2(n11_adj_5751), 
            .I3(n69921), .O(n70493));
    defparam i53403_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53397_4_lut (.I0(n21_adj_5745), .I1(n19_adj_5746), .I2(n17_adj_5747), 
            .I3(n70493), .O(n70487));
    defparam i53397_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54078_4_lut (.I0(current[15]), .I1(n23_adj_5744), .I2(duty[12]), 
            .I3(n70487), .O(n71168));
    defparam i54078_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1979 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n60571));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1979.LUT_INIT = 16'h2300;
    SB_LUT4 i52777_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n71168), .O(n69867));
    defparam i52777_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5756));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i52643_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5749), .O(n69733));
    defparam i52643_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n60570));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n60569));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n60568));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n60567));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i53435_3_lut (.I0(n4_adj_5756), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n70525));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53435_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51700_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n69775), .O(n68790));
    defparam i51700_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_11_i35_rep_184_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n72606));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_184_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54143_3_lut (.I0(n30), .I1(n10), .I2(n69733), .I3(GND_net), 
            .O(n71233));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52536_4_lut (.I0(n70525), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n69626));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52536_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n60566));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i53433_3_lut (.I0(n6_adj_5755), .I1(duty[10]), .I2(n21_adj_5745), 
            .I3(GND_net), .O(n70523));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53434_3_lut (.I0(n70523), .I1(duty[11]), .I2(n23_adj_5744), 
            .I3(GND_net), .O(n70524));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53383_4_lut (.I0(current[15]), .I1(n23_adj_5744), .I2(duty[12]), 
            .I3(n68899), .O(n70473));
    defparam i53383_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5753), .I1(duty[9]), .I2(n19_adj_5746), 
            .I3(GND_net), .O(n16_adj_5748));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54827 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(byte_transmit_counter[1]), .O(n71903));
    defparam byte_transmit_counter_0__bdd_4_lut_54827.LUT_INIT = 16'he4aa;
    SB_LUT4 i13575_3_lut (.I0(\data_in_frame[16] [0]), .I1(rx_data[0]), 
            .I2(n28113), .I3(GND_net), .O(n29436));   // verilog/coms.v(130[12] 305[6])
    defparam i13575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13578_3_lut (.I0(\data_in_frame[16] [1]), .I1(rx_data[1]), 
            .I2(n28113), .I3(GND_net), .O(n29439));   // verilog/coms.v(130[12] 305[6])
    defparam i13578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52538_3_lut (.I0(n70524), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n69628));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52538_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53724_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n69867), .O(n70814));
    defparam i53724_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i54306_4_lut (.I0(n69626), .I1(n71233), .I2(n72606), .I3(n68790), 
            .O(n71396));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54306_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53672_3_lut (.I0(n69628), .I1(n16_adj_5748), .I2(n70473), 
            .I3(GND_net), .O(n70762));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i53672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i54460_4_lut (.I0(n70762), .I1(n71396), .I2(n72606), .I3(n70814), 
            .O(n71550));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54460_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54128_4_lut (.I0(n71550), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n71218));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i54128_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i2_4_lut_adj_1985 (.I0(n71218), .I1(current[15]), .I2(duty[21]), 
            .I3(duty[20]), .O(n6));
    defparam i2_4_lut_adj_1985.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n60565));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_LUT4 i13581_3_lut (.I0(\data_in_frame[16] [2]), .I1(rx_data[2]), 
            .I2(n28113), .I3(GND_net), .O(n29442));   // verilog/coms.v(130[12] 305[6])
    defparam i13581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1987 (.I0(duty[22]), .I1(duty[23]), .I2(n6), 
            .I3(n260), .O(n9940));
    defparam i7_4_lut_adj_1987.LUT_INIT = 16'h3332;
    SB_LUT4 i13584_3_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(n28113), .I3(GND_net), .O(n29445));   // verilog/coms.v(130[12] 305[6])
    defparam i13584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n60564));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n60563));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n60562));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n60561));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n60560));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i51670_2_lut (.I0(n72086), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68429));
    defparam i51670_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n60559));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i13587_3_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(n28113), .I3(GND_net), .O(n29448));   // verilog/coms.v(130[12] 305[6])
    defparam i13587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n60558));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n60557));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n60556));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n60555));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n60554));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 i13590_3_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(n28113), .I3(GND_net), .O(n29451));   // verilog/coms.v(130[12] 305[6])
    defparam i13590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n60553));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 n71903_bdd_4_lut (.I0(n71903), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(byte_transmit_counter[1]), 
            .O(n71906));
    defparam n71903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n60475));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n60552));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5728), .I3(n15_adj_5790), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_91[6]), 
            .I2(n15_adj_5766), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(285[5] 288[10])
    defparam mux_243_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13758_3_lut_4_lut (.I0(\data_in_frame[23] [2]), .I1(rx_data[2]), 
            .I2(n37938), .I3(n39467), .O(n29619));   // verilog/coms.v(130[12] 305[6])
    defparam i13758_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22199_4_lut (.I0(n112), .I1(n60), .I2(rx_data[6]), .I3(\data_in_frame[16] [6]), 
            .O(n37982));   // verilog/coms.v(94[13:20])
    defparam i22199_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i22200_3_lut (.I0(n37982), .I1(\data_in_frame[16] [6]), .I2(reset), 
            .I3(GND_net), .O(n29456));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n60551));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n60550));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n60549));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 i13755_3_lut_4_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(n37938), .I3(n39467), .O(n29616));   // verilog/coms.v(130[12] 305[6])
    defparam i13755_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_2005 (.I0(\FRAME_MATCHER.i [5]), .I1(n8), .I2(GND_net), 
            .I3(GND_net), .O(n110));
    defparam i1_2_lut_adj_2005.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2006 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n60548));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2006.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2007 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n60547));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2007.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n60546));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 i22184_4_lut (.I0(n112), .I1(n60), .I2(rx_data[7]), .I3(\data_in_frame[16] [7]), 
            .O(n37967));   // verilog/coms.v(94[13:20])
    defparam i22184_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n60545));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i13253_3_lut (.I0(current[0]), .I1(data_adj_5928[0]), .I2(n27489), 
            .I3(GND_net), .O(n29114));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22185_3_lut (.I0(n37967), .I1(\data_in_frame[16] [7]), .I2(reset), 
            .I3(GND_net), .O(n29459));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i22185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n60544));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2011 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n60541));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2011.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2012 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n60540));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2012.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n60539));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2014 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n60538));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2014.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2015 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n60537));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2015.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2016 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n60536));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2016.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2017 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n60535));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2017.LUT_INIT = 16'h2300;
    SB_LUT4 i13768_3_lut_4_lut (.I0(\data_in_frame[23] [5]), .I1(rx_data[5]), 
            .I2(n37938), .I3(n39467), .O(n29629));   // verilog/coms.v(130[12] 305[6])
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13771_3_lut_4_lut (.I0(\data_in_frame[23] [6]), .I1(rx_data[6]), 
            .I2(n37938), .I3(n39467), .O(n29632));   // verilog/coms.v(130[12] 305[6])
    defparam i13771_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13774_3_lut_4_lut (.I0(\data_in_frame[23] [7]), .I1(rx_data[7]), 
            .I2(n37938), .I3(n39467), .O(n29635));   // verilog/coms.v(130[12] 305[6])
    defparam i13774_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i13857_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n22465), .I3(GND_net), .O(n29718));   // verilog/coms.v(130[12] 305[6])
    defparam i13857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_2018 (.I0(hall3), .I1(hall2), .I2(commutation_state[1]), 
            .I3(hall1), .O(n60302));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i1_3_lut_4_lut_adj_2018.LUT_INIT = 16'hc454;
    SB_LUT4 i13858_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n22465), .I3(GND_net), .O(n29719));   // verilog/coms.v(130[12] 305[6])
    defparam i13858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13859_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n22465), .I3(GND_net), .O(n29720));   // verilog/coms.v(130[12] 305[6])
    defparam i13859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13860_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n22465), .I3(GND_net), .O(n29721));   // verilog/coms.v(130[12] 305[6])
    defparam i13860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13861_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n22465), .I3(GND_net), .O(n29722));   // verilog/coms.v(130[12] 305[6])
    defparam i13861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13862_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n22465), .I3(GND_net), .O(n29723));   // verilog/coms.v(130[12] 305[6])
    defparam i13862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13863_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n22465), .I3(GND_net), .O(n29724));   // verilog/coms.v(130[12] 305[6])
    defparam i13863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27507), .O(n56754));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i13864_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n22465), .I3(GND_net), .O(n29725));   // verilog/coms.v(130[12] 305[6])
    defparam i13864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5863));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 i13865_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n22465), .I3(GND_net), .O(n29726));   // verilog/coms.v(130[12] 305[6])
    defparam i13865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1323), .I3(n39001), .O(n24_adj_5726));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i13866_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21] [6]), 
            .I2(n22465), .I3(GND_net), .O(n29727));   // verilog/coms.v(130[12] 305[6])
    defparam i13866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13867_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n22465), .I3(GND_net), .O(n29728));   // verilog/coms.v(130[12] 305[6])
    defparam i13867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13868_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n22465), .I3(GND_net), .O(n29729));   // verilog/coms.v(130[12] 305[6])
    defparam i13868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13353_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n28102), .I3(GND_net), .O(n29214));   // verilog/coms.v(130[12] 305[6])
    defparam i13353_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13869_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n22465), .I3(GND_net), .O(n29730));   // verilog/coms.v(130[12] 305[6])
    defparam i13869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13350_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n28102), .I3(GND_net), .O(n29211));   // verilog/coms.v(130[12] 305[6])
    defparam i13350_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13870_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n22465), .I3(GND_net), .O(n29731));   // verilog/coms.v(130[12] 305[6])
    defparam i13870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13871_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n22465), .I3(GND_net), .O(n29732));   // verilog/coms.v(130[12] 305[6])
    defparam i13871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13347_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n28102), .I3(GND_net), .O(n29208));   // verilog/coms.v(130[12] 305[6])
    defparam i13347_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12967_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5856), 
            .I2(commutation_state_prev[0]), .I3(n38983), .O(n28828));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i12967_2_lut_4_lut.LUT_INIT = 16'h00de;
    SB_LUT4 i23220_2_lut (.I0(n22661), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n38983));
    defparam i23220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_2019 (.I0(commutation_state[0]), .I1(n4_adj_5856), 
            .I2(commutation_state_prev[0]), .I3(n38983), .O(n27664));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2019.LUT_INIT = 16'hffde;
    SB_LUT4 i1_2_lut_4_lut_adj_2020 (.I0(commutation_state[0]), .I1(n4_adj_5856), 
            .I2(commutation_state_prev[0]), .I3(dti_N_404), .O(n27417));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2020.LUT_INIT = 16'hdeff;
    SB_LUT4 i13872_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n22465), .I3(GND_net), .O(n29733));   // verilog/coms.v(130[12] 305[6])
    defparam i13872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13873_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n22465), .I3(GND_net), .O(n29734));   // verilog/coms.v(130[12] 305[6])
    defparam i13873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13628_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n28117), .I3(GND_net), .O(n29489));   // verilog/coms.v(130[12] 305[6])
    defparam i13628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13875_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n22465), .I3(GND_net), .O(n29736));   // verilog/coms.v(130[12] 305[6])
    defparam i13875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13631_3_lut (.I0(\data_in_frame[18] [1]), .I1(rx_data[1]), 
            .I2(n28117), .I3(GND_net), .O(n29492));   // verilog/coms.v(130[12] 305[6])
    defparam i13631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13634_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n28117), .I3(GND_net), .O(n29495));   // verilog/coms.v(130[12] 305[6])
    defparam i13634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13637_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n28117), .I3(GND_net), .O(n29498));   // verilog/coms.v(130[12] 305[6])
    defparam i13637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13877_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n22465), .I3(GND_net), .O(n29738));   // verilog/coms.v(130[12] 305[6])
    defparam i13877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13878_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n22465), .I3(GND_net), .O(n29739));   // verilog/coms.v(130[12] 305[6])
    defparam i13878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut_adj_2021 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n39001), .O(n59166));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_4_lut_4_lut_adj_2021.LUT_INIT = 16'hb1f1;
    SB_LUT4 i13258_3_lut (.I0(CS_c), .I1(state_adj_5930[0]), .I2(state_adj_5930[1]), 
            .I3(GND_net), .O(n29119));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13258_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i54737_4_lut (.I0(n15_adj_5764), .I1(clk_out), .I2(state_adj_5930[0]), 
            .I3(state_adj_5930[1]), .O(n9_adj_5864));   // verilog/tli4970.v(35[10] 68[6])
    defparam i54737_4_lut.LUT_INIT = 16'hc8fc;
    coms neopxl_color_23__I_0 (.GND_net(GND_net), .n59876(n59876), .VCC_net(VCC_net), 
         .\data_in_frame[23] ({\data_in_frame[23] }), .clk16MHz(clk16MHz), 
         .n2881(n2881), .\data_out_frame[18] ({\data_out_frame[18] }), .n60534(n60534), 
         .n60533(n60533), .n29193(n29193), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n60532(n60532), .setpoint({setpoint}), .reset(reset), .n29619(n29619), 
         .n60531(n60531), .n28930(n28930), .n29616(n29616), .n60530(n60530), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n60474(n60474), 
         .n60529(n60529), .n60528(n60528), .n60527(n60527), .n60526(n60526), 
         .n60525(n60525), .n60524(n60524), .n60523(n60523), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n60522(n60522), .rx_data({rx_data}), .n60476(n60476), .n60521(n60521), 
         .n60520(n60520), .n60519(n60519), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .n60646(n60646), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .n60645(n60645), .\data_out_frame[3][7] (\data_out_frame[3] [7]), 
         .n60644(n60644), .n29613(n29613), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .n60643(n60643), .\data_in_frame[1] ({\data_in_frame[1] [7], Open_4, 
         Open_5, \data_in_frame[1] [4], Open_6, Open_7, \data_in_frame[1] [1], 
         Open_8}), .n60642(n60642), .n60658(n60658), .n60641(n60641), 
         .n60518(n60518), .\data_in_frame[8][6] (\data_in_frame[8] [6]), 
         .n17(n17_adj_5789), .control_mode({Open_9, Open_10, Open_11, 
         Open_12, Open_13, Open_14, control_mode[1:0]}), .n22(n22_adj_5786), 
         .\data_in_frame[8][2] (\data_in_frame[8] [2]), .n60517(n60517), 
         .n60516(n60516), .\data_in_frame[20] ({\data_in_frame[20] }), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n60515(n60515), .n60514(n60514), .n60513(n60513), .n60512(n60512), 
         .n60511(n60511), .n60510(n60510), .n60509(n60509), .n60508(n60508), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .n60507(n60507), 
         .n60506(n60506), .n60505(n60505), .n60504(n60504), .n60503(n60503), 
         .n60502(n60502), .n60501(n60501), .n60500(n60500), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .n60499(n60499), .n60640(n60640), .n60639(n60639), .n60638(n60638), 
         .n60498(n60498), .n60497(n60497), .n60496(n60496), .n60495(n60495), 
         .n60494(n60494), .n60493(n60493), .n60492(n60492), .n60637(n60637), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n60491(n60491), 
         .n60490(n60490), .n25647(n25647), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .displacement({displacement}), .n60489(n60489), .\data_in_frame[8][3] (\data_in_frame[8] [3]), 
         .n25732(n25732), .\data_out_frame[5] ({\data_out_frame[5] }), .n60636(n60636), 
         .n60635(n60635), .n60634(n60634), .n60633(n60633), .n60632(n60632), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .n60631(n60631), .n60630(n60630), 
         .n29196(n29196), .n60629(n60629), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .n60628(n60628), .n60488(n60488), .n60627(n60627), .n60626(n60626), 
         .n60625(n60625), .n60542(n60542), .n60487(n60487), .n60486(n60486), 
         .n60485(n60485), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n60484(n60484), .n60483(n60483), .n60482(n60482), .n60481(n60481), 
         .n60480(n60480), .n60479(n60479), .control_update(control_update), 
         .n27465(n27465), .\data_out_frame[7] ({\data_out_frame[7] }), .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), 
         .n60478(n60478), .n60477(n60477), .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), 
         .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), 
         .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), 
         .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .n60624(n60624), .byte_transmit_counter({Open_15, 
         Open_16, Open_17, byte_transmit_counter[4:0]}), .n60623(n60623), 
         .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), .n161(n161), 
         .\data_in_frame[16] ({\data_in_frame[16] }), .\data_in_frame[18] ({\data_in_frame[18] }), 
         .\encoder0_position_scaled[23] (encoder0_position_scaled[23]), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n60543(n60543), .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), 
         .n28096(n28096), .n8(n8), .tx_active(tx_active), .n31(n31_adj_5854), 
         .n60622(n60622), .pwm_setpoint({pwm_setpoint}), .\pwm_counter[15] (pwm_counter[15]), 
         .n31_adj_10(n31), .\data_in_frame[10] ({\data_in_frame[10] [7:4], 
         Open_18, Open_19, Open_20, Open_21}), .n60621(n60621), .\pwm_counter[16] (pwm_counter[16]), 
         .n33(n33), .n29199(n29199), .n60620(n60620), .n29020(n29020), 
         .n60619(n60619), .\data_in_frame[8][7] (\data_in_frame[8] [7]), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .n60896(n60896), .\data_out_frame[8][6] (\data_out_frame[8] [6]), 
         .\control_mode[6] (control_mode[6]), .n48532(n48532), .\control_mode[2] (control_mode[2]), 
         .\control_mode[4] (control_mode[4]), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .n29520(n29520), .n29513(n29513), .n59920(n59920), .\encoder0_position_scaled[21] (encoder0_position_scaled[21]), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .\data_in_frame[1][2] (\data_in_frame[1] [2]), 
         .n59922(n59922), .n29205(n29205), .n29501(n29501), .n29498(n29498), 
         .n29495(n29495), .n29492(n29492), .n29489(n29489), .n29486(n29486), 
         .n29483(n29483), .n29480(n29480), .n29477(n29477), .n29208(n29208), 
         .n29473(n29473), .n60618(n60618), .n29211(n29211), .n29214(n29214), 
         .n29466(n29466), .n29463(n29463), .n29460(n29460), .n29459(n29459), 
         .n29456(n29456), .n60617(n60617), .n29451(n29451), .n29448(n29448), 
         .n68429(n68429), .n29445(n29445), .n29442(n29442), .n29439(n29439), 
         .n29436(n29436), .n60616(n60616), .\data_in_frame[14][6] (\data_in_frame[14] [6]), 
         .\data_out_frame[8][1] (\data_out_frame[8] [1]), .n60615(n60615), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .n60657(n60657), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n60656(n60656), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n60655(n60655), 
         .\data_out_frame[1][0] (\data_out_frame[1] [0]), .n60654(n60654), 
         .\data_out_frame[1][1] (\data_out_frame[1] [1]), .n60653(n60653), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .n60652(n60652), 
         .\data_out_frame[1][5] (\data_out_frame[1] [5]), .n60651(n60651), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .n60650(n60650), 
         .\data_out_frame[1][7] (\data_out_frame[1] [7]), .n60649(n60649), 
         .\data_out_frame[3][1] (\data_out_frame[3] [1]), .n60648(n60648), 
         .\data_out_frame[3][3] (\data_out_frame[3] [3]), .n60647(n60647), 
         .\data_out_frame[8][2] (\data_out_frame[8] [2]), .n60614(n60614), 
         .\data_out_frame[8][3] (\data_out_frame[8] [3]), .n60613(n60613), 
         .\data_out_frame[8][4] (\data_out_frame[8] [4]), .n60612(n60612), 
         .\data_out_frame[8][5] (\data_out_frame[8] [5]), .n60611(n60611), 
         .n60610(n60610), .\data_out_frame[8][7] (\data_out_frame[8] [7]), 
         .n60609(n60609), .\data_out_frame[9] ({\data_out_frame[9] }), .n60608(n60608), 
         .n60607(n60607), .n60606(n60606), .n60605(n60605), .n60604(n60604), 
         .n60603(n60603), .n29002(n29002), .n60602(n60602), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n60601(n60601), .n60600(n60600), .n60599(n60599), .n60598(n60598), 
         .n60597(n60597), .n60596(n60596), .n60595(n60595), .n60594(n60594), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n60593(n60593), 
         .n60592(n60592), .n60591(n60591), .n60590(n60590), .n60589(n60589), 
         .n60588(n60588), .n60587(n60587), .n60586(n60586), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n60585(n60585), .n60584(n60584), .n60583(n60583), .n60582(n60582), 
         .n60581(n60581), .n60580(n60580), .n60579(n60579), .n60578(n60578), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n60577(n60577), 
         .n60576(n60576), .n60575(n60575), .n60574(n60574), .n60573(n60573), 
         .n60572(n60572), .n60571(n60571), .n60570(n60570), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n60569(n60569), .n60568(n60568), .n60567(n60567), .n60566(n60566), 
         .n60565(n60565), .n60564(n60564), .n60563(n60563), .n60562(n60562), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .n60561(n60561), 
         .n60560(n60560), .n60559(n60559), .n60558(n60558), .n60557(n60557), 
         .n60556(n60556), .n60555(n60555), .n60554(n60554), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n60553(n60553), .n60475(n60475), .n60552(n60552), .n60551(n60551), 
         .n60550(n60550), .n60549(n60549), .n60548(n60548), .n60547(n60547), 
         .n60546(n60546), .n60545(n60545), .n29236(n29236), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n60544(n60544), .n60541(n60541), .n60540(n60540), .n60539(n60539), 
         .LED_c(LED_c), .n8_adj_11(n8_adj_5810), .DE_c(DE_c), .\data_in_frame[1][6] (\data_in_frame[1] [6]), 
         .n39467(n39467), .n3483(n3483), .n37935(n37935), .n60700(n60700), 
         .n60538(n60538), .n56640(n56640), .n72152(n72152), .n60537(n60537), 
         .n59930(n59930), .deadband({deadband}), .IntegralLimit({IntegralLimit}), 
         .\Kp[0] (Kp[0]), .\Ki[0] (Ki[0]), .PWMLimit({PWMLimit}), .n29629(n29629), 
         .n29632(n29632), .n29635(n29635), .n29948(n29948), .n29945(n29945), 
         .n29942(n29942), .n29939(n29939), .n29936(n29936), .n29933(n29933), 
         .n29930(n29930), .n29927(n29927), .n29127(n29127), .n29130(n29130), 
         .n29133(n29133), .\data_in_frame[8][4] (\data_in_frame[8] [4]), 
         .n56696(n56696), .n29136(n29136), .\data_in_frame[8][5] (\data_in_frame[8] [5]), 
         .n29139(n29139), .n29142(n29142), .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), 
         .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
         .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
         .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .n60536(n60536), 
         .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), 
         .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
         .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
         .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
         .\Ki[15] (Ki[15]), .neopxl_color({neopxl_color}), .n60535(n60535), 
         .n29739(n29739), .n29738(n29738), .n29736(n29736), .n29734(n29734), 
         .n29733(n29733), .\control_mode[7] (control_mode[7]), .n29732(n29732), 
         .current_limit({current_limit}), .n29731(n29731), .n29730(n29730), 
         .n29729(n29729), .n29728(n29728), .n29727(n29727), .n29726(n29726), 
         .n29725(n29725), .n29724(n29724), .n29723(n29723), .n29722(n29722), 
         .n29721(n29721), .n29720(n29720), .n29719(n29719), .n29718(n29718), 
         .n29110(n29110), .n29172(n29172), .\data_in_frame[10][1] (\data_in_frame[10] [1]), 
         .n29175(n29175), .\data_in_frame[10][2] (\data_in_frame[10] [2]), 
         .n29178(n29178), .\data_in_frame[10][3] (\data_in_frame[10] [3]), 
         .n29181(n29181), .n29184(n29184), .n29187(n29187), .n29190(n29190), 
         .n39431(n39431), .n110(n110), .n112(n112), .n37941(n37941), 
         .n68422(n68422), .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), 
         .rx_data_ready(rx_data_ready), .n24820(n24820), .n34686(n34686), 
         .n34584(n34584), .n62686(n62686), .encoder1_position_scaled({encoder1_position_scaled}), 
         .n56501(n56501), .n56624(n56624), .n56565(n56565), .n25994(n25994), 
         .n55945(n55945), .n61288(n61288), .n26215(n26215), .n60951(n60951), 
         .n55578(n55578), .n61213(n61213), .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), 
         .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), 
         .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), 
         .\encoder0_position_scaled[2] (encoder0_position_scaled[2]), .n61461(n61461), 
         .n26311(n26311), .n56545(n56545), .n31_adj_12(n31_adj_5842), 
         .n25712(n25712), .n61442(n61442), .\encoder0_position_scaled[1] (encoder0_position_scaled[1]), 
         .n61245(n61245), .n22465(n22465), .n28(n28), .n6(n6_adj_5859), 
         .n28102(n28102), .n60771(n60771), .n60766(n60766), .n8_adj_13(n8_adj_5849), 
         .n115(n115), .ID({ID}), .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), 
         .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), 
         .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), .n72092(n72092), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .n72086(n72086), 
         .n72122(n72122), .n71906(n71906), .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), 
         .\current[7] (current[7]), .\current[6] (current[6]), .\current[5] (current[5]), 
         .\current[4] (current[4]), .\current[3] (current[3]), .\current[2] (current[2]), 
         .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), .\current[1] (current[1]), 
         .\current[0] (current[0]), .\current[15] (current[15]), .\current[11] (current[11]), 
         .\current[10] (current[10]), .\current[9] (current[9]), .\current[8] (current[8]), 
         .n61134(n61134), .n72026(n72026), .n15(n15_adj_5728), .n7(n7_adj_5840), 
         .n31_adj_14(n31_adj_5816), .n15_adj_15(n15_adj_5790), .n15_adj_16(n15_adj_5766), 
         .r_SM_Main({r_SM_Main_adj_5944}), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
         .n1(n1), .tx_o(tx_o), .\tx_data[0] (tx_data[0]), .n5227(n5227), 
         .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
         .n29(n29), .n23(n23_adj_5852), .n62322(n62322), .n27(n27), 
         .\r_Bit_Index[0] (r_Bit_Index_adj_5946[0]), .n60413(n60413), .n63831(n63831), 
         .r_Clock_Count({r_Clock_Count_adj_5945}), .n27514(n27514), .n29671(n29671), 
         .n61481(n61481), .n29123(n29123), .n72442(n72442), .n63819(n63819), 
         .n6_adj_17(n6_adj_5846), .tx_enable(tx_enable), .baudrate({baudrate}), 
         .r_Rx_Data(r_Rx_Data), .r_SM_Main_adj_31({r_SM_Main}), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .n5224(n5224), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .RX_N_2(RX_N_2), 
         .n25296(n25296), .r_Clock_Count_adj_32({r_Clock_Count}), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), 
         .\r_Bit_Index[0]_adj_29 (r_Bit_Index[0]), .n60415(n60415), .n63843(n63843), 
         .n27507(n27507), .n27511(n27511), .n29674(n29674), .n56754(n56754), 
         .n29679(n29679), .n29646(n29646), .n29645(n29645), .n29644(n29644), 
         .n29642(n29642), .n29641(n29641), .n29640(n29640), .n29639(n29639), 
         .n61483(n61483), .n6_adj_30(n6_adj_5866), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), 
         .n64131(n64131), .n64079(n64079), .n64167(n64167), .n64205(n64205), 
         .n64169(n64169), .n64151(n64151), .n64133(n64133), .n64097(n64097), 
         .n4(n4_adj_5759), .n63821(n63821)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i5248_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5248_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i5246_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i5246_3_lut_4_lut.LUT_INIT = 16'h21cc;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1792(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .\encoder1_position[31] (encoder1_position[31]), 
            .GND_net(GND_net), .\encoder1_position[30] (encoder1_position[30]), 
            .\encoder1_position[29] (encoder1_position[29]), .\encoder1_position[28] (encoder1_position[28]), 
            .\encoder1_position[27] (encoder1_position[27]), .\encoder1_position[26] (encoder1_position[26]), 
            .\encoder1_position[25] (encoder1_position[25]), .\encoder1_position[24] (encoder1_position[24]), 
            .\encoder1_position[23] (encoder1_position[23]), .\encoder1_position[22] (encoder1_position[22]), 
            .\encoder1_position[21] (encoder1_position[21]), .\encoder1_position[20] (encoder1_position[20]), 
            .\encoder1_position[19] (encoder1_position[19]), .\encoder1_position[18] (encoder1_position[18]), 
            .\encoder1_position[17] (encoder1_position[17]), .\encoder1_position[16] (encoder1_position[16]), 
            .\encoder1_position[15] (encoder1_position[15]), .\encoder1_position[14] (encoder1_position[14]), 
            .\encoder1_position[13] (encoder1_position[13]), .\encoder1_position[12] (encoder1_position[12]), 
            .\encoder1_position[11] (encoder1_position[11]), .\encoder1_position[10] (encoder1_position[10]), 
            .\encoder1_position[9] (encoder1_position[9]), .\encoder1_position[8] (encoder1_position[8]), 
            .\encoder1_position[7] (encoder1_position[7]), .\encoder1_position[6] (encoder1_position[6]), 
            .\encoder1_position[5] (encoder1_position[5]), .\encoder1_position[4] (encoder1_position[4]), 
            .\encoder1_position[3] (encoder1_position[3]), .\encoder1_position[2] (encoder1_position[2]), 
            .n1829(n1829), .n1831(n1831), .VCC_net(VCC_net), .b_prev(b_prev_adj_5770), 
            .\a_new[1] (a_new_adj_5908[1]), .\b_new[1] (b_new_adj_5909[1]), 
            .n29239(n29239), .a_prev(a_prev_adj_5769), .position_31__N_3836(position_31__N_3836_adj_5772), 
            .n29125(n29125), .n29124(n29124), .n1797(n1797), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5771)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i642_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2881));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i642_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_2022 (.I0(n94), .I1(n115), .I2(n37941), 
            .I3(GND_net), .O(n28117));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_adj_2022.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_2023 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n94));
    defparam i1_2_lut_adj_2023.LUT_INIT = 16'h2222;
    SB_LUT4 i117_2_lut (.I0(reset), .I1(n39431), .I2(GND_net), .I3(GND_net), 
            .O(n115));
    defparam i117_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i10_2_lut_adj_2024 (.I0(PWMLimit[18]), .I1(setpoint[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i10_2_lut_adj_2024.LUT_INIT = 16'h6666;
    TLI4970 tli (.\data[15] (data_adj_5928[15]), .\state[1] (state_adj_5930[1]), 
            .\state[0] (state_adj_5930[0]), .n27489(n27489), .GND_net(GND_net), 
            .\data[12] (data_adj_5928[12]), .clk16MHz(clk16MHz), .n6(n6_adj_5762), 
            .n5(n5_adj_5763), .n5_adj_8(n5_adj_5791), .n6_adj_9(n6_adj_5761), 
            .n39133(n39133), .n39146(n39146), .\current[15] (current[15]), 
            .n29320(n29320), .\current[1] (current[1]), .n29319(n29319), 
            .\current[2] (current[2]), .n29318(n29318), .\current[3] (current[3]), 
            .n29317(n29317), .\current[4] (current[4]), .n29316(n29316), 
            .\current[5] (current[5]), .n29315(n29315), .\current[6] (current[6]), 
            .n29314(n29314), .\current[7] (current[7]), .n29313(n29313), 
            .\current[8] (current[8]), .n29312(n29312), .\current[9] (current[9]), 
            .n29311(n29311), .\current[10] (current[10]), .n29310(n29310), 
            .\current[11] (current[11]), .n15(n15_adj_5764), .n11(n11_adj_5765), 
            .n29880(n29880), .n29879(n29879), .n29878(n29878), .\data[11] (data_adj_5928[11]), 
            .n29877(n29877), .\data[10] (data_adj_5928[10]), .n29875(n29875), 
            .\data[9] (data_adj_5928[9]), .n29874(n29874), .\data[8] (data_adj_5928[8]), 
            .n29872(n29872), .\data[7] (data_adj_5928[7]), .n29871(n29871), 
            .\data[6] (data_adj_5928[6]), .n29869(n29869), .\data[5] (data_adj_5928[5]), 
            .n29868(n29868), .\data[4] (data_adj_5928[4]), .n29866(n29866), 
            .\data[3] (data_adj_5928[3]), .n29865(n29865), .\data[2] (data_adj_5928[2]), 
            .n29840(n29840), .\data[1] (data_adj_5928[1]), .n9(n9_adj_5864), 
            .clk_out(clk_out), .n29119(n29119), .CS_c(CS_c), .n29114(n29114), 
            .\current[0] (current[0]), .n29683(n29683), .\data[0] (data_adj_5928[0]), 
            .VCC_net(VCC_net), .n25298(n25298), .n25289(n25289), .state_7__N_4319(state_7__N_4319), 
            .CS_CLK_c(CS_CLK_c), .n25328(n25328), .n25345(n25345), .n25316(n25316)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(405[11] 411[4])
    SB_LUT4 i1_2_lut_3_lut_adj_2025 (.I0(n94), .I1(n115), .I2(n110), .I3(GND_net), 
            .O(n28113));   // verilog/TinyFPGA_B.v(359[10] 389[6])
    defparam i1_2_lut_3_lut_adj_2025.LUT_INIT = 16'h0202;
    SB_LUT4 i18760_3_lut (.I0(n8_adj_5812), .I1(PWMLimit[4]), .I2(setpoint[4]), 
            .I3(GND_net), .O(n10_adj_5813));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i18760_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i18721_3_lut (.I0(n10_adj_5813), .I1(PWMLimit[5]), .I2(setpoint[5]), 
            .I3(GND_net), .O(n12_adj_5814));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i18721_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_adj_2026 (.I0(n37938), .I1(n39467), .I2(GND_net), 
            .I3(GND_net), .O(n28127));
    defparam i1_2_lut_adj_2026.LUT_INIT = 16'h8888;
    SB_LUT4 i18967_3_lut (.I0(n20_adj_5815), .I1(PWMLimit[10]), .I2(setpoint[10]), 
            .I3(GND_net), .O(n34791));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i18967_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i11_4_lut_adj_2027 (.I0(\data_in_frame[23] [3]), .I1(n60700), 
            .I2(n28127), .I3(rx_data[3]), .O(n59876));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_2027.LUT_INIT = 16'hca0a;
    EEPROM eeprom (.GND_net(GND_net), .enable_slow_N_4213(enable_slow_N_4213), 
           .clk16MHz(clk16MHz), .\state_7__N_4110[0] (state_7__N_4110[0]), 
           .ID({ID}), .baudrate({baudrate}), .n29328(n29328), .n29327(n29327), 
           .n29326(n29326), .n29325(n29325), .n29324(n29324), .n29323(n29323), 
           .n29322(n29322), .n29321(n29321), .data_ready(data_ready), 
           .\state_7__N_3918[0] (state_7__N_3918[0]), .n63193(n63193), .data({data_adj_5921}), 
           .\state[0] (state_adj_5954[0]), .\state_7__N_4126[3] (state_7__N_4126[3]), 
           .scl_enable(scl_enable), .scl(scl), .n6714(n6714), .sda_enable(sda_enable), 
           .n29668(n29668), .n6(n6_adj_5865), .VCC_net(VCC_net), .n29663(n29663), 
           .n29661(n29661), .n29660(n29660), .n29659(n29659), .n29658(n29658), 
           .n29654(n29654), .n29652(n29652), .sda_out(sda_out), .n39034(n39034), 
           .n10(n10_adj_5760), .n25302(n25302), .n25348(n25348), .n4(n4_adj_5757), 
           .n4_adj_6(n4_adj_5758), .n39188(n39188), .n10_adj_7(n10_adj_5844)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(391[10] 403[6])
    motorControl control (.setpoint({setpoint}), .GND_net(GND_net), .\Kp[1] (Kp[1]), 
            .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Ki[4] (Ki[4]), .n358(n358), 
            .PWMLimit({PWMLimit}), .\motor_state[9] (motor_state[9]), .\Kp[3] (Kp[3]), 
            .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .duty({duty}), .n39420(n39420), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .n284(n284), 
            .IntegralLimit({IntegralLimit}), .n258(n258), .n359(n359), 
            .\Ki[0] (Ki[0]), .control_update(control_update), .n22(n22_adj_5786), 
            .\Ki[3] (Ki[3]), .n348(n348), .n337(n337), .n338(n338), 
            .n339(n339), .n341(n341), .n342(n342), .n343(n343), .n344(n344), 
            .n345(n345), .clk16MHz(clk16MHz), .reset(reset), .n349(n349), 
            .n350(n350), .n351(n351), .n352(n352), .n353(n353), .n354(n354), 
            .n355(n355), .n356(n356), .n357(n357), .\control_mode[7] (control_mode[7]), 
            .n17(n17_adj_5789), .n48532(n48532), .\control_mode[1] (control_mode[1]), 
            .\control_mode[0] (control_mode[0]), .\motor_state[8] (motor_state[8]), 
            .n238(n238), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .\motor_state[7] (motor_state[7]), .n336(n336), .\motor_state[6] (motor_state[6]), 
            .\motor_state[5] (motor_state[5]), .\Ki[5] (Ki[5]), .\motor_state[4] (motor_state[4]), 
            .\Ki[6] (Ki[6]), .n290(n290), .n39(n39_adj_5817), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .deadband({deadband}), 
            .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .n29864(n29864), .n29863(n29863), 
            .n29862(n29862), .n29861(n29861), .n29860(n29860), .n29859(n29859), 
            .n29858(n29858), .n29857(n29857), .n29856(n29856), .n29855(n29855), 
            .n29854(n29854), .n29853(n29853), .n29852(n29852), .n29851(n29851), 
            .n29850(n29850), .n29849(n29849), .n29848(n29848), .n29847(n29847), 
            .n29846(n29846), .n29845(n29845), .n29844(n29844), .n29843(n29843), 
            .n29839(n29839), .n29097(n29097), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
            .\Ki[15] (Ki[15]), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), .n346(n346), 
            .n347(n347), .n34584(n34584), .n34686(n34686), .VCC_net(VCC_net), 
            .\motor_state[3] (motor_state[3]), .\motor_state[2] (motor_state[2]), 
            .\motor_state[1] (motor_state[1]), .\Kp[13] (Kp[13]), .n17_adj_1(n17_adj_5853), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .n3(n3_adj_5841), .\motor_state[10] (motor_state[10]), 
            .\Kp[14] (Kp[14]), .n20628(n20628), .n20682(n20682), .n20719(n20719), 
            .n34395(n34395), .n6(n6_adj_5847), .\Kp[15] (Kp[15]), .\encoder1_position_scaled[0] (encoder1_position_scaled[0]), 
            .n15(n15_adj_5766), .n68243(n68243), .n15_adj_2(n15_adj_5728), 
            .n53436(n53436), .n131(n131), .n204(n204), .n4(n4_adj_5848), 
            .n4_adj_3(n4_adj_5811), .n8(n8_adj_5812), .n12(n12_adj_5814), 
            .n20(n20_adj_5815), .n31(n31_adj_5816), .n37(n37), .n34791(n34791)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 303[4])
    pwm PWM (.GND_net(GND_net), .\pwm_counter[16] (pwm_counter[16]), .\pwm_counter[19] (pwm_counter[19]), 
        .\pwm_counter[15] (pwm_counter[15]), .\pwm_counter[22] (pwm_counter[22]), 
        .\pwm_counter[21] (pwm_counter[21]), .\pwm_counter[20] (pwm_counter[20]), 
        .n2881(n2881), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .pwm_setpoint({pwm_setpoint}), 
        .n31(n31), .n33(n33), .n45(n45), .n43(n43), .VCC_net(VCC_net), 
        .n39(n39), .n41(n41), .reset(reset), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
        .\rx_data[7] (rx_data[7]), .n60771(n60771), .n29190(n29190), .\data_in_frame[10][6] (\data_in_frame[10] [6]), 
        .n25647(n25647), .n25732(n25732), .n60896(n60896)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, GND_net, state, 
            timer, VCC_net, n29377, bit_ctr, n5, n29347, t0, n29346, 
            n29345, n27645, n29344, n29343, n29342, n29341, n29340, 
            n29339, n29338, n35689, \bit_ctr[0] , NEOPXL_c, n29126, 
            neopxl_color, LED_c, n39530, n3172, n23) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    input GND_net;
    output [1:0]state;
    output [10:0]timer;
    input VCC_net;
    input n29377;
    output [4:0]bit_ctr;
    input n5;
    input n29347;
    output [10:0]t0;
    input n29346;
    input n29345;
    output n27645;
    input n29344;
    input n29343;
    input n29342;
    input n29341;
    input n29340;
    input n29339;
    input n29338;
    output n35689;
    output \bit_ctr[0] ;
    output NEOPXL_c;
    input n29126;
    input [23:0]neopxl_color;
    input LED_c;
    output n39530;
    output n3172;
    output n23;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n63032, \neo_pixel_transmitter.done , 
        start_N_507, n7, start, n25322, n50, n61673, n6, n63, 
        n4, n65195, n56, n66, n68282, n39054, n68281, n59, n1;
    wire [10:0]n49;
    
    wire n54460, n54459, n54458, n61, n61581, n44, n12, n54457, 
        n54456, n54455, n54454, n54453, n54452, n54451;
    wire [5:0]color_bit_N_502;
    
    wire n65635, n65636, n72017, n65459, n65458, n72020;
    wire [31:0]n149;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    
    wire n29064, n63103, n68474, n62802, n57_adj_5701, n43, n32, 
        one_wire_N_499, n6_adj_5702, n71852, n72116, n70583, n20767, 
        n27639, n28538;
    wire [1:0]state_1__N_451;
    
    wire n28537, n68432, n61487, n70904, n55684, n65371, n65372, 
        n65375, n65374, n71840;
    wire [10:0]n13;
    
    wire n53860, n53859, n53858, n53857, n53856, n53855, n53854, 
        n53853, n53852, n53851, n71849, n39155, n14, n72113, n7200, 
        n39007, n68464, n41, n71915, n71918;
    
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n63032), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i3_4_lut (.I0(t1[3]), .I1(t1[1]), .I2(t1[4]), .I3(t1[0]), 
            .O(n25322));   // verilog/neopixel.v(60[15:45])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(t1[4]), .I1(t1[0]), .I2(t1[2]), .I3(n50), 
            .O(n61673));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(n25322), .I1(t1[10]), .I2(t1[8]), .I3(n6), 
            .O(n63));
    defparam i4_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i48114_3_lut_4_lut (.I0(t1[4]), .I1(t1[0]), .I2(t1[10]), .I3(n4), 
            .O(n65195));
    defparam i48114_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(t1[2]), .I1(t1[4]), .I2(GND_net), .I3(GND_net), 
            .O(n56));   // verilog/neopixel.v(13[8] 16[4])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i83_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(n63), .I2(GND_net), 
            .I3(GND_net), .O(n66));
    defparam i83_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i51866_3_lut (.I0(n25322), .I1(n50), .I2(t1[2]), .I3(GND_net), 
            .O(n68282));   // verilog/neopixel.v(19[11:16])
    defparam i51866_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i52504_4_lut (.I0(n56), .I1(n50), .I2(n39054), .I3(t1[0]), 
            .O(n68281));   // verilog/neopixel.v(19[11:16])
    defparam i52504_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n68281), .I2(n68282), 
            .I3(state[0]), .O(n59));   // verilog/neopixel.v(19[11:16])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i15_4_lut (.I0(n59), .I1(n1), .I2(state[1]), .I3(start), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i54666_2_lut (.I0(state[1]), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i54666_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 timer_2039_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n54460), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2039_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n54459), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_11 (.CI(n54459), .I0(GND_net), .I1(timer[9]), 
            .CO(n54460));
    SB_LUT4 timer_2039_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n54458), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1754 (.I0(t1[5]), .I1(t1[6]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1754.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1755 (.I0(t1[9]), .I1(t1[7]), .I2(GND_net), .I3(GND_net), 
            .O(n61));
    defparam i1_2_lut_adj_1755.LUT_INIT = 16'heeee;
    SB_LUT4 i23291_2_lut (.I0(t1[1]), .I1(t1[3]), .I2(GND_net), .I3(GND_net), 
            .O(n39054));
    defparam i23291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i44543_2_lut (.I0(t1[3]), .I1(t1[1]), .I2(GND_net), .I3(GND_net), 
            .O(n61581));
    defparam i44543_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(t1[2]), .I1(t1[8]), .I2(n44), .I3(n61), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i2_4_lut (.I0(state[1]), .I1(n65195), .I2(start), .I3(n12), 
            .O(n63032));
    defparam i2_4_lut.LUT_INIT = 16'hfbfa;
    SB_CARRY timer_2039_add_4_10 (.CI(n54458), .I0(GND_net), .I1(timer[8]), 
            .CO(n54459));
    SB_LUT4 timer_2039_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n54457), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19908_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(19[11:16])
    defparam i19908_3_lut.LUT_INIT = 16'hc1c1;
    SB_CARRY timer_2039_add_4_9 (.CI(n54457), .I0(GND_net), .I1(timer[7]), 
            .CO(n54458));
    SB_LUT4 timer_2039_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n54456), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_8 (.CI(n54456), .I0(GND_net), .I1(timer[6]), 
            .CO(n54457));
    SB_LUT4 timer_2039_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n54455), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_7 (.CI(n54455), .I0(GND_net), .I1(timer[5]), 
            .CO(n54456));
    SB_LUT4 timer_2039_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n54454), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_6 (.CI(n54454), .I0(GND_net), .I1(timer[4]), 
            .CO(n54455));
    SB_LUT4 timer_2039_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n54453), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_5 (.CI(n54453), .I0(GND_net), .I1(timer[3]), 
            .CO(n54454));
    SB_LUT4 timer_2039_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n54452), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_4 (.CI(n54452), .I0(GND_net), .I1(timer[2]), 
            .CO(n54453));
    SB_LUT4 timer_2039_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n54451), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_3 (.CI(n54451), .I0(GND_net), .I1(timer[1]), 
            .CO(n54452));
    SB_LUT4 timer_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n54451));
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(color_bit_N_502[1]), .I1(n65635), 
            .I2(n65636), .I3(color_bit_N_502[2]), .O(n72017));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n72017_bdd_4_lut (.I0(n72017), .I1(n65459), .I2(n65458), .I3(color_bit_N_502[2]), 
            .O(n72020));
    defparam n72017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(VCC_net), .D(n29377));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n5));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n29347));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n29346));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n4), .I1(n61), .I2(t1[2]), .I3(GND_net), 
            .O(n6));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF timer_2039__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n29345));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n27645), 
            .D(n149[2]), .R(n29064));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr_c[3]), .C(clk16MHz), .E(n27645), 
            .D(n149[3]), .R(n29064));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr_c[4]), .C(clk16MHz), .E(n27645), 
            .D(n149[4]), .R(n29064));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n29344));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n29343));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n29342));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n29341));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n29340));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n29339));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n29338));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1756 (.I0(n4), .I1(n61), .I2(t1[8]), .I3(t1[10]), 
            .O(n50));
    defparam i2_3_lut_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1757 (.I0(state[1]), .I1(state[0]), .I2(n63), 
            .I3(\neo_pixel_transmitter.done ), .O(n63103));   // verilog/neopixel.v(34[12] 113[6])
    defparam i2_4_lut_adj_1757.LUT_INIT = 16'h0020;
    SB_LUT4 i52341_3_lut (.I0(n63), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n68474));
    defparam i52341_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_4_lut_adj_1758 (.I0(n61581), .I1(n61673), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n62802));
    defparam i2_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 i61_4_lut (.I0(n62802), .I1(n68474), .I2(state[1]), .I3(start), 
            .O(n57_adj_5701));
    defparam i61_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i54741_3_lut (.I0(n43), .I1(n57_adj_5701), .I2(n61673), .I3(GND_net), 
            .O(n32));
    defparam i54741_3_lut.LUT_INIT = 16'h3131;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));   // verilog/neopixel.v(34[12] 113[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(n35689), .I1(n66), .I2(state[1]), .I3(state[0]), 
            .O(n6_adj_5702));
    defparam i14_4_lut.LUT_INIT = 16'hfa3a;
    SB_LUT4 i53493_3_lut (.I0(n71852), .I1(n72116), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n70583));
    defparam i53493_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR bit_ctr_i0 (.Q(\bit_ctr[0] ), .C(clk16MHz), .E(n27639), 
            .D(n20767), .R(n28538));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n6_adj_5702), .D(state_1__N_451[0]), 
            .S(n28537));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i23240_4_lut (.I0(n68432), .I1(n61487), .I2(n70904), .I3(n55684), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i23240_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n32), .D(one_wire_N_499), 
            .R(n63103));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n29126));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2039__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 i48281_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n65371));
    defparam i48281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48282_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n65372));
    defparam i48282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48285_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n65375));
    defparam i48285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48284_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n65374));
    defparam i48284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71837_bdd_4_lut_4_lut_4_lut_4_lut (.I0(t1[3]), .I1(t1[1]), 
            .I2(state[0]), .I3(\neo_pixel_transmitter.done ), .O(n71840));
    defparam n71837_bdd_4_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h1881;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n53860), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n13[9]), 
            .I3(n53859), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n53859), .I0(timer[9]), .I1(n13[9]), 
            .CO(n53860));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n53858), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n53858), .I0(timer[8]), .I1(n13[8]), 
            .CO(n53859));
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n53857), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n53857), .I0(timer[7]), .I1(n13[7]), 
            .CO(n53858));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n13[6]), 
            .I3(n53856), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n53856), .I0(timer[6]), .I1(n13[6]), 
            .CO(n53857));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n13[5]), 
            .I3(n53855), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n53855), .I0(timer[5]), .I1(n13[5]), 
            .CO(n53856));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n53854), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n53854), .I0(timer[4]), .I1(n13[4]), 
            .CO(n53855));
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n53853), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n53853), .I0(timer[3]), .I1(n13[3]), 
            .CO(n53854));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n53852), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n53852), .I0(timer[2]), .I1(n13[2]), 
            .CO(n53853));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n13[1]), 
            .I3(n53851), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n53851), .I0(timer[1]), .I1(n13[1]), 
            .CO(n53852));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n13[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n53851));
    SB_LUT4 bit_ctr_0__bdd_4_lut_54971_4_lut_4_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n71849));   // verilog/neopixel.v(65[23:32])
    defparam bit_ctr_0__bdd_4_lut_54971_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 i2215_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(\bit_ctr[0] ), .I3(bit_ctr_c[3]), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2215_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i23391_2_lut_3_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n39155));
    defparam i23391_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1759 (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), 
            .I2(bit_ctr_c[2]), .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1759.LUT_INIT = 16'h1e1e;
    SB_LUT4 i6_3_lut_4_lut (.I0(t1[8]), .I1(t1[5]), .I2(t1[6]), .I3(n56), 
            .O(n14));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2208_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2208_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(\bit_ctr[0] ), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n72113));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 n72113_bdd_4_lut (.I0(n72113), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n72116));
    defparam n72113_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2203_2_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n7200));   // verilog/neopixel.v(65[23:32])
    defparam i2203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n61487), .I2(LED_c), .I3(state[1]), 
            .O(n27639));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i12677_2_lut_4_lut (.I0(state[0]), .I1(n61487), .I2(LED_c), 
            .I3(state[1]), .O(n28538));   // verilog/neopixel.v(35[4] 112[11])
    defparam i12677_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23759_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n39155), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n39530));
    defparam i23759_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1760 (.I0(bit_ctr_c[3]), .I1(n39155), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n55684));
    defparam i1_2_lut_3_lut_adj_1760.LUT_INIT = 16'h7878;
    SB_LUT4 i23244_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n39007));
    defparam i23244_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53194_4_lut (.I0(n39007), .I1(n61), .I2(t1[10]), .I3(n71840), 
            .O(n68464));   // verilog/neopixel.v(19[11:16])
    defparam i53194_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i44_4_lut (.I0(n68464), .I1(state[1]), .I2(start), .I3(n14), 
            .O(n3172));   // verilog/neopixel.v(19[11:16])
    defparam i44_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i2222_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n7200), .I2(bit_ctr_c[3]), 
            .I3(bit_ctr_c[4]), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2222_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i52_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr_c[3]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41));
    defparam i52_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 i3_4_lut_adj_1761 (.I0(n55684), .I1(n41), .I2(bit_ctr[1]), 
            .I3(\bit_ctr[0] ), .O(n23));
    defparam i3_4_lut_adj_1761.LUT_INIT = 16'h0008;
    SB_LUT4 i44457_2_lut (.I0(n23), .I1(n39530), .I2(GND_net), .I3(GND_net), 
            .O(n61487));
    defparam i44457_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1762 (.I0(start), .I1(n59), .I2(GND_net), .I3(GND_net), 
            .O(n35689));   // verilog/neopixel.v(19[11:16])
    defparam i1_2_lut_adj_1762.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(n27639), .I1(n35689), .I2(state[1]), .I3(GND_net), 
            .O(n27645));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13204_2_lut (.I0(n27645), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29064));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_54892 (.I0(color_bit_N_502[1]), .I1(n65374), 
            .I2(n65375), .I3(color_bit_N_502[2]), .O(n71915));
    defparam color_bit_N_502_1__bdd_4_lut_54892.LUT_INIT = 16'he4aa;
    SB_LUT4 n71915_bdd_4_lut (.I0(n71915), .I1(n65372), .I2(n65371), .I3(color_bit_N_502[2]), 
            .O(n71918));
    defparam n71915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48368_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n65458));
    defparam i48368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48369_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n65459));
    defparam i48369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48546_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n65636));
    defparam i48546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48545_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(\bit_ctr[0] ), .I3(GND_net), .O(n65635));
    defparam i48545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2201_2_lut (.I0(bit_ctr[1]), .I1(\bit_ctr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_502[1]));   // verilog/neopixel.v(65[23:32])
    defparam i2201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n71849_bdd_4_lut_4_lut (.I0(color_bit_N_502[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n71849), .O(n71852));   // verilog/neopixel.v(65[23:32])
    defparam n71849_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 i16_2_lut_3_lut (.I0(start), .I1(n59), .I2(\bit_ctr[0] ), 
            .I3(GND_net), .O(n20767));   // verilog/neopixel.v(20[11:18])
    defparam i16_2_lut_3_lut.LUT_INIT = 16'hb4b4;
    SB_LUT4 i12_3_lut_4_lut (.I0(start), .I1(n59), .I2(n1), .I3(state[1]), 
            .O(n28537));   // verilog/neopixel.v(34[12] 113[6])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0f44;
    SB_LUT4 i60_4_lut_4_lut (.I0(t1[1]), .I1(t1[3]), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n43));
    defparam i60_4_lut_4_lut.LUT_INIT = 16'h1880;
    SB_LUT4 i63_4_lut_4_lut (.I0(t1[3]), .I1(t1[1]), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n44));
    defparam i63_4_lut_4_lut.LUT_INIT = 16'h1881;
    SB_LUT4 i85_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n63), .I3(GND_net), .O(n1));
    defparam i85_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i51496_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n39155), .I2(n72020), 
            .I3(GND_net), .O(n68432));
    defparam i51496_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i53814_3_lut_4_lut (.I0(bit_ctr_c[3]), .I1(n39155), .I2(n71918), 
            .I3(n70583), .O(n70904));
    defparam i53814_3_lut_4_lut.LUT_INIT = 16'hf960;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1792, ENCODER0_A_N_keep, 
            \a_new[1] , \b_new[1] , n29238, n1747, n29237, a_prev, 
            n29235, b_prev, position_31__N_3836, \encoder0_position[0] , 
            \encoder0_position[1] , \encoder0_position[2] , \encoder0_position[3] , 
            \encoder0_position[4] , \encoder0_position[5] , \encoder0_position[6] , 
            \encoder0_position[7] , \encoder0_position[8] , \encoder0_position[9] , 
            \encoder0_position[10] , \encoder0_position[11] , \encoder0_position[12] , 
            \encoder0_position[13] , \encoder0_position[14] , \encoder0_position[15] , 
            \encoder0_position[16] , \encoder0_position[17] , \encoder0_position[18] , 
            \encoder0_position[19] , \encoder0_position[20] , \encoder0_position[21] , 
            \encoder0_position[22] , n1765, n1763, n1761, n1759, n1757, 
            n1755, n1753, n1751, n1749, debounce_cnt_N_3833, GND_net, 
            VCC_net) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1792;
    input ENCODER0_A_N_keep;
    output \a_new[1] ;
    output \b_new[1] ;
    input n29238;
    output n1747;
    input n29237;
    output a_prev;
    input n29235;
    output b_prev;
    output position_31__N_3836;
    output \encoder0_position[0] ;
    output \encoder0_position[1] ;
    output \encoder0_position[2] ;
    output \encoder0_position[3] ;
    output \encoder0_position[4] ;
    output \encoder0_position[5] ;
    output \encoder0_position[6] ;
    output \encoder0_position[7] ;
    output \encoder0_position[8] ;
    output \encoder0_position[9] ;
    output \encoder0_position[10] ;
    output \encoder0_position[11] ;
    output \encoder0_position[12] ;
    output \encoder0_position[13] ;
    output \encoder0_position[14] ;
    output \encoder0_position[15] ;
    output \encoder0_position[16] ;
    output \encoder0_position[17] ;
    output \encoder0_position[18] ;
    output \encoder0_position[19] ;
    output \encoder0_position[20] ;
    output \encoder0_position[21] ;
    output \encoder0_position[22] ;
    output n1765;
    output n1763;
    output n1761;
    output n1759;
    output n1757;
    output n1755;
    output n1753;
    output n1751;
    output n1749;
    output debounce_cnt_N_3833;
    input GND_net;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n54616, n54615, n54614, n54613, n54612, 
        n54611, n54610, n54609, n54608, n54607, n54606, n54605, 
        n54604, n54603, n54602, n54601, n54600, n54599, n54598, 
        n54597, n54596, n54595, n54594, n54593, n54592, n54591, 
        n54590, n54589, n54588, n54587, n54586;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1792), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1792), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1792), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1792), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1747), .C(n1792), .D(n29238));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1792), .D(n29237));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1792), .D(n29235));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i0 (.Q(\encoder0_position[0] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(\encoder0_position[1] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(\encoder0_position[2] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(\encoder0_position[3] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(\encoder0_position[4] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(\encoder0_position[5] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(\encoder0_position[6] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(\encoder0_position[7] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(\encoder0_position[8] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(\encoder0_position[9] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(\encoder0_position[10] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(\encoder0_position[11] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(\encoder0_position[12] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(\encoder0_position[13] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(\encoder0_position[14] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(\encoder0_position[15] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(\encoder0_position[16] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(\encoder0_position[17] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(\encoder0_position[18] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(\encoder0_position[19] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(\encoder0_position[20] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(\encoder0_position[21] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(\encoder0_position[22] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(n1765), .C(n1792), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(n1763), .C(n1792), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(n1761), .C(n1792), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(n1759), .C(n1792), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(n1757), .C(n1792), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(n1755), .C(n1792), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(n1753), .C(n1792), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(n1751), .C(n1792), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i31 (.Q(n1749), .C(n1792), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1749), .I3(n54616), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1751), .I3(n54615), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n54615), .I0(direction_N_3840), 
            .I1(n1751), .CO(n54616));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1753), .I3(n54614), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n54614), .I0(direction_N_3840), 
            .I1(n1753), .CO(n54615));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1755), .I3(n54613), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n54613), .I0(direction_N_3840), 
            .I1(n1755), .CO(n54614));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1757), .I3(n54612), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n54612), .I0(direction_N_3840), 
            .I1(n1757), .CO(n54613));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1759), .I3(n54611), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n54611), .I0(direction_N_3840), 
            .I1(n1759), .CO(n54612));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1761), .I3(n54610), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n54610), .I0(direction_N_3840), 
            .I1(n1761), .CO(n54611));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1763), .I3(n54609), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n54609), .I0(direction_N_3840), 
            .I1(n1763), .CO(n54610));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1765), .I3(n54608), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n54608), .I0(direction_N_3840), 
            .I1(n1765), .CO(n54609));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[22] ), .I3(n54607), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n54607), .I0(direction_N_3840), 
            .I1(\encoder0_position[22] ), .CO(n54608));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n54606), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n54606), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n54607));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n54605), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n54605), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n54606));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n54604), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n54604), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n54605));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n54603), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n54603), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n54604));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n54602), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n54602), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n54603));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n54601), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n54601), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n54602));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n54600), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n54600), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n54601));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n54599), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n54599), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n54600));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n54598), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n54598), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n54599));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n54597), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n54597), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n54598));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n54596), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n54596), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n54597));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n54595), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n54595), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n54596));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n54594), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n54594), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n54595));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n54593), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n54593), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n54594));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n54592), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n54592), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n54593));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n54591), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n54591), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n54592));
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n54590), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n54590), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n54591));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n54589), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_6 (.CI(n54589), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n54590));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n54588), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n54588), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n54589));
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n54587), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n54587), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n54588));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n54586), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n54586), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n54587));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n54586));
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (GND_net, n59876, VCC_net, \data_in_frame[23] , clk16MHz, 
            n2881, \data_out_frame[18] , n60534, n60533, n29193, \data_in_frame[11] , 
            n60532, setpoint, reset, n29619, n60531, n28930, n29616, 
            n60530, \data_out_frame[19] , n60474, n60529, n60528, 
            n60527, n60526, n60525, n60524, n60523, \data_out_frame[20] , 
            n60522, rx_data, n60476, n60521, n60520, n60519, \data_out_frame[3][4] , 
            n60646, \data_out_frame[3][6] , n60645, \data_out_frame[3][7] , 
            n60644, n29613, \data_out_frame[4] , n60643, \data_in_frame[1] , 
            n60642, n60658, n60641, n60518, \data_in_frame[8][6] , 
            n17, control_mode, n22, \data_in_frame[8][2] , n60517, 
            n60516, \data_in_frame[20] , \data_out_frame[21] , n60515, 
            n60514, n60513, n60512, n60511, n60510, n60509, n60508, 
            \data_out_frame[22] , n60507, n60506, n60505, n60504, 
            n60503, n60502, n60501, n60500, \data_out_frame[23] , 
            n60499, n60640, n60639, n60638, n60498, n60497, n60496, 
            n60495, n60494, n60493, n60492, n60637, \data_out_frame[24] , 
            n60491, n60490, n25647, \FRAME_MATCHER.i_31__N_2509 , displacement, 
            n60489, \data_in_frame[8][3] , n25732, \data_out_frame[5] , 
            n60636, n60635, n60634, n60633, n60632, \data_in_frame[21] , 
            n60631, n60630, n29196, n60629, \data_out_frame[6] , n60628, 
            n60488, n60627, n60626, n60625, n60542, n60487, n60486, 
            n60485, \data_out_frame[25] , n60484, n60483, n60482, 
            n60481, n60480, n60479, control_update, n27465, \data_out_frame[7] , 
            \encoder0_position_scaled[12] , n60478, n60477, \encoder0_position_scaled[11] , 
            \encoder0_position_scaled[10] , \FRAME_MATCHER.i[5] , \FRAME_MATCHER.i[4] , 
            \encoder0_position_scaled[9] , \FRAME_MATCHER.i[3] , n60624, 
            byte_transmit_counter, n60623, \encoder0_position_scaled[8] , 
            n161, \data_in_frame[16] , \data_in_frame[18] , \encoder0_position_scaled[23] , 
            \FRAME_MATCHER.state[3] , n60543, \encoder0_position_scaled[22] , 
            n28096, n8, tx_active, n31, n60622, pwm_setpoint, \pwm_counter[15] , 
            n31_adj_10, \data_in_frame[10] , n60621, \pwm_counter[16] , 
            n33, n29199, n60620, n29020, n60619, \data_in_frame[8][7] , 
            \data_in_frame[17] , n60896, \data_out_frame[8][6] , \control_mode[6] , 
            n48532, \control_mode[2] , \control_mode[4] , \data_in_frame[2] , 
            n29520, n29513, n59920, \encoder0_position_scaled[21] , 
            \data_out_frame[0][2] , \data_in_frame[1][2] , n59922, n29205, 
            n29501, n29498, n29495, n29492, n29489, n29486, n29483, 
            n29480, n29477, n29208, n29473, n60618, n29211, n29214, 
            n29466, n29463, n29460, n29459, n29456, n60617, n29451, 
            n29448, n68429, n29445, n29442, n29439, n29436, n60616, 
            \data_in_frame[14][6] , \data_out_frame[8][1] , n60615, \data_out_frame[17] , 
            n60657, \data_out_frame[0][3] , n60656, \data_out_frame[0][4] , 
            n60655, \data_out_frame[1][0] , n60654, \data_out_frame[1][1] , 
            n60653, \data_out_frame[1][3] , n60652, \data_out_frame[1][5] , 
            n60651, \data_out_frame[1][6] , n60650, \data_out_frame[1][7] , 
            n60649, \data_out_frame[3][1] , n60648, \data_out_frame[3][3] , 
            n60647, \data_out_frame[8][2] , n60614, \data_out_frame[8][3] , 
            n60613, \data_out_frame[8][4] , n60612, \data_out_frame[8][5] , 
            n60611, n60610, \data_out_frame[8][7] , n60609, \data_out_frame[9] , 
            n60608, n60607, n60606, n60605, n60604, n60603, n29002, 
            n60602, \data_out_frame[10] , n60601, n60600, n60599, 
            n60598, n60597, n60596, n60595, n60594, \data_out_frame[11] , 
            n60593, n60592, n60591, n60590, n60589, n60588, n60587, 
            n60586, \data_out_frame[12] , n60585, n60584, n60583, 
            n60582, n60581, n60580, n60579, n60578, \data_out_frame[13] , 
            n60577, n60576, n60575, n60574, n60573, n60572, n60571, 
            n60570, \data_out_frame[14] , n60569, n60568, n60567, 
            n60566, n60565, n60564, n60563, n60562, \data_out_frame[15] , 
            n60561, n60560, n60559, n60558, n60557, n60556, n60555, 
            n60554, \data_out_frame[16] , n60553, n60475, n60552, 
            n60551, n60550, n60549, n60548, n60547, n60546, n60545, 
            n29236, \FRAME_MATCHER.rx_data_ready_prev , n60544, n60541, 
            n60540, n60539, LED_c, n8_adj_11, DE_c, \data_in_frame[1][6] , 
            n39467, n3483, n37935, n60700, n60538, n56640, n72152, 
            n60537, n59930, deadband, IntegralLimit, \Kp[0] , \Ki[0] , 
            PWMLimit, n29629, n29632, n29635, n29948, n29945, n29942, 
            n29939, n29936, n29933, n29930, n29927, n29127, n29130, 
            n29133, \data_in_frame[8][4] , n56696, n29136, \data_in_frame[8][5] , 
            n29139, n29142, \Kp[1] , \Kp[2] , \Kp[3] , \Kp[4] , 
            \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , \Kp[10] , 
            \Kp[11] , \Kp[12] , \Kp[13] , n60536, \Kp[14] , \Kp[15] , 
            \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , 
            \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , \Ki[12] , 
            \Ki[13] , \Ki[14] , \Ki[15] , neopxl_color, n60535, n29739, 
            n29738, n29736, n29734, n29733, \control_mode[7] , n29732, 
            current_limit, n29731, n29730, n29729, n29728, n29727, 
            n29726, n29725, n29724, n29723, n29722, n29721, n29720, 
            n29719, n29718, n29110, n29172, \data_in_frame[10][1] , 
            n29175, \data_in_frame[10][2] , n29178, \data_in_frame[10][3] , 
            n29181, n29184, n29187, n29190, n39431, n110, n112, 
            n37941, n68422, \encoder0_position_scaled[20] , rx_data_ready, 
            n24820, n34686, n34584, n62686, encoder1_position_scaled, 
            n56501, n56624, n56565, n25994, n55945, n61288, n26215, 
            n60951, n55578, n61213, \encoder0_position_scaled[7] , \encoder0_position_scaled[6] , 
            \encoder0_position_scaled[5] , \encoder0_position_scaled[4] , 
            \encoder0_position_scaled[3] , \encoder0_position_scaled[2] , 
            n61461, n26311, n56545, n31_adj_12, n25712, n61442, 
            \encoder0_position_scaled[1] , n61245, n22465, n28, n6, 
            n28102, n60771, n60766, n8_adj_13, n115, ID, \encoder0_position_scaled[19] , 
            \encoder0_position_scaled[18] , \encoder0_position_scaled[17] , 
            \encoder0_position_scaled[16] , n72092, \encoder0_position_scaled[15] , 
            n72086, n72122, n71906, \encoder0_position_scaled[14] , 
            \current[7] , \current[6] , \current[5] , \current[4] , 
            \current[3] , \current[2] , \encoder0_position_scaled[13] , 
            \current[1] , \current[0] , \current[15] , \current[11] , 
            \current[10] , \current[9] , \current[8] , n61134, n72026, 
            n15, n7, n31_adj_14, n15_adj_15, n15_adj_16, r_SM_Main, 
            \r_SM_Main_2__N_3536[1] , n1, tx_o, \tx_data[0] , n5227, 
            \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , n29, n23, n62322, 
            n27, \r_Bit_Index[0] , n60413, n63831, r_Clock_Count, 
            n27514, n29671, n61481, n29123, n72442, n63819, n6_adj_17, 
            tx_enable, baudrate, r_Rx_Data, r_SM_Main_adj_31, \r_SM_Main_2__N_3446[1] , 
            n5224, \o_Rx_DV_N_3488[8] , RX_N_2, n25296, r_Clock_Count_adj_32, 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[7] , \r_Bit_Index[0]_adj_29 , n60415, n63843, 
            n27507, n27511, n29674, n56754, n29679, n29646, n29645, 
            n29644, n29642, n29641, n29640, n29639, n61483, n6_adj_30, 
            \o_Rx_DV_N_3488[0] , n64131, n64079, n64167, n64205, n64169, 
            n64151, n64133, n64097, n4, n63821) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n59876;
    input VCC_net;
    output [7:0]\data_in_frame[23] ;
    input clk16MHz;
    input n2881;
    output [7:0]\data_out_frame[18] ;
    input n60534;
    input n60533;
    input n29193;
    output [7:0]\data_in_frame[11] ;
    input n60532;
    output [23:0]setpoint;
    input reset;
    input n29619;
    input n60531;
    input n28930;
    input n29616;
    input n60530;
    output [7:0]\data_out_frame[19] ;
    input n60474;
    input n60529;
    input n60528;
    input n60527;
    input n60526;
    input n60525;
    input n60524;
    input n60523;
    output [7:0]\data_out_frame[20] ;
    input n60522;
    output [7:0]rx_data;
    input n60476;
    input n60521;
    input n60520;
    input n60519;
    output \data_out_frame[3][4] ;
    input n60646;
    output \data_out_frame[3][6] ;
    input n60645;
    output \data_out_frame[3][7] ;
    input n60644;
    input n29613;
    output [7:0]\data_out_frame[4] ;
    input n60643;
    output [7:0]\data_in_frame[1] ;
    input n60642;
    input n60658;
    input n60641;
    input n60518;
    output \data_in_frame[8][6] ;
    output n17;
    output [7:0]control_mode;
    output n22;
    output \data_in_frame[8][2] ;
    input n60517;
    input n60516;
    output [7:0]\data_in_frame[20] ;
    output [7:0]\data_out_frame[21] ;
    input n60515;
    input n60514;
    input n60513;
    input n60512;
    input n60511;
    input n60510;
    input n60509;
    input n60508;
    output [7:0]\data_out_frame[22] ;
    input n60507;
    input n60506;
    input n60505;
    input n60504;
    input n60503;
    input n60502;
    input n60501;
    input n60500;
    output [7:0]\data_out_frame[23] ;
    input n60499;
    input n60640;
    input n60639;
    input n60638;
    input n60498;
    input n60497;
    input n60496;
    input n60495;
    input n60494;
    input n60493;
    input n60492;
    input n60637;
    output [7:0]\data_out_frame[24] ;
    input n60491;
    input n60490;
    output n25647;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]displacement;
    input n60489;
    output \data_in_frame[8][3] ;
    output n25732;
    output [7:0]\data_out_frame[5] ;
    input n60636;
    input n60635;
    input n60634;
    input n60633;
    input n60632;
    output [7:0]\data_in_frame[21] ;
    input n60631;
    input n60630;
    input n29196;
    input n60629;
    output [7:0]\data_out_frame[6] ;
    input n60628;
    input n60488;
    input n60627;
    input n60626;
    input n60625;
    input n60542;
    input n60487;
    input n60486;
    input n60485;
    output [7:0]\data_out_frame[25] ;
    input n60484;
    input n60483;
    input n60482;
    input n60481;
    input n60480;
    input n60479;
    input control_update;
    output n27465;
    output [7:0]\data_out_frame[7] ;
    input \encoder0_position_scaled[12] ;
    input n60478;
    input n60477;
    input \encoder0_position_scaled[11] ;
    input \encoder0_position_scaled[10] ;
    output \FRAME_MATCHER.i[5] ;
    output \FRAME_MATCHER.i[4] ;
    input \encoder0_position_scaled[9] ;
    output \FRAME_MATCHER.i[3] ;
    input n60624;
    output [7:0]byte_transmit_counter;
    input n60623;
    input \encoder0_position_scaled[8] ;
    output n161;
    output [7:0]\data_in_frame[16] ;
    output [7:0]\data_in_frame[18] ;
    input \encoder0_position_scaled[23] ;
    output \FRAME_MATCHER.state[3] ;
    input n60543;
    input \encoder0_position_scaled[22] ;
    output n28096;
    output n8;
    output tx_active;
    input n31;
    input n60622;
    input [23:0]pwm_setpoint;
    input \pwm_counter[15] ;
    output n31_adj_10;
    output [7:0]\data_in_frame[10] ;
    input n60621;
    input \pwm_counter[16] ;
    output n33;
    input n29199;
    input n60620;
    input n29020;
    input n60619;
    output \data_in_frame[8][7] ;
    output [7:0]\data_in_frame[17] ;
    input n60896;
    output \data_out_frame[8][6] ;
    output \control_mode[6] ;
    output n48532;
    output \control_mode[2] ;
    output \control_mode[4] ;
    output [7:0]\data_in_frame[2] ;
    input n29520;
    input n29513;
    input n59920;
    input \encoder0_position_scaled[21] ;
    output \data_out_frame[0][2] ;
    output \data_in_frame[1][2] ;
    input n59922;
    input n29205;
    input n29501;
    input n29498;
    input n29495;
    input n29492;
    input n29489;
    input n29486;
    input n29483;
    input n29480;
    input n29477;
    input n29208;
    input n29473;
    input n60618;
    input n29211;
    input n29214;
    input n29466;
    input n29463;
    input n29460;
    input n29459;
    input n29456;
    input n60617;
    input n29451;
    input n29448;
    input n68429;
    input n29445;
    input n29442;
    input n29439;
    input n29436;
    input n60616;
    output \data_in_frame[14][6] ;
    output \data_out_frame[8][1] ;
    input n60615;
    output [7:0]\data_out_frame[17] ;
    input n60657;
    output \data_out_frame[0][3] ;
    input n60656;
    output \data_out_frame[0][4] ;
    input n60655;
    output \data_out_frame[1][0] ;
    input n60654;
    output \data_out_frame[1][1] ;
    input n60653;
    output \data_out_frame[1][3] ;
    input n60652;
    output \data_out_frame[1][5] ;
    input n60651;
    output \data_out_frame[1][6] ;
    input n60650;
    output \data_out_frame[1][7] ;
    input n60649;
    output \data_out_frame[3][1] ;
    input n60648;
    output \data_out_frame[3][3] ;
    input n60647;
    output \data_out_frame[8][2] ;
    input n60614;
    output \data_out_frame[8][3] ;
    input n60613;
    output \data_out_frame[8][4] ;
    input n60612;
    output \data_out_frame[8][5] ;
    input n60611;
    input n60610;
    output \data_out_frame[8][7] ;
    input n60609;
    output [7:0]\data_out_frame[9] ;
    input n60608;
    input n60607;
    input n60606;
    input n60605;
    input n60604;
    input n60603;
    input n29002;
    input n60602;
    output [7:0]\data_out_frame[10] ;
    input n60601;
    input n60600;
    input n60599;
    input n60598;
    input n60597;
    input n60596;
    input n60595;
    input n60594;
    output [7:0]\data_out_frame[11] ;
    input n60593;
    input n60592;
    input n60591;
    input n60590;
    input n60589;
    input n60588;
    input n60587;
    input n60586;
    output [7:0]\data_out_frame[12] ;
    input n60585;
    input n60584;
    input n60583;
    input n60582;
    input n60581;
    input n60580;
    input n60579;
    input n60578;
    output [7:0]\data_out_frame[13] ;
    input n60577;
    input n60576;
    input n60575;
    input n60574;
    input n60573;
    input n60572;
    input n60571;
    input n60570;
    output [7:0]\data_out_frame[14] ;
    input n60569;
    input n60568;
    input n60567;
    input n60566;
    input n60565;
    input n60564;
    input n60563;
    input n60562;
    output [7:0]\data_out_frame[15] ;
    input n60561;
    input n60560;
    input n60559;
    input n60558;
    input n60557;
    input n60556;
    input n60555;
    input n60554;
    output [7:0]\data_out_frame[16] ;
    input n60553;
    input n60475;
    input n60552;
    input n60551;
    input n60550;
    input n60549;
    input n60548;
    input n60547;
    input n60546;
    input n60545;
    input n29236;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n60544;
    input n60541;
    input n60540;
    input n60539;
    output LED_c;
    output n8_adj_11;
    output DE_c;
    output \data_in_frame[1][6] ;
    output n39467;
    output n3483;
    output n37935;
    output n60700;
    input n60538;
    output n56640;
    output n72152;
    input n60537;
    input n59930;
    output [23:0]deadband;
    output [23:0]IntegralLimit;
    output \Kp[0] ;
    output \Ki[0] ;
    output [23:0]PWMLimit;
    input n29629;
    input n29632;
    input n29635;
    input n29948;
    input n29945;
    input n29942;
    input n29939;
    input n29936;
    input n29933;
    input n29930;
    input n29927;
    input n29127;
    input n29130;
    input n29133;
    output \data_in_frame[8][4] ;
    output n56696;
    input n29136;
    output \data_in_frame[8][5] ;
    input n29139;
    input n29142;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    output \Kp[13] ;
    input n60536;
    output \Kp[14] ;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    output [23:0]neopxl_color;
    input n60535;
    input n29739;
    input n29738;
    input n29736;
    input n29734;
    input n29733;
    output \control_mode[7] ;
    input n29732;
    output [15:0]current_limit;
    input n29731;
    input n29730;
    input n29729;
    input n29728;
    input n29727;
    input n29726;
    input n29725;
    input n29724;
    input n29723;
    input n29722;
    input n29721;
    input n29720;
    input n29719;
    input n29718;
    input n29110;
    input n29172;
    output \data_in_frame[10][1] ;
    input n29175;
    output \data_in_frame[10][2] ;
    input n29178;
    output \data_in_frame[10][3] ;
    input n29181;
    input n29184;
    input n29187;
    input n29190;
    input n39431;
    input n110;
    output n112;
    output n37941;
    output n68422;
    input \encoder0_position_scaled[20] ;
    output rx_data_ready;
    input n24820;
    output n34686;
    output n34584;
    input n62686;
    input [23:0]encoder1_position_scaled;
    output n56501;
    input n56624;
    input n56565;
    output n25994;
    input n55945;
    output n61288;
    output n26215;
    output n60951;
    output n55578;
    input n61213;
    input \encoder0_position_scaled[7] ;
    input \encoder0_position_scaled[6] ;
    input \encoder0_position_scaled[5] ;
    input \encoder0_position_scaled[4] ;
    input \encoder0_position_scaled[3] ;
    input \encoder0_position_scaled[2] ;
    output n61461;
    input n26311;
    output n56545;
    output n31_adj_12;
    output n25712;
    input n61442;
    input \encoder0_position_scaled[1] ;
    input n61245;
    output n22465;
    input n28;
    output n6;
    output n28102;
    output n60771;
    output n60766;
    output n8_adj_13;
    input n115;
    input [7:0]ID;
    input \encoder0_position_scaled[19] ;
    input \encoder0_position_scaled[18] ;
    input \encoder0_position_scaled[17] ;
    input \encoder0_position_scaled[16] ;
    output n72092;
    input \encoder0_position_scaled[15] ;
    output n72086;
    input n72122;
    input n71906;
    input \encoder0_position_scaled[14] ;
    input \current[7] ;
    input \current[6] ;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \encoder0_position_scaled[13] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    input n61134;
    input n72026;
    output n15;
    output n7;
    output n31_adj_14;
    output n15_adj_15;
    output n15_adj_16;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    output n1;
    output tx_o;
    input \tx_data[0] ;
    input n5227;
    output \o_Rx_DV_N_3488[12] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    input n62322;
    output n27;
    output \r_Bit_Index[0] ;
    output n60413;
    input n63831;
    output [8:0]r_Clock_Count;
    output n27514;
    input n29671;
    output n61481;
    input n29123;
    input n72442;
    output n63819;
    output n6_adj_17;
    output tx_enable;
    input [31:0]baudrate;
    output r_Rx_Data;
    output [2:0]r_SM_Main_adj_31;
    input \r_SM_Main_2__N_3446[1] ;
    input n5224;
    output \o_Rx_DV_N_3488[8] ;
    input RX_N_2;
    output n25296;
    output [7:0]r_Clock_Count_adj_32;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0]_adj_29 ;
    output n60415;
    input n63843;
    output n27507;
    output n27511;
    input n29674;
    input n56754;
    input n29679;
    input n29646;
    input n29645;
    input n29644;
    input n29642;
    input n29641;
    input n29640;
    input n29639;
    output n61483;
    output n6_adj_30;
    output \o_Rx_DV_N_3488[0] ;
    input n64131;
    output n64079;
    input n64167;
    output n64205;
    output n64169;
    output n64151;
    output n64133;
    output n64097;
    output n4;
    output n63821;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n54525, n28031;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire n54526;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    
    wire n64693, n2, n2_adj_5297, n10, n61254, n25746, n16;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    
    wire n18, n2_adj_5298;
    wire [23:0]n4939;
    
    wire n27414, n2_adj_5299, n2_adj_5300, n2_adj_5301, n2_adj_5302, 
        n2_adj_5303, n2_adj_5304, n2_adj_5305, n2_adj_5306, n2_adj_5307, 
        n27778, n54524, n68360, n2_adj_5308, n25598, n60855, n61415, 
        n26126, n17_c, n2_adj_5309, n2_adj_5310, n8_c, n60760;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    
    wire n29999, n2_adj_5311, n2_adj_5312, n2_adj_5313, n30002, n2_adj_5314, 
        n30005, n2_adj_5315, n27776, n54523, n68363, n2_adj_5316, 
        n30008, n2_adj_5317, n30011, n2_adj_5318;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    
    wire n60890, n10_adj_5319, n2_adj_5320, n30014, n30017, n2_adj_5321, 
        n30020, n29610;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5322, n2_adj_5323, n56705, Kp_23__N_974, n65144, n21, 
        n26220, n26250, n56127, n26089, n65225, n25718, n26621, 
        n4_c, n2_adj_5325, n2_adj_5326, n8_adj_5327, n60740, n29539, 
        n2_adj_5328, n2_adj_5329, n2_adj_5330, n2_adj_5331, n29542, 
        n29545, n2_adj_5332, n2_adj_5333, n2_adj_5334, n2_adj_5335, 
        n2_adj_5336, n2_adj_5337, n2_adj_5338, n2_adj_5339, n2_adj_5340, 
        n2_adj_5341, n2_adj_5342, n2_adj_5343, n2_adj_5344, n2_adj_5345, 
        n2_adj_5346, n29607, n2_adj_5347, n2_adj_5348, n2_adj_5349, 
        n2_adj_5350, n2_adj_5351, n2_adj_5352, n2_adj_5353, n2_adj_5354, 
        n56707;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n18_adj_5355, n29604, n2_adj_5356, n2_adj_5357, n2_adj_5358, 
        n29549, n26077, n71572, n7_c, n26;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5359, n2_adj_5360, n29601, Kp_23__N_869, n65247, n29552, 
        n29555, n27774, n54522, n68364, n27772, n54521, n68365, 
        n2_adj_5361, n29598, n2_adj_5362, n29595, n2_adj_5363, n29592, 
        n2_adj_5364, n29589, n8_adj_5365, n29586, n29558, n2_adj_5366, 
        n29583, n2_adj_5367, n2_adj_5368, n29579, n2_adj_5369, n2_adj_5370, 
        n29576, n2_adj_5371, n29573, n2_adj_5372, n29570, n2_adj_5373, 
        n2_adj_5374, n2_adj_5375, n2_adj_5376, n29567, n2_adj_5377, 
        n2_adj_5378, n2_adj_5379, n2_adj_5380, n2_adj_5381, n2_adj_5382, 
        n2_adj_5383, n29561, n37468, n2_adj_5384, n29564, n17_adj_5385, 
        n25249, n2_adj_5386, n2_adj_5387, n2_adj_5388, n3;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n60693, n3_adj_5389, n60690, n3_adj_5390, n60689, n2_adj_5391, 
        n3_adj_5392, n60688, n27770, n54520, n68366, n3_adj_5393, 
        n60687, n3_adj_5394, n60680, n3_adj_5395, n60694, n27768, 
        n54519, n68367, n27766, n54518, n68369, n3_adj_5396, n60683, 
        n3_adj_5397;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n60691, n3_adj_5398, n60682, n2_adj_5399, n27764, n54517, 
        n68375, n27762, n54516, n68377, n3_adj_5400, n60681, n2_adj_5401, 
        n27760, n54515, n68380, n3_adj_5402, n60685, n3_adj_5403, 
        n60686, n3_adj_5404, n60679, n70567, n68462, n72059, n71954, 
        n7_adj_5405;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n2_adj_5406, n2_adj_5407;
    wire [31:0]n133;
    
    wire Kp_23__N_1067, n29975, n3_adj_5408, n60692, n29978, n61335, 
        n56563, Kp_23__N_1271, n61439, n70513, n68444, n72047, n3_adj_5409, 
        n60684, n2075, Kp_23__N_1748, n71936, n65337, n29981, n29984, 
        n61310, n10_adj_5410, n2_adj_5411, n1_c, n60673, n29987, 
        n29990, n1_adj_5412, n60672, n60785, n55989, n29993, n29996, 
        n71960, n72134, n70710, n71870, \FRAME_MATCHER.i_31__N_2511 , 
        n1_adj_5413, \FRAME_MATCHER.i_31__N_2514 , n60730;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n1_adj_5414, n1_adj_5415, n60671, n1_adj_5416, n60670, n1_adj_5417, 
        n60669, n1_adj_5418, n60668, n72041, n1958, n62539, n4452, 
        n20871, n22473, n64994, n26846, n3303, \FRAME_MATCHER.i_31__N_2512 , 
        n2067, n60674, Kp_23__N_1080, n64711, n72396, \FRAME_MATCHER.i_31__N_2507 , 
        n26843, \FRAME_MATCHER.i_31__N_2508 , n2_adj_5419, n2055, n2056, 
        n20876, n59808, \FRAME_MATCHER.i_31__N_2513 , n1961, n1964, 
        n64990, n62727, n1962, n25260, n771, n5, n60128, n25281, 
        n25150;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n60833, n27402, n63171, n25265;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n6_c;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n6_adj_5421, n25313, n20, n25163;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n19, n24870, n60985, n60987, n65189, n25394, n18_adj_5422, 
        n25325, n20_adj_5423, n15_c;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n39028, n4_adj_5424, n4_adj_5425, n39534, n32327, n16_adj_5426, 
        n17_adj_5427, n10_adj_5428, n14, n15_adj_5429, n16_adj_5430, 
        n17_adj_5431, n62533, n6_adj_5432, n72044, n26178, n55997, 
        n6_adj_5434, n61412;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    
    wire n60969;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    
    wire n25501, n29536;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    
    wire n29533, n29530, n29527, n29524, n29521, n23700, n60979, 
        n26123, Kp_23__N_878, n56744, n56678, n56555;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n25825, n61313, n60858, n37, n55521;
    wire [7:0]control_mode_c;   // verilog/TinyFPGA_B.v(246[14:26])
    
    wire n44, n42, n43, n41, n40, n39, n50, n45, n61326, n61012, 
        n56505, n56535, n25564, n56675, n60816, n72080, n71978, 
        n62519, n6_adj_5435, n60825, n61030, n26057, n61433, n29517, 
        n26120, n26447, n61329, n26154, n25591, n26451, n60841, 
        n29514, n55574, n61129, n60871, n56614, n61125, n61104, 
        n60837, Kp_23__N_772, n61261, n68446, n26274, n56634, n56529, 
        n25687, n65354, n65355, n65353, n72140, n61122, n64917, 
        n72188, n71876, n64873, n25987, n63380, n61458, n64921, 
        n61361, n64925, n5_adj_5436, n56559, n62964, n26599, n8_adj_5437, 
        n29951, n2_adj_5438, n29217, n29220, n6_adj_5439, n2_adj_5440, 
        n70717, n72209, n29433, n29954, n29430, n29427, n29424, 
        n2_adj_5441, n29421, n29418, n29415, n29412, n29409;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    
    wire n29406, n29403, n29400, n29397, n25658, n61048, n60927, 
        n64931, n29394, n71924, n7_adj_5442, n29224, n29229, n29232, 
        n29240, n23704, n63425, n65623, n65624, n72005, n65309, 
        n65308, n72008, n29243, n29957, n29246, n29249, n61436, 
        n64933, n64939, n70699, n68453, n72197, n29252, n29255, 
        n29258, n29261, n29264, n29267, n29270, n29273, n29276, 
        n61141, n24953, n29960, n29963, n29966, n29969, n2_adj_5443, 
        n55540, n55580, n64961, n60903, n25817, n56075, n6_adj_5444, 
        n56684, n55705, n55503, n60960, n60880, n60932, n61201, 
        n61018, n61295, n14_adj_5445, n60828, n13, n10_adj_5446, 
        n61455, n12, n14_adj_5447, n10_adj_5448, n25556, n71987, 
        n29972, n25950, n60963, n60118, n56561, n61107, n6_adj_5449, 
        n60822, Kp_23__N_1389, n10_adj_5450, n61178, n64883, Kp_23__N_1518, 
        n61388, n61174, n61367, n7_adj_5451, n71990, n61282, n5_adj_5452, 
        n2_adj_5453, n2_adj_5454, n2_adj_5455, n2_adj_5456, n2_adj_5457, 
        n2_adj_5458, n2_adj_5459, n2_adj_5460, n2_adj_5461, n2_adj_5462, 
        n2_adj_5463, n2_adj_5464, n2_adj_5465, n2_adj_5466, n2_adj_5467, 
        n2_adj_5468, n2_adj_5469, n2_adj_5470, n2_adj_5471, n2_adj_5472, 
        n2_adj_5473, n2_adj_5474, n2_adj_5475, n2_adj_5476, n2_adj_5477, 
        n2_adj_5478, n2_adj_5479, n2_adj_5480, n2_adj_5481, n2_adj_5482, 
        n2_adj_5483, n2_adj_5484, n2_adj_5485, n2_adj_5486, n2_adj_5487, 
        n2_adj_5488, n2_adj_5489, n2_adj_5490, n2_adj_5491, n2_adj_5492, 
        n2_adj_5493, n2_adj_5494, n2_adj_5495, n2_adj_5496, n2_adj_5497, 
        n2_adj_5498, n2_adj_5499, n29309, n2_adj_5500, n29308, n2_adj_5501, 
        n29307, n2_adj_5502, n29306, n2_adj_5503, n29305, n2_adj_5504, 
        n29304, n2_adj_5505, n29303, n2_adj_5506, n29302, n2_adj_5507, 
        n29301, n2_adj_5508, n29300, n2_adj_5509, n29299, n2_adj_5510, 
        n29298, n2_adj_5511, n29297, n2_adj_5512, n29296, n2_adj_5513, 
        n29295, n2_adj_5514, n29294, n2_adj_5515, n29293, n2_adj_5516, 
        n29292, n2_adj_5517, n29291, n2_adj_5518, n29290, n2_adj_5519, 
        n29289, n2_adj_5520, n29288, n2_adj_5521, n29287, n2_adj_5522, 
        n29286, n2_adj_5523, n29285, n2_adj_5524, n29284, n2_adj_5525, 
        n29283, n29282, n2_adj_5526, n29281, n29280, n29279, n2_adj_5527, 
        n2_adj_5528, n2_adj_5529, n2_adj_5530, n2_adj_5531, n2_adj_5532, 
        n2_adj_5533, n2_adj_5534, n2_adj_5535, n2_adj_5536, n68321, 
        n2_adj_5537, n2_adj_5538, n2_adj_5539, n2_adj_5540, n72191, 
        n9, n12_adj_5541, n11, n68319, n68320, n5_adj_5542, n4_adj_5543, 
        n72194, n61323, n65402, n27827, n65403, n65401, n72104, 
        n68434, n55137, n61344, n65016, n60947, n61298, n62580, 
        n63286, n62654, n6_adj_5544, n63297, n64829, n4_adj_5545, 
        n64831, n6_adj_5546, n63036, n56596, n64835, n55682, n62755, 
        n27733, n72110, n70681, n5_adj_5547, n28610, n25765, n29903, 
        n26729, n28603, n64903, n60966, n64839, n55692, n64841, 
        n25461, n1244, n1_adj_5549, n28599, n60993, Kp_23__N_872, 
        n6_adj_5550, n29906, n8_adj_5551, n61285, n60906, n62556, 
        n29909, n29912, n61355, n62822, n1516, n72185, n63143, 
        n26198, n64705, n29915, n29918, n71975, n2_adj_5552, n29921, 
        n29924, n60667, n61267, n62899, n72179, n64645, n64647, 
        n61098, n64657, n72182, n60861, n60844, n64659, n25540, 
        n64665, n61224, n63034, n64663, n64671, n64685, n25669, 
        n55544, n64783, n56575, n64909, n60990, n64791, n63330, 
        n60883, n64793, n72167, n71930, n7_adj_5553, n64799, n72161, 
        n65333, n61198, n61102, n64805, n72155, n55511, n61185, 
        n60973, n64811, n72149, n61381, n64817, n72143, n55970, 
        n72146, n10_adj_5554, n59688, n64845, n64881, n61051, n62406, 
        n33_adj_5555, n29104, n29105, n29106, n29107;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29111, n29694, n29098, n29680, n30065, n30062, n30059, 
        n30056, n30053, n30050, n30047, n30044, n30041, n30038, 
        n30035, n30032, n30029, n30026, n30023, n29695, n29900, 
        n29897, n29894, n29891, n29888, n29885, n29882, n61113, 
        n56591, n56507, n72137, n55576, n29838, n29837, n29836, 
        n29835, n29834, n29833, n29832, n29831, n29830, n29829, 
        n29828, n29827, n29826, n29825, n29696, n56581, n10_adj_5556, 
        n29824, n29823, n29822, n29821, n29820, n29819, n29818, 
        n29817, n29816, n29815, n29814, n29813, n29812, n29811, 
        n29810, n29809, n29808, n29807, n29806, n29805, n29804, 
        n29803, n29802, n29801, n29800, n29799, n29798, n29797, 
        n29796, n29795, n29794, n29793, n29792, n29791, n29790, 
        n29789, n29788, n29787, n29786, n29785, n29784, n29783, 
        n29782, n29781, n29780, n29697, n29779, n29778, n29777, 
        n29776, n29775, n29774, n29773, n29772, n29771, n29770, 
        n29769, n29768, n29698, n29767, n29766, n29765, n29764, 
        n29763, n29762, n29761, n64765, n64771, n29760, n29759, 
        n29758, n29757, n55700, n26262, n29756, n26258, n29755, 
        n29754, n29753, n61119, n29752, n29751, n29750, n29749, 
        n29748, n29747, n61332, n29746, n29745, n29744, n29743, 
        n29121, n29700, n2_adj_5557, n29742, n29741, n29740, n29737, 
        n29735, n29717, n29716, n29715, n29714, n29713, n29712, 
        n12_adj_5558, n27780, n27782, n27784, n27786, n27788, n27790, 
        n27792, n27794, n27796, n27798, n27800, n27802, n27804, 
        n27806, n27808, n27810, n27812, n27814, n27816, n27818, 
        n27820, n29711, n29710, n29709, n29708, n29707, n29706, 
        n29705, n29704, n29703, n29702, n29701, n29145, n29148, 
        n29151, n29154, n29157, n29160, n29109, n29108, n29163, 
        n61430, n25662, n71568, n18_adj_5559, n29166, n29169, n60924, 
        n61352, n19_adj_5560, n25781, Kp_23__N_1301, n60996, n60938, 
        n16_adj_5561, n17_adj_5562, tx_transmit_N_3416, n25923, n55679, 
        n61073, n6_adj_5563, n27713, n65348, n65349, n65347, n68456, 
        n71948, n70569, n1_adj_5564, n65332, n65383, n65384, n65456, 
        n65455, n65389, n65390, n65438, n65437, n65425, n65426, 
        n65393, n65392, n65452, n65453, n65465, n65464, n65434, 
        n65435, n65342, n65341, n68359, n6_adj_5565, n68358, n68357, 
        n68346, n68345, n32330, n68342, n68337, n68332, n68295, 
        n68294, n68293, n68278, n68273, n68269, n68268, n68267, 
        n68265, n68264, n68263, n68262, n68261, n64849, n64677, 
        n64851, n61027, n53699, n60666, n53698, n53697, n32326, 
        n53696, n53695, n53694, n53693, n60940, n59626, n55617, 
        n61301, n64729, n54545, n54544, n54543, n54542, n54541, 
        n60779, n6_adj_5566, n54540, Kp_23__N_799, n54539, n54538, 
        n54537, n54536, n54535, n72131, n54534, n54533, n54532, 
        n54531, n10_adj_5567, n60769, n54530, n5_adj_5568, n63365, 
        n63147, n56541, n6_adj_5569, n60790, n6_adj_5570, n60900, 
        n61137, n55646, n63372, n61452, n55517, n14_adj_5571, n56573, 
        n25874, n55696, n15_adj_5572, n72125, n61378, n61195, n65364, 
        n61216, n55893, n26398, n61427, n61009, n61349, n14_adj_5573, 
        n26560, n61375, n61307, n26555, n13_adj_5574, n55519, n14_adj_5575, 
        n60957, n15_adj_5576, n55631, n7_adj_5577, n62513, n55598, 
        n61251, n62642, n61421, n4_adj_5578, n61156, n62684, n56626, 
        n10_adj_5579, n61227, n56578, n61233, n10_adj_5580, n18_adj_5581, 
        n25927, n6_adj_5582, n61188, n55650, n25465, n54529, n61385, 
        n60793, n61230, n55644, n6_adj_5583, n55639, n12_adj_5584, 
        n55515, n61089, n20_adj_5585, n56632, n55534, n56492, n19_adj_5586, 
        n62914, n21_adj_5587, n54528, n26_adj_5588, n54527, n34, 
        n60819, n61042, n32, n31_adj_5589, n55731, n35, n37_adj_5590, 
        n61110, n61358, n10_adj_5591, n6_adj_5592, n56543, n61207, 
        n25879, n14_adj_5593, n61006, n61391, n6_adj_5594, n6_adj_5595, 
        n55523, n4_adj_5596, n55741, n55368, n26185, n61147, n1168, 
        n60864, n10_adj_5597, n1130, n8_adj_5598, n61181, n10_adj_5599, 
        n62824, n61150, n26405, n14_adj_5600, n61039, n61062, n61418, 
        n61291, n10_adj_5601, n26147, n23471, n61000, n60850, n60803, 
        n9_adj_5602, n61276, n61159, n56069, n23430, n61273, n26304, 
        n61364, n10_adj_5603, n55499, n61024, n6_adj_5604, n56583, 
        n6_adj_5605, n60944, n10_adj_5606, n55715, n25490, n6_adj_5607, 
        n24849, n10_adj_5608, n56537, n61162, n6_adj_5609, n60867, 
        n61270, n7_adj_5610, n56192, n62635, n62923, n68385, n12_adj_5611, 
        n55388, n6_adj_5612, n61204, n10_adj_5613, n61144, n61165, 
        n10_adj_5614, n56728, n25700, n26181, n25604, n1720, n25683, 
        n61248, n6_adj_5615, n55761, n54, n61424, n52, n60982, 
        n53, n51, n48, n50_adj_5616, n60976, n1655, n56308, n49, 
        n60, n61316, n55, n21_adj_5617, n56531, n60954, n12_adj_5618, 
        n56739, n72107, n26289, n26293, n12_adj_5619, n15_adj_5620, 
        n26323, n6_adj_5621, n56006, n61400, n61015, n1191, n12_adj_5622, 
        n8_adj_5623, n6_adj_5624, n55525, n6_adj_5625, n60912, n14_adj_5626, 
        n61239, n25458, n16_adj_5627, n55572, n13_adj_5628, n27721, 
        n65411, n18_adj_5629, n26038, n62886, n65412, n61394, n60799, 
        n65410, n18_adj_5631, n61406, n61242, n6_adj_5632, n20_adj_5633, 
        n26609, n61397, n15_adj_5634, n26308, n13_adj_5635, n26136, 
        n10_adj_5636, n12_adj_5637, n25528, n61279, n14_adj_5638, 
        n60874, n61082, n60921, n61264, n61446, n62942, n26457, 
        n14_adj_5639, n10_adj_5640, n61403, n61319, n10_adj_5641, 
        n1180, n61003, n61236, n60877, n63014, n61449, n10_adj_5642, 
        n63376, n60782, n63283, n26691, n28_c, n71957, n31_adj_5643, 
        n22_adj_5644, n30, n34_adj_5645, n15_adj_5646, n55595, n6_adj_5647, 
        n60796, n10_adj_5649, n61153, n14_adj_5650, n12_adj_5651, 
        n60806, n63420, n71951, n14_adj_5652, n12_adj_5654, n72098, 
        n71900, n19_adj_5655, n71945, n65414, n65415, n65413, n22_adj_5657, 
        n63172, n16_adj_5658, n61409, n17_adj_5659, n14_adj_5660, 
        n63189, n72101, n12_adj_5661, n56553, n14_adj_5662, n13_adj_5663, 
        n72095, n6_adj_5664, n8_adj_5665, n10_adj_5666, n11_adj_5667, 
        n25614, n9_adj_5668, n71933, n64955, n27719, n65405, n65406, 
        n65404, n71927, n63317, n71921, n61116, n72089, n72083, 
        n61070, n61036, n61092, n61055, Kp_23__N_748, n64947, n72077, 
        n26_adj_5669, n24, n55550, n72071, n71897, n63255, n30_adj_5670, 
        n65433, n56748, n28_adj_5671, n71873, n71867, n64725, n64727, 
        n72065, n29_c, n65181, n64735, n64741, n64747, n64753, 
        n64759, n64679, n63040, n7_adj_5672, n10_adj_5673;
    
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_13  (.CI(n54525), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n54526));
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[6] [4]), .I3(GND_net), .O(n64693));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n59876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2), .S(n60534));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5297), .S(n60533));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n29193));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n10), .I3(n61254), .O(n25746));   // verilog/coms.v(80[16:43])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(\data_in_frame[6] [4]), .I1(n16), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n18));   // verilog/coms.v(81[16:27])
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5298), .S(n60532));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27414), 
            .D(n4939[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5299), .S(n60531));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5300), .S(n28930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5301), .S(n60530));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5302), .S(n60474));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5303), .S(n60529));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5304), .S(n60528));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5305), .S(n60527));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5306), .S(n60526));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5307), .S(n60525));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27414), 
            .D(n4939[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_12_lut  (.I0(n68360), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n54524), .O(n27778)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27414), 
            .D(n4939[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27414), 
            .D(n4939[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27414), 
            .D(n4939[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5308), .S(n60524));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut (.I0(n25598), .I1(n60855), .I2(n61415), .I3(n26126), 
            .O(n17_c));   // verilog/coms.v(81[16:27])
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5309), .S(n60523));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5310), .S(n60522));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14138_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n29999));
    defparam i14138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5311), .S(n60476));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5312), .S(n60521));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5313), .S(n60520));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14141_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n30002));
    defparam i14141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27414), 
            .D(n4939[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_12  (.CI(n54524), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n54525));
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27414), 
            .D(n4939[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5314), .S(n60519));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27414), 
            .D(n4939[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27414), 
            .D(n4939[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14144_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n30005));
    defparam i14144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27414), 
            .D(n4939[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27414), 
            .D(n4939[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27414), 
            .D(n4939[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27414), 
            .D(n4939[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5315), .S(n60646));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_11_lut  (.I0(n68363), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n54523), .O(n27776)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_11  (.CI(n54523), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n54524));
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5316), .S(n60645));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14147_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n30008));
    defparam i14147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5317), .S(n60644));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29613));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14150_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n30011));
    defparam i14150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5318), .S(n60643));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[4] [1]), .I3(n60890), .O(n10_adj_5319));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5320), .S(n60642));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14153_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n30014));
    defparam i14153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14156_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n30017));
    defparam i14156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5321), .S(n60658));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14159_3_lut_4_lut (.I0(n8_c), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n30020));
    defparam i14159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29610));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5322), .S(n60641));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5323), .S(n60518));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i48065_4_lut (.I0(n56705), .I1(Kp_23__N_974), .I2(\data_in_frame[8] [0]), 
            .I3(\data_in_frame[8][6] ), .O(n65144));
    defparam i48065_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n21), .I1(n17), .I2(control_mode[0]), .I3(control_mode[1]), 
            .O(n22));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i48144_4_lut (.I0(n26220), .I1(n26250), .I2(n56127), .I3(n26089), 
            .O(n65225));
    defparam i48144_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(n25718), .I1(n26621), .I2(\data_in_frame[8][2] ), 
            .I3(GND_net), .O(n4_c));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5325), .S(n60517));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5326), .S(n60516));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13678_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29539));
    defparam i13678_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5328), .S(n60515));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5329), .S(n60514));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5330), .S(n60513));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5331), .S(n60512));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13681_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n29542));
    defparam i13681_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13684_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n29545));
    defparam i13684_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5332), .S(n60511));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5333), .S(n60510));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5334), .S(n60509));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5335), .S(n60508));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5336), .S(n60507));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5337), .S(n60506));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5338), .S(n60505));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5339), .S(n60504));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5340), .S(n60503));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5341), .S(n60502));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5342), .S(n60501));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5343), .S(n60500));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5344), .S(n60499));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5345), .S(n60640));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5346), .S(n60639));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29607));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5347), .S(n60638));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5348), .S(n60498));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5349), .S(n60497));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5350), .S(n60496));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5351), .S(n60495));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5352), .S(n60494));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5353), .S(n60493));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5354), .S(n60492));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut (.I0(n56707), .I1(n17_c), .I2(\data_in_frame[7] [7]), 
            .I3(n18), .O(n18_adj_5355));
    defparam i2_4_lut.LUT_INIT = 16'h4812;
    SB_DFFE data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29604));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5356), .S(n60637));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5357), .S(n60491));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5358), .S(n60490));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13688_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29549));
    defparam i13688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut (.I0(n26077), .I1(n71572), .I2(n25647), .I3(n7_c), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 select_787_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5360), .S(n60489));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29601));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1087 (.I0(\data_in_frame[8][3] ), .I1(Kp_23__N_869), 
            .I2(\data_in_frame[6] [2]), .I3(n25718), .O(n26220));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i48166_4_lut (.I0(n65225), .I1(n25732), .I2(n65144), .I3(n4_c), 
            .O(n65247));
    defparam i48166_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13691_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29552));
    defparam i13691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13694_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29555));
    defparam i13694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_10_lut  (.I0(n68364), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n54522), .O(n27774)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_10  (.CI(n54522), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n54523));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_9_lut  (.I0(n68365), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n54521), .O(n27772)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5361), .S(n60636));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29598));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5362), .S(n60635));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29595));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5363), .S(n60634));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29592));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5364), .S(n60633));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29589));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2881), .D(n8_adj_5365), .S(n60632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29586));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13697_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29558));
    defparam i13697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5366), .S(n60631));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29583));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5367), .S(n60630));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n29196));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_9  (.CI(n54521), .I0(n28031), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n54522));
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5368), .S(n60629));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29579));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5369), .S(n60628));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5370), .S(n60488));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29576));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5371), .S(n60627));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29573));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5372), .S(n60626));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29570));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5373), .S(n60625));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27414), 
            .D(n4939[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5374), .S(n60542));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5375), .S(n60487));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5376), .S(n60486));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29567));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5377), .S(n60485));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5378), .S(n60484));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5379), .S(n60483));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5380), .S(n60482));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5381), .S(n60481));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5382), .S(n60480));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5383), .S(n60479));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13700_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60740), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29561));
    defparam i13700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23236_3_lut_4_lut (.I0(n37468), .I1(control_mode[0]), .I2(control_update), 
            .I3(control_mode[1]), .O(n27465));   // verilog/coms.v(130[12] 305[6])
    defparam i23236_3_lut_4_lut.LUT_INIT = 16'hb0f0;
    SB_LUT4 select_787_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29564));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i15_4_lut (.I0(n17_adj_5385), .I1(n65247), .I2(n26), .I3(n18_adj_5355), 
            .O(n25249));
    defparam i15_4_lut.LUT_INIT = 16'h2000;
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5386), .S(n60478));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5387), .S(n60477));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [3]), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2881), .D(n3), .S(n60693));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5389), .S(n60690));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5390), .S(n60689));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5392), .S(n60688));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_8_lut  (.I0(n68366), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n54520), .O(n27770)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5393), .S(n60687));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_8  (.CI(n54520), .I0(n28031), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n54521));
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5394), .S(n60680));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5395), .S(n60694));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27414), 
            .D(n4939[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_7_lut  (.I0(n68367), .I1(n28031), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n54519), .O(n27768)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_7  (.CI(n54519), .I0(n28031), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n54520));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_6_lut  (.I0(n68369), .I1(n28031), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n54518), .O(n27766)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27414), 
            .D(n4939[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5396), .S(n60683));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5397), .S(n60691));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5398), .S(n60682));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_6  (.CI(n54518), .I0(n28031), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n54519));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_5_lut  (.I0(n68375), .I1(n28031), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n54517), .O(n27764)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_5  (.CI(n54517), .I0(n28031), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n54518));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_4_lut  (.I0(n68377), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n54516), .O(n27762)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_4  (.CI(n54516), .I0(n28031), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n54517));
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5400), .S(n60681));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5401), .S(n60624));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_3_lut  (.I0(n68380), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n54515), .O(n27760)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_3  (.CI(n54515), .I0(n28031), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n54516));
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5402), .S(n60685));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5403), .S(n60686));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5404), .S(n60679));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54931 (.I0(byte_transmit_counter[3]), 
            .I1(n70567), .I2(n68462), .I3(byte_transmit_counter[4]), .O(n72059));
    defparam byte_transmit_counter_3__bdd_4_lut_54931.LUT_INIT = 16'he4aa;
    SB_LUT4 n72059_bdd_4_lut (.I0(n72059), .I1(n71954), .I2(n7_adj_5405), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n72059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5406), .S(n60623));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n54515));
    SB_LUT4 i1_2_lut (.I0(n25647), .I1(n25732), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14114_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29975));
    defparam i14114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5408), .S(n60692));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14117_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29978));
    defparam i14117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1088 (.I0(\data_in_frame[16] [2]), .I1(n61335), 
            .I2(n56563), .I3(Kp_23__N_1271), .O(n61439));
    defparam i3_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_54926 (.I0(byte_transmit_counter[3]), 
            .I1(n70513), .I2(n68444), .I3(byte_transmit_counter[4]), .O(n72047));
    defparam byte_transmit_counter_3__bdd_4_lut_54926.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2881), .D(n3_adj_5409), .S(n60684));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2075), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29561));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n72047_bdd_4_lut (.I0(n72047), .I1(n71936), .I2(n65337), .I3(byte_transmit_counter[4]), 
            .O(tx_data[4]));
    defparam n72047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14120_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29981));
    defparam i14120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14123_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29984));
    defparam i14123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1089 (.I0(n61310), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[21] [0]), .I3(n61439), .O(n10_adj_5410));
    defparam i4_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[6] [7]), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'ha088;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27414), 
            .D(n4939[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2881), .D(n1_c), .S(n60673));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14126_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29987));
    defparam i14126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14129_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29990));
    defparam i14129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2881), .D(n1_adj_5412), .S(n60672));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(n60785), .I1(n10_adj_5410), .I2(\data_in_frame[20] [6]), 
            .I3(GND_net), .O(n55989));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14132_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29993));
    defparam i14132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14135_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29996));
    defparam i14135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i53620_4_lut (.I0(n71960), .I1(n72134), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n70710));
    defparam i53620_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i48223_3_lut (.I0(n71870), .I1(n70710), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i48223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_789_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1091 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n60730));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1091.LUT_INIT = 16'hfefe;
    SB_LUT4 select_789_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[7]), 
            .I3(GND_net), .O(n1_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFFE data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29558));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2881), .D(n1_adj_5415), .S(n60671));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2881), .D(n1_adj_5416), .S(n60670));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), 
            .C(clk16MHz), .E(n2881), .D(n1_adj_5417), .S(n60669));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), 
            .C(clk16MHz), .E(n2881), .D(n1_adj_5418), .S(n60668));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54921 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n72041));
    defparam byte_transmit_counter_0__bdd_4_lut_54921.LUT_INIT = 16'he4aa;
    SB_LUT4 i5359_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1958), 
            .I2(n62539), .I3(n4452), .O(n20871));   // verilog/coms.v(148[4] 304[11])
    defparam i5359_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1092 (.I0(n20871), .I1(n1958), .I2(n22473), .I3(n64994), 
            .O(n26846));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1092.LUT_INIT = 16'hbbba;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2067));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), 
            .C(clk16MHz), .E(n2881), .D(n1_adj_5414), .S(n60674));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1093 (.I0(Kp_23__N_1080), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n64711));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n72396), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n26843), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29555));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5419), .S(n60543));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2055), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2056), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20876), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n59808), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2067), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n26846), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i47918_4_lut (.I0(n1958), .I1(n1961), .I2(n3303), .I3(n1964), 
            .O(n64990));   // verilog/coms.v(139[4] 141[7])
    defparam i47918_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1094 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1961), 
            .I2(n64990), .I3(n62727), .O(n59808));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1094.LUT_INIT = 16'hb3a0;
    SB_LUT4 i5364_4_lut (.I0(n1962), .I1(\FRAME_MATCHER.state[3] ), .I2(n1964), 
            .I3(n25260), .O(n20876));   // verilog/coms.v(148[4] 304[11])
    defparam i5364_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2056));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2055));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_787_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[6]), 
            .I3(GND_net), .O(n1_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i23434_4_lut (.I0(n5), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i23434_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i54473_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[8] [1]), .I2(n28096), 
            .I3(GND_net), .O(n60128));   // verilog/coms.v(94[13:20])
    defparam i54473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\FRAME_MATCHER.i[4] ), .I1(n25281), .I2(GND_net), 
            .I3(GND_net), .O(n25150));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1]_c [0]), .I3(\data_in_frame[3] [2]), .O(n60833));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[5]), 
            .I3(GND_net), .O(n1_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i23435_4_lut (.I0(n8), .I1(\FRAME_MATCHER.i [31]), .I2(n25150), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i23435_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n22473));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_789_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i3_2_lut (.I0(n25260), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27402));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1097 (.I0(n4452), .I1(n27402), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22473), .O(n63171));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1097.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1098 (.I0(n25265), .I1(n1964), .I2(n1962), .I3(n63171), 
            .O(n26843));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1098.LUT_INIT = 16'hbaaa;
    SB_LUT4 select_789_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_2_lut_adj_1099 (.I0(\data_in[3] [3]), .I1(\data_in[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_c));
    defparam i2_2_lut_adj_1099.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1100 (.I0(\data_in[3] [6]), .I1(\data_in[2] [1]), 
            .I2(n6_c), .I3(\data_in[3] [5]), .O(n6_adj_5421));   // verilog/coms.v(142[7:80])
    defparam i1_4_lut_adj_1100.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_1101 (.I0(\data_in[2] [3]), .I1(\data_in[3] [1]), 
            .I2(\data_in[0] [2]), .I3(n6_adj_5421), .O(n25313));   // verilog/coms.v(142[7:80])
    defparam i4_4_lut_adj_1101.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), .I2(n25313), 
            .I3(\data_in[0] [5]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1102 (.I0(n25163), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19));
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1103 (.I0(n7_c), .I1(n24870), .I2(n64711), .I3(n60985), 
            .O(n60987));
    defparam i1_4_lut_adj_1103.LUT_INIT = 16'h9669;
    SB_LUT4 i48108_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[1] [3]), .I2(\data_in[0] [1]), 
            .I3(\data_in[3] [2]), .O(n65189));
    defparam i48108_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n65189), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n1958));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1104 (.I0(\data_in[2] [4]), .I1(n25313), .I2(\data_in[1] [5]), 
            .I3(n25394), .O(n18_adj_5422));
    defparam i7_4_lut_adj_1104.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(\data_in[0] [6]), .I1(n18_adj_5422), .I2(\data_in[3] [0]), 
            .I3(n25325), .O(n20_adj_5423));
    defparam i9_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_c));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1105 (.I0(n15_c), .I1(n20_adj_5423), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1961));
    defparam i10_4_lut_adj_1105.LUT_INIT = 16'hfeff;
    SB_LUT4 i23265_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n39028));
    defparam i23265_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5424));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1107 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_5425));
    defparam i1_4_lut_adj_1107.LUT_INIT = 16'ha8a0;
    SB_LUT4 i23763_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter_c[7]), 
            .I2(n4_adj_5425), .I3(n4_adj_5424), .O(n39534));
    defparam i23763_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n32327));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'heeee;
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5411), .S(n31));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), .I2(\data_in[3] [2]), 
            .I3(\data_in[0] [5]), .O(n16_adj_5426));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1109 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5427));
    defparam i7_4_lut_adj_1109.LUT_INIT = 16'hfffd;
    SB_DFFE data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29552));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i9_4_lut_adj_1110 (.I0(n17_adj_5427), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5426), .I3(\data_in[2] [6]), .O(n25325));
    defparam i9_4_lut_adj_1110.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1111 (.I0(\data_in[0] [4]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [7]), .I3(\data_in[3] [4]), .O(n10_adj_5428));
    defparam i4_4_lut_adj_1111.LUT_INIT = 16'hdfff;
    SB_LUT4 i5_3_lut_adj_1112 (.I0(\data_in[1] [1]), .I1(n10_adj_5428), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n25394));
    defparam i5_3_lut_adj_1112.LUT_INIT = 16'hefef;
    SB_LUT4 select_787_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_adj_1113 (.I0(\data_in[0] [3]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [0]), .I3(GND_net), .O(n14));
    defparam i5_3_lut_adj_1113.LUT_INIT = 16'hdfdf;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5407), .S(n60622));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1114 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(n25394), .I3(\data_in[1] [5]), .O(n15_adj_5429));
    defparam i6_4_lut_adj_1114.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1115 (.I0(n15_adj_5429), .I1(\data_in[1] [0]), 
            .I2(n14), .I3(\data_in[2] [2]), .O(n25163));
    defparam i8_4_lut_adj_1115.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n25163), .O(n16_adj_5430));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(n25325), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_5431));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1118 (.I0(n17_adj_5431), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5430), .I3(\data_in[3] [1]), .O(n1964));
    defparam i9_4_lut_adj_1118.LUT_INIT = 16'hfbff;
    SB_LUT4 i366_2_lut (.I0(n1961), .I1(n1958), .I2(GND_net), .I3(GND_net), 
            .O(n1962));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1119 (.I0(n39534), .I1(n62533), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n39028), .O(n6_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1119.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(n32327), .I1(n6_adj_5432), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n72396));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'hefee;
    SB_LUT4 n72041_bdd_4_lut (.I0(n72041), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n72044));
    defparam n72041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1_c));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i13_2_lut (.I0(pwm_setpoint[15]), .I1(\pwm_counter[15] ), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_10));   // verilog/pwm.v(11[19:30])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29549));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1121 (.I0(n26178), .I1(n60987), .I2(n25732), 
            .I3(\data_in_frame[10] [6]), .O(n55997));
    defparam i1_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5399), .S(n60621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1122 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[7] [4]), 
            .I2(n60833), .I3(n6_adj_5434), .O(n61412));
    defparam i4_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[13] [2]), .I1(n55997), 
            .I2(GND_net), .I3(GND_net), .O(n60969));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i12_2_lut (.I0(\pwm_counter[16] ), .I1(pwm_setpoint[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(95[20:32])
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n29199));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5391), .S(n60620));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29545));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29542));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25501));
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29539));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i160 (.Q(\data_in_frame[19] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29536));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5388), .S(n29020));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29533));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5384), .S(n60619));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i158 (.Q(\data_in_frame[19] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29530));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i157 (.Q(\data_in_frame[19] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29527));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i156 (.Q(\data_in_frame[19] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29524));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29521));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1125 (.I0(\data_in_frame[11] [6]), .I1(n23700), 
            .I2(n25501), .I3(n26250), .O(n60979));
    defparam i3_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(n26123), .I1(n60855), .I2(Kp_23__N_878), 
            .I3(\data_in_frame[8][7] ), .O(n7_c));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(n56744), .I1(n56678), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n56555));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1126 (.I0(\data_in_frame[12] [7]), .I1(n60896), 
            .I2(\data_in_frame[15] [2]), .I3(n25825), .O(n61313));
    defparam i3_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n60858));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[4] [2]), .O(n37));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1128 (.I0(n26123), .I1(n60855), .I2(Kp_23__N_878), 
            .I3(n71572), .O(n55521));
    defparam i1_2_lut_4_lut_adj_1128.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(control_mode_c[5]), .I1(\control_mode[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n48532));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1130 (.I0(control_mode_c[3]), .I1(\control_mode[2] ), 
            .I2(\control_mode[4] ), .I3(GND_net), .O(n17));
    defparam i1_3_lut_adj_1130.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(n17), .I1(n21), .I2(GND_net), .I3(GND_net), 
            .O(n37468));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(157[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(157[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1132 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1132.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut_adj_1133 (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(157[7:23])
    defparam i13_2_lut_adj_1133.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(157[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(157[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n25281));   // verilog/coms.v(157[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23436_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25281), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i23436_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2075));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1134 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [1]), 
            .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1134.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[1]_c [3]), .I1(n60858), .I2(n61326), 
            .I3(n61012), .O(n25718));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1135 (.I0(n61313), .I1(n60969), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[12] [6]), .O(n56505));
    defparam i1_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1136 (.I0(n56535), .I1(n56678), .I2(\data_in_frame[15] [5]), 
            .I3(GND_net), .O(n25564));
    defparam i1_3_lut_adj_1136.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_223_i3_4_lut (.I0(n56675), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n60816), .I3(\data_out_frame[25] [6]), .O(n3_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_223_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i51785_2_lut (.I0(n72044), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68444));
    defparam i51785_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i53423_3_lut (.I0(n72080), .I1(n71978), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70513));
    defparam i53423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1137 (.I0(\data_in_frame[15] [3]), .I1(n56505), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n62519));
    defparam i1_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_222_i3_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5435), .I3(n60816), 
            .O(n3_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_222_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60825));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61030));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26057));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n29520));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[8][7] ), .I1(\data_in_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61433));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29517));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1142 (.I0(n26120), .I1(n26447), .I2(GND_net), 
            .I3(GND_net), .O(n61329));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1143 (.I0(\data_in_frame[4] [4]), .I1(n25598), 
            .I2(n26154), .I3(GND_net), .O(n26123));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_in_frame[6] [7]), .I1(n25591), 
            .I2(GND_net), .I3(GND_net), .O(n26451));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_in_frame[8] [1]), .I1(n56705), 
            .I2(GND_net), .I3(GND_net), .O(n60841));
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h9999;
    SB_DFFE data_in_frame_0___i153 (.Q(\data_in_frame[19] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29514));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29513));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1146 (.I0(\data_in_frame[13] [7]), .I1(n55574), 
            .I2(GND_net), .I3(GND_net), .O(n61129));
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1147 (.I0(n61329), .I1(n60871), .I2(Kp_23__N_878), 
            .I3(n61433), .O(n10));
    defparam i4_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[1]_c [3]), .I1(n60858), .I2(n56614), 
            .I3(n61125), .O(n56705));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61104));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1149 (.I0(n60837), .I1(Kp_23__N_772), .I2(\data_in_frame[1] [4]), 
            .I3(GND_net), .O(n61261));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n59920));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51721_2_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n68446));
    defparam i51721_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(n26274), .I1(n56634), .I2(GND_net), 
            .I3(GND_net), .O(n56529));
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25687));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i48264_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65354));
    defparam i48264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48265_4_lut (.I0(n65354), .I1(n68446), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n65355));
    defparam i48265_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i48263_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65353));
    defparam i48263_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n59922));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n29205));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i52193_2_lut (.I0(n72140), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68462));
    defparam i52193_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1152 (.I0(n61122), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[12] [1]), .O(n64917));
    defparam i1_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i53477_3_lut (.I0(n72188), .I1(n71876), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70567));
    defparam i53477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1153 (.I0(n26447), .I1(n64873), .I2(n25591), 
            .I3(n25987), .O(n63380));   // verilog/coms.v(88[17:70])
    defparam i1_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i54482_2_lut (.I0(n63380), .I1(\data_in_frame[7] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n71572));   // verilog/coms.v(99[12:25])
    defparam i54482_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1154 (.I0(n26451), .I1(n61329), .I2(n61030), 
            .I3(\data_in_frame[4] [5]), .O(n26077));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29501));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29498));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1155 (.I0(n61458), .I1(n64921), .I2(n64917), 
            .I3(n61361), .O(n64925));
    defparam i1_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29495));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1156 (.I0(n63380), .I1(n26057), .I2(\data_in_frame[10] [7]), 
            .I3(n60896), .O(n5_adj_5436));
    defparam i1_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29492));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1157 (.I0(n62519), .I1(n56555), .I2(\data_in_frame[19] [6]), 
            .I3(GND_net), .O(n56559));
    defparam i1_2_lut_3_lut_adj_1157.LUT_INIT = 16'h9696;
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29489));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29486));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29483));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29480));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29477));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1158 (.I0(n62519), .I1(n56555), .I2(n62964), 
            .I3(GND_net), .O(n26599));
    defparam i1_2_lut_3_lut_adj_1158.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n29208));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29473));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14090_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29951));
    defparam i14090_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5438), .S(n60618));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n29211));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n29214));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n29217));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n29220));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29466));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29463));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29460));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1159 (.I0(\data_in_frame[11] [2]), .I1(n5_adj_5436), 
            .I2(\data_in_frame[7] [3]), .I3(\data_in_frame[8][2] ), .O(n6_adj_5439));
    defparam i1_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29459));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29456));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5440), .S(n60617));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29451));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29448));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n70717), .I2(n68429), .I3(byte_transmit_counter[4]), .O(n72209));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFFE data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29445));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29442));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29439));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29436));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29433));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14093_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29954));
    defparam i14093_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29430));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29427));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29424));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5441), .S(n60616));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29421));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29418));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29415));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29412));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29409));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29406));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29403));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29400));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29397));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1160 (.I0(n25658), .I1(n61048), .I2(n60927), 
            .I3(n64925), .O(n64931));
    defparam i1_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29394));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n72209_bdd_4_lut (.I0(n72209), .I1(n71924), .I2(n7_adj_5442), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n72209_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n29224));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n29229));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n29232));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n29240));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1161 (.I0(n23704), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[11] [1]), .I3(n6_adj_5439), .O(n63425));
    defparam i4_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55001 (.I0(byte_transmit_counter[1]), 
            .I1(n65623), .I2(n65624), .I3(byte_transmit_counter[2]), .O(n72005));
    defparam byte_transmit_counter_1__bdd_4_lut_55001.LUT_INIT = 16'he4aa;
    SB_LUT4 n72005_bdd_4_lut (.I0(n72005), .I1(n65309), .I2(n65308), .I3(byte_transmit_counter[2]), 
            .O(n72008));
    defparam n72005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n29243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27414), 
            .D(n4939[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i14096_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29957));
    defparam i14096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27414), 
            .D(n4939[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27414), 
            .D(n4939[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27414), 
            .D(n4939[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27414), 
            .D(n4939[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27414), 
            .D(n4939[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27414), 
            .D(n4939[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n29246));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n29249));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1162 (.I0(n61436), .I1(n63425), .I2(n64933), 
            .I3(n64931), .O(n64939));
    defparam i1_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55046 (.I0(byte_transmit_counter[3]), 
            .I1(n70699), .I2(n68453), .I3(byte_transmit_counter[4]), .O(n72197));
    defparam byte_transmit_counter_3__bdd_4_lut_55046.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n29252));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n29255));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n29258));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n29261));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n29264));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n29267));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
           .D(n29270));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
           .D(n29273));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
           .D(n29276));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1163 (.I0(n64939), .I1(n56529), .I2(n60841), 
            .I3(n61141), .O(n24953));
    defparam i1_4_lut_adj_1163.LUT_INIT = 16'h9669;
    SB_LUT4 i14099_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29960));
    defparam i14099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14102_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29963));
    defparam i14102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14105_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29966));
    defparam i14105_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14108_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29969));
    defparam i14108_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8][1] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5443), .S(n60615));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1271));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1164 (.I0(n55540), .I1(n26077), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n55580));
    defparam i2_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n64961));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1166 (.I0(n55580), .I1(n60903), .I2(n25817), 
            .I3(n64961), .O(n56075));
    defparam i1_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(\data_in_frame[18] [3]), .I1(n56075), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5444));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1168 (.I0(n56684), .I1(n55705), .I2(n61104), 
            .I3(n6_adj_5444), .O(n55503));
    defparam i4_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1169 (.I0(n55503), .I1(\data_in_frame[20] [5]), 
            .I2(\data_in_frame[20] [6]), .I3(GND_net), .O(n60960));
    defparam i2_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1170 (.I0(\data_in_frame[4] [4]), .I1(n60880), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[1] [7]), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1171 (.I0(Kp_23__N_878), .I1(n60932), .I2(\data_in_frame[6] [4]), 
            .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(GND_net), .I3(GND_net), .O(n61048));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n61201), .I1(n61018), .I2(n61295), 
            .I3(n60871), .O(n14_adj_5445));
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[9] [0]), .I1(n60828), .I2(n60932), 
            .I3(\data_in_frame[5] [0]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1174 (.I0(n13), .I1(n10_adj_5446), .I2(n61455), 
            .I3(n14_adj_5445), .O(n12));
    defparam i5_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1175 (.I0(n61412), .I1(n12), .I2(\data_in_frame[14] [2]), 
            .I3(n61361), .O(n56563));
    defparam i6_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1176 (.I0(n61295), .I1(\data_in_frame[11] [5]), 
            .I2(n55521), .I3(\data_in_frame[13] [7]), .O(n14_adj_5447));
    defparam i6_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1177 (.I0(\data_in_frame[14] [1]), .I1(n14_adj_5447), 
            .I2(n10_adj_5448), .I3(n25556), .O(n56684));
    defparam i7_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54912 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[1]), .O(n71987));
    defparam byte_transmit_counter_0__bdd_4_lut_54912.LUT_INIT = 16'he4aa;
    SB_LUT4 i14111_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29972));
    defparam i14111_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_in_frame[16] [3]), .I1(n25950), 
            .I2(GND_net), .I3(GND_net), .O(n60963));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i54472_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[8] [0]), .I2(n28096), 
            .I3(GND_net), .O(n60118));   // verilog/coms.v(94[13:20])
    defparam i54472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(n56684), .I1(n56563), .I2(GND_net), 
            .I3(GND_net), .O(n56561));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(\data_in_frame[10] [5]), .I1(n25732), 
            .I2(n26220), .I3(GND_net), .O(n61107));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5449));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1182 (.I0(\data_in_frame[20] [2]), .I1(n60822), 
            .I2(Kp_23__N_1389), .I3(\data_in_frame[18] [0]), .O(n10_adj_5450));
    defparam i4_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1183 (.I0(n56678), .I1(n10_adj_5450), .I2(\data_in_frame[13] [4]), 
            .I3(GND_net), .O(n61178));
    defparam i5_3_lut_adj_1183.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(n55503), .I1(n60785), .I2(GND_net), 
            .I3(GND_net), .O(n64883));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1185 (.I0(Kp_23__N_1518), .I1(n61388), .I2(n61174), 
            .I3(n64883), .O(n61367));
    defparam i1_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 n72197_bdd_4_lut (.I0(n72197), .I1(n72008), .I2(n7_adj_5451), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n72197_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n71987_bdd_4_lut (.I0(n71987), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[1]), 
            .O(n71990));
    defparam n71987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1186 (.I0(n25647), .I1(n61107), .I2(n26178), 
            .I3(n6_adj_5449), .O(n61282));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1187 (.I0(\data_in_frame[20] [3]), .I1(n55503), 
            .I2(\data_in_frame[20] [4]), .I3(GND_net), .O(n5_adj_5452));
    defparam i1_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5454), .S(n60657));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5455), .S(n60656));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5456), .S(n60655));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5457), .S(n60654));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5458), .S(n60653));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5459), .S(n60652));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5460), .S(n60651));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5461), .S(n60650));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5462), .S(n60649));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5463), .S(n60648));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5464), .S(n60647));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8][2] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5465), .S(n60614));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8][3] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5466), .S(n60613));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8][4] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5467), .S(n60612));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8][5] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5468), .S(n60611));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8][6] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5469), .S(n60610));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8][7] ), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5470), .S(n60609));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5471), .S(n60608));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5472), .S(n60607));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5473), .S(n60606));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5474), .S(n60605));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5475), .S(n60604));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5476), .S(n60603));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5477), .S(n29002));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5478), .S(n60602));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5479), .S(n60601));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5480), .S(n60600));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5481), .S(n60599));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5482), .S(n60598));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5483), .S(n60597));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5484), .S(n60596));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5485), .S(n60595));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5486), .S(n60594));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5487), .S(n60593));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5488), .S(n60592));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5489), .S(n60591));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5490), .S(n60590));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5491), .S(n60589));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5492), .S(n60588));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5493), .S(n60587));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5494), .S(n60586));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5495), .S(n60585));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5496), .S(n60584));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5497), .S(n60583));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5498), .S(n60582));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5499), .S(n60581));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n29309));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5500), .S(n60580));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n29308));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5501), .S(n60579));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n29307));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5502), .S(n60578));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n29306));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5503), .S(n60577));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n29305));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5504), .S(n60576));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n29304));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5505), .S(n60575));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n29303));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5506), .S(n60574));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n29302));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5507), .S(n60573));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n29301));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5508), .S(n60572));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n29300));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5509), .S(n60571));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n29299));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5510), .S(n60570));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n29298));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5511), .S(n60569));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n29297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5512), .S(n60568));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n29296));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5513), .S(n60567));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n29295));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5514), .S(n60566));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n29294));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5515), .S(n60565));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n29293));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5516), .S(n60564));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n29292));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5517), .S(n60563));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n29291));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5518), .S(n60562));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n29290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5519), .S(n60561));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n29289));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5520), .S(n60560));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n29288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5521), .S(n60559));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n29287));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5522), .S(n60558));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n29286));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5523), .S(n60557));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n29285));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5524), .S(n60556));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n29284));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5525), .S(n60555));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n29283));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n29282));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5526), .S(n60554));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n29281));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n29280));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n29279));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5527), .S(n60553));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5528), .S(n60475));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5529), .S(n60552));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5530), .S(n60551));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5531), .S(n60550));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5532), .S(n60549));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5533), .S(n60548));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5534), .S(n60547));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5535), .S(n60546));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5536), .S(n60545));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i51625_2_lut (.I0(\data_out_frame[9] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n68321));
    defparam i51625_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29236));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5537), .S(n60544));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5538), .S(n60541));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5539), .S(n60540));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5540), .S(n60539));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n72191));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i9_3_lut (.I0(\data_out_frame[10] [0]), 
            .I1(\data_out_frame[11] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1188 (.I0(\data_in_frame[15] [3]), .I1(n61282), 
            .I2(n60969), .I3(\data_in_frame[13] [1]), .O(n56744));
    defparam i1_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i18870_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n12_adj_5541));   // verilog/coms.v(105[12:33])
    defparam i18870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i11_3_lut (.I0(\data_out_frame[12] [0]), 
            .I1(\data_out_frame[13] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51626_2_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n68319));
    defparam i51626_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51786_2_lut (.I0(\data_out_frame[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n68320));
    defparam i51786_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5542));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32773_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n4_adj_5543));   // verilog/coms.v(105[12:33])
    defparam i32773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n72191_bdd_4_lut (.I0(n72191), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n72194));
    defparam n72191_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n61323));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i48312_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65402));
    defparam i48312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48313_4_lut (.I0(n65402), .I1(n27827), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][5] ), .O(n65403));
    defparam i48313_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i48311_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65401));
    defparam i48311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51797_2_lut (.I0(n72104), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68434));
    defparam i51797_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i47942_4_lut (.I0(n5_adj_5452), .I1(n55137), .I2(n61344), 
            .I3(\data_in_frame[22] [5]), .O(n65016));
    defparam i47942_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i2_3_lut_adj_1190 (.I0(n60947), .I1(n61298), .I2(\data_in_frame[23] [4]), 
            .I3(GND_net), .O(n62580));
    defparam i2_3_lut_adj_1190.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1191 (.I0(\data_in_frame[20] [5]), .I1(n61174), 
            .I2(\data_in_frame[22] [6]), .I3(\data_in_frame[20] [4]), .O(n63286));
    defparam i3_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1192 (.I0(n62654), .I1(\data_in_frame[20] [3]), 
            .I2(\data_in_frame[22] [4]), .I3(n6_adj_5544), .O(n63297));
    defparam i4_4_lut_adj_1192.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1193 (.I0(n63297), .I1(n63286), .I2(n62580), 
            .I3(n65016), .O(n64829));
    defparam i1_4_lut_adj_1193.LUT_INIT = 16'h0080;
    SB_LUT4 i1_3_lut_adj_1194 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[23] [3]), 
            .I2(n61298), .I3(GND_net), .O(n4_adj_5545));
    defparam i1_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1195 (.I0(\data_in_frame[21] [1]), .I1(n64829), 
            .I2(\data_in_frame[23] [2]), .I3(n55989), .O(n64831));
    defparam i1_4_lut_adj_1195.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5546));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1197 (.I0(n63036), .I1(n56596), .I2(n64831), 
            .I3(n4_adj_5545), .O(n64835));
    defparam i1_4_lut_adj_1197.LUT_INIT = 16'h8020;
    SB_LUT4 i4_4_lut_adj_1198 (.I0(\data_in_frame[22] [0]), .I1(n55682), 
            .I2(n56559), .I3(n6_adj_5546), .O(n62755));
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_DFFR \FRAME_MATCHER.i_2043__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n27733), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i53591_3_lut (.I0(n72110), .I1(n71990), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70681));
    defparam i53591_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2881), .D(n5_adj_5547), 
            .S(n28610));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1199 (.I0(n60979), .I1(\data_in_frame[14] [0]), 
            .I2(n25765), .I3(GND_net), .O(n61335));
    defparam i2_3_lut_adj_1199.LUT_INIT = 16'h9696;
    SB_LUT4 i14042_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[1]_c [0]), .O(n29903));
    defparam i14042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2881), .D(n26729), 
            .S(n28603));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1200 (.I0(n61344), .I1(\data_in_frame[20] [0]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[22] [2]), .O(n64903));
    defparam i1_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1201 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(n10_adj_5319), .I3(\data_in_frame[3] [6]), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1202 (.I0(\data_in_frame[23] [7]), .I1(n62755), 
            .I2(n60966), .I3(n64835), .O(n64839));
    defparam i1_4_lut_adj_1202.LUT_INIT = 16'h4800;
    SB_LUT4 i1_4_lut_adj_1203 (.I0(\data_in_frame[23] [5]), .I1(n64839), 
            .I2(n60947), .I3(n55692), .O(n64841));
    defparam i1_4_lut_adj_1203.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n25461), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[6] [3]), .O(n1244));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2881), .D(n1_adj_5549), .S(n28599));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[3] [7]), .O(n61326));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1205 (.I0(n26154), .I1(n60993), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[6] [5]), .O(n60932));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1206 (.I0(n26154), .I1(n60993), .I2(\data_in_frame[2] [0]), 
            .I3(Kp_23__N_872), .O(n6_adj_5550));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i14045_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29906));
    defparam i14045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5551));
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i3_4_lut_adj_1207 (.I0(\data_in_frame[21] [7]), .I1(n61285), 
            .I2(n60906), .I3(\data_in_frame[22] [1]), .O(n62556));
    defparam i3_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i23699_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n39467));
    defparam i23699_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i14048_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[1][2] ), .O(n29909));
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14051_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n29912));
    defparam i14051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1208 (.I0(n61355), .I1(n62822), .I2(\data_out_frame[10] [3]), 
            .I3(\data_out_frame[6] [1]), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55036 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n72185));
    defparam byte_transmit_counter_0__bdd_4_lut_55036.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1209 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2513 ), .I3(n60730), .O(n63143));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1209.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1210 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3483));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1210.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1211 (.I0(n161), .I1(n37935), .I2(n3483), 
            .I3(n39467), .O(n60700));
    defparam i2_3_lut_4_lut_adj_1211.LUT_INIT = 16'h8000;
    SB_LUT4 n72185_bdd_4_lut (.I0(n72185), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n72188));
    defparam n72185_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1212 (.I0(n161), .I1(n37935), .I2(reset), 
            .I3(n28031), .O(n60740));
    defparam i2_3_lut_4_lut_adj_1212.LUT_INIT = 16'hfff7;
    SB_LUT4 i13728_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n29589));
    defparam i13728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13731_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29592));
    defparam i13731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1213 (.I0(n60785), .I1(n26198), .I2(\data_in_frame[18] [1]), 
            .I3(\data_in_frame[20] [1]), .O(n64705));
    defparam i1_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i14054_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29915));
    defparam i14054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14057_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[1]_c [5]), .O(n29918));
    defparam i14057_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13734_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n29595));
    defparam i13734_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13737_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29598));
    defparam i13737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13740_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29601));
    defparam i13740_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13743_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29604));
    defparam i13743_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54867 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n71975));
    defparam byte_transmit_counter_0__bdd_4_lut_54867.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5552), .S(n60538));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13746_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29607));
    defparam i13746_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13749_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60740), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29610));
    defparam i13749_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14060_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[1][6] ), .O(n29921));
    defparam i14060_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14063_3_lut_4_lut (.I0(n8_adj_11), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29924));
    defparam i14063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n71975_bdd_4_lut (.I0(n71975), .I1(\data_out_frame[21] [4]), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n71978));
    defparam n71975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2881), .D(n1_adj_5413), .S(n60667));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1214 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [0]), 
            .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1214.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [7]), 
            .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1216 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1216.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_304_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_11));   // verilog/coms.v(157[7:23])
    defparam equal_304_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[1]_c [5]), .I1(\data_in_frame[1]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60837));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n61267));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1219 (.I0(n56555), .I1(Kp_23__N_1518), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n62899));
    defparam i1_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55031 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n72179));
    defparam byte_transmit_counter_0__bdd_4_lut_55031.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1220 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[5] [6]), .O(n64645));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1221 (.I0(n64645), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[2] [2]), .O(n64647));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1222 (.I0(n60890), .I1(n61267), .I2(n60858), 
            .I3(n61098), .O(n64657));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1223 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1958), .I3(n1961), .O(n25265));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1223.LUT_INIT = 16'h4000;
    SB_LUT4 n72179_bdd_4_lut (.I0(n72179), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n72182));
    defparam n72179_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1224 (.I0(n25591), .I1(n64647), .I2(n60861), 
            .I3(n60844), .O(n64659));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1225 (.I0(n64659), .I1(n25540), .I2(n64657), 
            .I3(GND_net), .O(n64665));   // verilog/coms.v(73[16:27])
    defparam i1_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1226 (.I0(n61224), .I1(n62899), .I2(n63034), 
            .I3(n64705), .O(n61388));
    defparam i1_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1227 (.I0(n26120), .I1(n60880), .I2(n64665), 
            .I3(n64663), .O(n64671));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1228 (.I0(n25987), .I1(n64685), .I2(n64671), 
            .I3(n25669), .O(n55544));   // verilog/coms.v(73[16:27])
    defparam i1_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1229 (.I0(n1958), .I1(n4452), .I2(n1961), 
            .I3(n1964), .O(n62539));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1229.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_1230 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[14][6] ), .I3(\data_in_frame[17] [1]), .O(n64783));
    defparam i1_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1231 (.I0(n61285), .I1(n56575), .I2(n64903), 
            .I3(n62519), .O(n64909));
    defparam i1_4_lut_adj_1231.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1958), .I1(n4452), .I2(n64994), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n62727));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_1232 (.I0(n64783), .I1(n60990), .I2(\data_in_frame[16] [3]), 
            .I3(\data_in_frame[13] [7]), .O(n64791));
    defparam i1_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1233 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[5] [3]), .I3(GND_net), .O(n64685));
    defparam i1_2_lut_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1234 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[7] [2]), .I3(\data_in_frame[5] [1]), .O(n63330));
    defparam i2_3_lut_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(\data_in_frame[8][6] ), .I1(\data_in_frame[11] [0]), 
            .I2(Kp_23__N_974), .I3(GND_net), .O(n26178));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1236 (.I0(n60883), .I1(n61323), .I2(n61104), 
            .I3(Kp_23__N_1389), .O(n64793));
    defparam i1_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55041 (.I0(byte_transmit_counter[3]), 
            .I1(n70681), .I2(n68434), .I3(byte_transmit_counter[4]), .O(n72167));
    defparam byte_transmit_counter_3__bdd_4_lut_55041.LUT_INIT = 16'he4aa;
    SB_LUT4 n72167_bdd_4_lut (.I0(n72167), .I1(n71930), .I2(n7_adj_5553), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n72167_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(n61335), .I1(n61313), .I2(n64793), 
            .I3(n64791), .O(n64799));
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55026 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(byte_transmit_counter[1]), 
            .O(n72161));
    defparam byte_transmit_counter_0__bdd_4_lut_55026.LUT_INIT = 16'he4aa;
    SB_LUT4 n72161_bdd_4_lut (.I0(n72161), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(byte_transmit_counter[1]), 
            .O(n65333));
    defparam n72161_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1238 (.I0(n61198), .I1(n56640), .I2(n64799), 
            .I3(n61102), .O(n64805));
    defparam i1_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5543), .I2(n5_adj_5542), .I3(byte_transmit_counter[2]), 
            .O(n72155));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n72155_bdd_4_lut (.I0(n72155), .I1(n68320), .I2(n68319), .I3(byte_transmit_counter[2]), 
            .O(n65337));
    defparam n72155_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1239 (.I0(n55511), .I1(n61185), .I2(n60973), 
            .I3(n64805), .O(n64811));
    defparam i1_4_lut_adj_1239.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_55006 (.I0(byte_transmit_counter[1]), 
            .I1(n11), .I2(n12_adj_5541), .I3(byte_transmit_counter[2]), 
            .O(n72149));
    defparam byte_transmit_counter_1__bdd_4_lut_55006.LUT_INIT = 16'he4aa;
    SB_LUT4 n72149_bdd_4_lut (.I0(n72149), .I1(n9), .I2(n68321), .I3(byte_transmit_counter[2]), 
            .O(n72152));
    defparam n72149_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1240 (.I0(n56561), .I1(n56744), .I2(n61381), 
            .I3(n64811), .O(n64817));
    defparam i1_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_55011 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n72143));
    defparam byte_transmit_counter_0__bdd_4_lut_55011.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1241 (.I0(n25564), .I1(n26599), .I2(n55970), 
            .I3(n64817), .O(Kp_23__N_1518));
    defparam i1_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 n72143_bdd_4_lut (.I0(n72143), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n72146));
    defparam n72143_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1242 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n10_adj_5554), .I3(n59688), .O(n61298));   // verilog/coms.v(81[16:27])
    defparam i5_3_lut_4_lut_adj_1242.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1243 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n60785));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1243.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1244 (.I0(n64909), .I1(n62556), .I2(n61367), 
            .I3(n64841), .O(n64845));
    defparam i1_4_lut_adj_1244.LUT_INIT = 16'h1200;
    SB_LUT4 i1_2_lut_3_lut_adj_1245 (.I0(n26220), .I1(n4_c), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n25825));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1245.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5453), .S(n60537));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1246 (.I0(n56575), .I1(n61178), .I2(\data_in_frame[19] [7]), 
            .I3(\data_in_frame[22] [3]), .O(n64881));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1247 (.I0(n56596), .I1(n61051), .I2(\data_in_frame[23] [1]), 
            .I3(GND_net), .O(n62406));
    defparam i1_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n59930));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13243_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n29104));   // verilog/coms.v(148[4] 304[11])
    defparam i13243_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13244_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n29105));   // verilog/coms.v(148[4] 304[11])
    defparam i13244_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5552));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13245_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [0]), 
            .I3(\Kp[0] ), .O(n29106));   // verilog/coms.v(148[4] 304[11])
    defparam i13245_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13246_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n29107));   // verilog/coms.v(148[4] 304[11])
    defparam i13246_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18876_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10]_c [0]), 
            .I3(PWMLimit[0]), .O(n29111));   // verilog/coms.v(148[4] 304[11])
    defparam i18876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13833_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][7] ), 
            .I3(PWMLimit[23]), .O(n29694));   // verilog/coms.v(148[4] 304[11])
    defparam i13833_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29629));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29632));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n29098));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n60118));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
           .D(n29680));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30065));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30062));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30059));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30056));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30053));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30050));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30047));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30044));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30041));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i54 (.Q(\data_in_frame[6] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30038));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30035));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30032));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30029));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30026));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i49 (.Q(\data_in_frame[6] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30023));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30020));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n30017));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n30014));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n30011));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30008));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30005));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30002));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29999));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29996));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29993));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13834_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][6] ), 
            .I3(PWMLimit[22]), .O(n29695));   // verilog/coms.v(148[4] 304[11])
    defparam i13834_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29990));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29984));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29981));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29978));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29975));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29972));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29966));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29963));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i28 (.Q(\data_in_frame[3] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29960));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29957));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29954));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i25 (.Q(\data_in_frame[3] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29951));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29948));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29945));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29942));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29936));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29933));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29930));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29924));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1]_c [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29918));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1][2] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29909));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29906));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1]_c [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29897));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26198));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29888));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29882));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n60128));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1249 (.I0(\data_in_frame[5] [4]), .I1(n60833), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n25540));
    defparam i1_3_lut_adj_1249.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8][2] ), .C(clk16MHz), 
           .D(n29127));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8][3] ), .C(clk16MHz), 
           .D(n29130));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8][4] ), .C(clk16MHz), 
           .D(n29133));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\data_in_frame[16] [4]), .I1(n56696), 
            .I2(GND_net), .I3(GND_net), .O(n61113));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1251 (.I0(\data_in_frame[12] [2]), .I1(n61201), 
            .I2(n56591), .I3(GND_net), .O(n56507));
    defparam i2_3_lut_adj_1251.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54996 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n72137));
    defparam byte_transmit_counter_0__bdd_4_lut_54996.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1252 (.I0(n61439), .I1(\data_in_frame[16] [3]), 
            .I2(n62654), .I3(GND_net), .O(n55576));
    defparam i2_3_lut_adj_1252.LUT_INIT = 16'h6969;
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8][5] ), .C(clk16MHz), 
           .D(n29136));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8][6] ), .C(clk16MHz), 
           .D(n29139));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8][7] ), .C(clk16MHz), 
           .D(n29142));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29838), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29837), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29836), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29835), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29834), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29833), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29832), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29831), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29830), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29829), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29828), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29827), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29826), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29825), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_in_frame[1]_c [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60890));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i13835_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][5] ), 
            .I3(PWMLimit[21]), .O(n29696));   // verilog/coms.v(148[4] 304[11])
    defparam i13835_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[8][4] ), .I1(Kp_23__N_872), 
            .I2(GND_net), .I3(GND_net), .O(n60927));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[5] [2]), .O(n60861));   // verilog/coms.v(88[17:70])
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[6] [0]), .I1(n61415), 
            .I2(GND_net), .I3(GND_net), .O(n61018));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1257 (.I0(n56581), .I1(n55540), .I2(\data_in_frame[11] [7]), 
            .I3(\data_in_frame[12] [1]), .O(n10_adj_5556));
    defparam i4_4_lut_adj_1257.LUT_INIT = 16'h9669;
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29824), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29823), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29822), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29821), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29820), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29819), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29818), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29817), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29816), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29815), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29814), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29813), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29812), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29811), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29810), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29809), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29808), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29807), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29806), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29805), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29804), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29803), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29802), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29801), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29800), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29799), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29798), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29797), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29796), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29795), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29794), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29793), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29792), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29791), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29790), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29789), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29788), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29787), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29786), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29785), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29784), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29783), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29782), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29781), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29780), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5359), .S(n60536));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13836_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][4] ), 
            .I3(PWMLimit[20]), .O(n29697));   // verilog/coms.v(148[4] 304[11])
    defparam i13836_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29779), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29778), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29777), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29776), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29775), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[4] [5]), .I1(n55544), 
            .I2(GND_net), .I3(GND_net), .O(n61455));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29774), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n61361));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29773), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29772), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29771), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29770), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29769), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29768), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13837_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][3] ), 
            .I3(PWMLimit[19]), .O(n29698));   // verilog/coms.v(148[4] 304[11])
    defparam i13837_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29767), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29766), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29765), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29764), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29763), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29762));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29761));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1260 (.I0(n64765), .I1(Kp_23__N_1067), .I2(n26077), 
            .I3(Kp_23__N_974), .O(n64771));   // verilog/coms.v(74[16:27])
    defparam i1_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29760));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29759));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29758));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29757));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1261 (.I0(n61436), .I1(n55700), .I2(n26262), 
            .I3(n64771), .O(n24870));   // verilog/coms.v(74[16:27])
    defparam i1_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1262 (.I0(n25647), .I1(n24870), .I2(\data_in_frame[9] [0]), 
            .I3(GND_net), .O(n26258));
    defparam i1_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29755));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29754));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29753));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1263 (.I0(\data_in_frame[9] [3]), .I1(n61119), 
            .I2(\data_in_frame[9] [6]), .I3(n25501), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29752));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29751));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1264 (.I0(Kp_23__N_1080), .I1(n26258), .I2(GND_net), 
            .I3(GND_net), .O(n60985));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29750));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29749));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1265 (.I0(n23700), .I1(n23704), .I2(GND_net), 
            .I3(GND_net), .O(n26262));
    defparam i1_2_lut_adj_1265.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29748));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29747));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_in_frame[8][7] ), .I1(\data_in_frame[8][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n61332));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29746));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29745));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29744));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[8][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n61458));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29743));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n61122));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29121));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13839_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8][2] ), 
            .I3(PWMLimit[18]), .O(n29700));   // verilog/coms.v(148[4] 304[11])
    defparam i13839_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2881), .D(n2_adj_5557), .S(n60535));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29742));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29741));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29739));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(\control_mode[2] ), .C(clk16MHz), .D(n29738));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode_c[3]), .C(clk16MHz), .D(n29737));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(\control_mode[4] ), .C(clk16MHz), .D(n29736));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode_c[5]), .C(clk16MHz), .D(n29735));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(\control_mode[6] ), .C(clk16MHz), .D(n29734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(\control_mode[7] ), .C(clk16MHz), .D(n29733));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n29732));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n29731));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n29730));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n29729));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n29728));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29727));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29726));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29725));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29724));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29723));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29722));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29721));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29720));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29719));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29718));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29717), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29716), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29715), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29714), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29713), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29712), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_2043__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n27760), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n27762), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_3_lut_adj_1269 (.I0(\data_in_frame[1][6] ), .I1(n56581), 
            .I2(n61122), .I3(GND_net), .O(n12_adj_5558));   // verilog/coms.v(99[12:25])
    defparam i1_3_lut_adj_1269.LUT_INIT = 16'h6969;
    SB_DFFR \FRAME_MATCHER.i_2043__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n27764), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n27766), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n27768), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n27770), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n27772), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n27774), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n27776), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n27778), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n27780), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n27782), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n27784), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n27786), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n27788), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n27790), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n27792), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n27794), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n27796), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n27798), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n27800), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n27802), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n27804), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n27806), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n27808), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n27810), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n27812), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n27814), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n27816), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n27818), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n27820), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29711), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29710), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29709), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29708), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29707), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29706), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29705), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29704), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29703), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n29702), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n29701), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n29700), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n29145));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n29698), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n29697), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n29696), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n29695), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n29694), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n29148));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n29151));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n29154));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n29157));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n29160));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29111), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29110));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29109));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29108));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29107), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29106), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29105), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n29163));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1270 (.I0(n61430), .I1(n61332), .I2(n25662), 
            .I3(n71568), .O(n18_adj_5559));   // verilog/coms.v(99[12:25])
    defparam i7_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n29166));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10]_c [0]), .C(clk16MHz), 
           .D(n29169));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10][1] ), .C(clk16MHz), 
           .D(n29172));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10][2] ), .C(clk16MHz), 
           .D(n29175));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10][3] ), .C(clk16MHz), 
           .D(n29178));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n29181));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
           .D(n29184));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n29187));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
           .D(n29190));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29104), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i8_4_lut_adj_1271 (.I0(n61458), .I1(n60924), .I2(n61352), 
            .I3(\data_in_frame[8][4] ), .O(n19_adj_5560));   // verilog/coms.v(99[12:25])
    defparam i8_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1272 (.I0(n19_adj_5560), .I1(\data_in_frame[8] [0]), 
            .I2(n18_adj_5559), .I3(n12_adj_5558), .O(n61295));   // verilog/coms.v(99[12:25])
    defparam i10_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 n72137_bdd_4_lut (.I0(n72137), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n72140));
    defparam n72137_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1273 (.I0(n25781), .I1(Kp_23__N_1301), .I2(\data_in_frame[15] [6]), 
            .I3(GND_net), .O(n60822));
    defparam i2_3_lut_adj_1273.LUT_INIT = 16'h9696;
    SB_LUT4 i19375_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n29701));   // verilog/coms.v(148[4] 304[11])
    defparam i19375_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60990));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60996));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(n25746), .I1(n60938), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1301));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1277 (.I0(n24953), .I1(n60990), .I2(n25817), 
            .I3(\data_in_frame[13] [2]), .O(n55574));
    defparam i3_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1278 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[16] [1]), 
            .I2(n60996), .I3(\data_in_frame[13] [6]), .O(n16_adj_5561));
    defparam i6_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1279 (.I0(n55574), .I1(n60979), .I2(n61323), 
            .I3(Kp_23__N_1301), .O(n17_adj_5562));
    defparam i7_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 select_1745_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5549));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut_adj_1280 (.I0(n17_adj_5562), .I1(\data_in_frame[14] [0]), 
            .I2(n16_adj_5561), .I3(n55705), .O(n62654));
    defparam i9_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i53119_3_lut (.I0(n61102), .I1(n56696), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n59688));
    defparam i53119_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(\data_in_frame[21] [2]), .I1(n25950), 
            .I2(n25923), .I3(\data_in_frame[19] [0]), .O(n10_adj_5554));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1282 (.I0(\data_in_frame[16] [0]), .I1(n61129), 
            .I2(n56075), .I3(n55679), .O(n61073));
    defparam i3_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5563));
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1284 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[15] [5]), 
            .I2(n61073), .I3(n6_adj_5563), .O(n61344));
    defparam i4_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1285 (.I0(\data_in_frame[20] [0]), .I1(n26599), 
            .I2(\data_in_frame[19] [7]), .I3(\data_in_frame[19] [5]), .O(n60906));
    defparam i1_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i11853_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27713));   // verilog/coms.v(109[34:55])
    defparam i11853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48258_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65348));
    defparam i48258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48259_4_lut (.I0(n65348), .I1(n27713), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n65349));
    defparam i48259_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48257_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65347));
    defparam i48257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51669_2_lut (.I0(n72146), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68456));
    defparam i51669_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i53479_3_lut (.I0(n72194), .I1(n71948), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70569));
    defparam i53479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5564));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19488_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n29702));   // verilog/coms.v(148[4] 304[11])
    defparam i19488_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48242_4_lut (.I0(n1_adj_5564), .I1(\data_out_frame[3][3] ), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n65332));
    defparam i48242_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i18021_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n29703));   // verilog/coms.v(148[4] 304[11])
    defparam i18021_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13843_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n29704));   // verilog/coms.v(148[4] 304[11])
    defparam i13843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48293_3_lut (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65383));
    defparam i48293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48294_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65384));
    defparam i48294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48366_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65456));
    defparam i48366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48365_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65455));
    defparam i48365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48299_3_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65389));
    defparam i48299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48300_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65390));
    defparam i48300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48348_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65438));
    defparam i48348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48347_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65437));
    defparam i48347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48335_3_lut (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65425));
    defparam i48335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1286 (.I0(\FRAME_MATCHER.i[4] ), .I1(n39431), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n110), .O(n112));
    defparam i1_2_lut_4_lut_adj_1286.LUT_INIT = 16'hfff7;
    SB_LUT4 i48336_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65426));
    defparam i48336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48303_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65393));
    defparam i48303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48302_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65392));
    defparam i48302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48362_3_lut (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65452));
    defparam i48362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48363_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65453));
    defparam i48363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48375_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65465));
    defparam i48375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48374_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65464));
    defparam i48374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48344_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65434));
    defparam i48344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48345_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65435));
    defparam i48345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48252_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65342));
    defparam i48252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48251_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65341));
    defparam i48251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51689_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68359));   // verilog/coms.v(158[12:15])
    defparam i51689_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1287 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5565), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n26729));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'haaa8;
    SB_LUT4 i51683_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68358));   // verilog/coms.v(158[12:15])
    defparam i51683_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51512_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68357));   // verilog/coms.v(158[12:15])
    defparam i51512_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51659_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68346));   // verilog/coms.v(158[12:15])
    defparam i51659_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51716_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68345));   // verilog/coms.v(158[12:15])
    defparam i51716_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16470_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n32330));   // verilog/coms.v(118[11:12])
    defparam i16470_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i13844_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n29705));   // verilog/coms.v(148[4] 304[11])
    defparam i13844_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51469_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68342));   // verilog/coms.v(158[12:15])
    defparam i51469_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13845_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n29706));   // verilog/coms.v(148[4] 304[11])
    defparam i13845_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i52021_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68337));   // verilog/coms.v(158[12:15])
    defparam i52021_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51468_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68332));   // verilog/coms.v(158[12:15])
    defparam i51468_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13846_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n29707));   // verilog/coms.v(148[4] 304[11])
    defparam i13846_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51690_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68360));   // verilog/coms.v(158[12:15])
    defparam i51690_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51577_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68295));   // verilog/coms.v(158[12:15])
    defparam i51577_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51653_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68294));   // verilog/coms.v(158[12:15])
    defparam i51653_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51568_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68293));   // verilog/coms.v(158[12:15])
    defparam i51568_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51517_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68278));   // verilog/coms.v(158[12:15])
    defparam i51517_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51543_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68273));   // verilog/coms.v(158[12:15])
    defparam i51543_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11872_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3483), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n27733));   // verilog/coms.v(158[12:15])
    defparam i11872_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i51492_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68269));   // verilog/coms.v(158[12:15])
    defparam i51492_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51732_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68268));   // verilog/coms.v(158[12:15])
    defparam i51732_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51678_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68267));   // verilog/coms.v(158[12:15])
    defparam i51678_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51489_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68265));   // verilog/coms.v(158[12:15])
    defparam i51489_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51488_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68264));   // verilog/coms.v(158[12:15])
    defparam i51488_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51487_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68263));   // verilog/coms.v(158[12:15])
    defparam i51487_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51782_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68262));   // verilog/coms.v(158[12:15])
    defparam i51782_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51714_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68261));   // verilog/coms.v(158[12:15])
    defparam i51714_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1288 (.I0(n62406), .I1(n64881), .I2(n64845), 
            .I3(n61367), .O(n64849));
    defparam i1_4_lut_adj_1288.LUT_INIT = 16'h8020;
    SB_LUT4 i1_4_lut_adj_1289 (.I0(\data_in_frame[18] [5]), .I1(n60960), 
            .I2(n56575), .I3(\data_in_frame[22] [7]), .O(n64677));
    defparam i1_4_lut_adj_1289.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1290 (.I0(\data_in_frame[23] [0]), .I1(n64849), 
            .I2(n55989), .I3(n61051), .O(n64851));
    defparam i1_4_lut_adj_1290.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5540));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18959_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n29708));   // verilog/coms.v(148[4] 304[11])
    defparam i18959_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13848_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n29709));   // verilog/coms.v(148[4] 304[11])
    defparam i13848_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[8][2] ), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61430));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i13849_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n29710));   // verilog/coms.v(148[4] 304[11])
    defparam i13849_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut_adj_1292 (.I0(n64851), .I1(n64677), .I2(n55989), 
            .I3(n61051), .O(n33_adj_5555));
    defparam i1_4_lut_adj_1292.LUT_INIT = 16'h8228;
    SB_LUT4 select_787_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5306));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5539));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5538));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5304));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5537));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13850_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n29711));   // verilog/coms.v(148[4] 304[11])
    defparam i13850_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18673_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n29712));   // verilog/coms.v(148[4] 304[11])
    defparam i18673_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1293 (.I0(\data_in_frame[7] [7]), .I1(n61027), 
            .I2(\data_in_frame[1]_c [5]), .I3(GND_net), .O(n25662));
    defparam i2_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5536));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5535));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5534));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18716_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n29713));   // verilog/coms.v(148[4] 304[11])
    defparam i18716_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5533));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i18762_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n29714));   // verilog/coms.v(148[4] 304[11])
    defparam i18762_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1194_9_lut (.I0(n60666), .I1(byte_transmit_counter_c[7]), 
            .I2(GND_net), .I3(n53699), .O(n60674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1194_8_lut (.I0(n60666), .I1(byte_transmit_counter_c[6]), 
            .I2(GND_net), .I3(n53698), .O(n60668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_8 (.CI(n53698), .I0(byte_transmit_counter_c[6]), .I1(GND_net), 
            .CO(n53699));
    SB_LUT4 add_1194_7_lut (.I0(n60666), .I1(byte_transmit_counter_c[5]), 
            .I2(GND_net), .I3(n53697), .O(n60669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_7 (.CI(n53697), .I0(byte_transmit_counter_c[5]), .I1(GND_net), 
            .CO(n53698));
    SB_LUT4 i13897_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [5]), 
            .I3(neopxl_color[5]), .O(n29758));   // verilog/coms.v(130[12] 305[6])
    defparam i13897_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 add_1194_6_lut (.I0(n60666), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n53696), .O(n60670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_6 (.CI(n53696), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n53697));
    SB_LUT4 add_1194_5_lut (.I0(n60666), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n53695), .O(n60671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_5 (.CI(n53695), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n53696));
    SB_LUT4 add_1194_4_lut (.I0(n60666), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n53694), .O(n60672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_4 (.CI(n53694), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n53695));
    SB_LUT4 add_1194_3_lut (.I0(n60666), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n53693), .O(n60673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_3 (.CI(n53693), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n53694));
    SB_LUT4 add_1194_2_lut (.I0(n60666), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n60667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n53693));
    SB_LUT4 i13854_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10][3] ), 
            .I3(PWMLimit[3]), .O(n29715));   // verilog/coms.v(148[4] 304[11])
    defparam i13854_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5531));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13855_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10][2] ), 
            .I3(PWMLimit[2]), .O(n29716));   // verilog/coms.v(148[4] 304[11])
    defparam i13855_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5530));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13856_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[10][1] ), 
            .I3(PWMLimit[1]), .O(n29717));   // verilog/coms.v(148[4] 304[11])
    defparam i13856_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i51804_2_lut_4_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(n39431), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n37941), .O(n68422));
    defparam i51804_2_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 select_787_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5529));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13886_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [0]), 
            .I3(neopxl_color[16]), .O(n29747));   // verilog/coms.v(130[12] 305[6])
    defparam i13886_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_787_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5528));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5527));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13898_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [4]), 
            .I3(neopxl_color[4]), .O(n29759));   // verilog/coms.v(130[12] 305[6])
    defparam i13898_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13902_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n29763));   // verilog/coms.v(148[4] 304[11])
    defparam i13902_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_1294 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[2] [1]), .O(n61352));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5526));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13882_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [4]), 
            .I3(neopxl_color[20]), .O(n29743));   // verilog/coms.v(130[12] 305[6])
    defparam i13882_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13894_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [0]), 
            .I3(neopxl_color[8]), .O(n29755));   // verilog/coms.v(130[12] 305[6])
    defparam i13894_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1295 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1] [1]), 
            .I2(n61261), .I3(\data_in_frame[1]_c [0]), .O(n25669));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i22020_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [5]), 
            .I3(neopxl_color[13]), .O(n29750));   // verilog/coms.v(130[12] 305[6])
    defparam i22020_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(\data_in_frame[10] [7]), .I1(n60987), 
            .I2(n60938), .I3(GND_net), .O(n60940));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5525));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13883_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [3]), 
            .I3(neopxl_color[19]), .O(n29744));   // verilog/coms.v(130[12] 305[6])
    defparam i13883_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n37935));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h0404;
    SB_LUT4 i15_2_lut_3_lut (.I0(\data_in_frame[10] [7]), .I1(n60987), .I2(n25746), 
            .I3(GND_net), .O(n59626));
    defparam i15_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13895_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [7]), 
            .I3(neopxl_color[7]), .O(n29756));   // verilog/coms.v(130[12] 305[6])
    defparam i13895_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13888_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [6]), 
            .I3(neopxl_color[14]), .O(n29749));   // verilog/coms.v(130[12] 305[6])
    defparam i13888_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_787_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5524));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19376_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [0]), 
            .I3(neopxl_color[0]), .O(n29108));   // verilog/coms.v(130[12] 305[6])
    defparam i19376_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13881_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [5]), 
            .I3(neopxl_color[21]), .O(n29742));   // verilog/coms.v(130[12] 305[6])
    defparam i13881_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13893_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [1]), 
            .I3(neopxl_color[9]), .O(n29754));   // verilog/coms.v(130[12] 305[6])
    defparam i13893_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1298 (.I0(n60947), .I1(n55617), .I2(\data_in_frame[21] [4]), 
            .I3(GND_net), .O(n61301));
    defparam i1_2_lut_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5523));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i22015_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [4]), 
            .I3(neopxl_color[12]), .O(n29751));   // verilog/coms.v(130[12] 305[6])
    defparam i22015_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13903_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n29764));   // verilog/coms.v(148[4] 304[11])
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_4_lut_adj_1299 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[20] [3]), .I3(\data_in_frame[20] [4]), .O(n64729));
    defparam i1_3_lut_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1300 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n61412), .O(n23700));
    defparam i1_2_lut_3_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5522));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_33_lut  (.I0(n68261), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n54545), .O(n27820)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_32_lut  (.I0(n68262), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n54544), .O(n27818)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13884_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [2]), 
            .I3(neopxl_color[18]), .O(n29745));   // verilog/coms.v(130[12] 305[6])
    defparam i13884_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_32  (.CI(n54544), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n54545));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_31_lut  (.I0(n68263), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n54543), .O(n27816)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_31  (.CI(n54543), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n54544));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_30_lut  (.I0(n68264), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n54542), .O(n27814)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13896_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [6]), 
            .I3(neopxl_color[6]), .O(n29757));   // verilog/coms.v(130[12] 305[6])
    defparam i13896_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_30  (.CI(n54542), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n54543));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_29_lut  (.I0(n68265), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n54541), .O(n27812)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_4_lut_adj_1301 (.I0(\data_in_frame[10][3] ), .I1(n60779), 
            .I2(n61326), .I3(n6_adj_5566), .O(n26274));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_29  (.CI(n54541), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n54542));
    SB_LUT4 i13887_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [7]), 
            .I3(neopxl_color[15]), .O(n29748));   // verilog/coms.v(130[12] 305[6])
    defparam i13887_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_28_lut  (.I0(n68267), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n54540), .O(n27810)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_28  (.CI(n54540), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n54541));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1302 (.I0(n25598), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[0] [1]), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_27_lut  (.I0(n68268), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n54539), .O(n27808)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_27  (.CI(n54539), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n54540));
    SB_LUT4 i13904_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n29765));   // verilog/coms.v(148[4] 304[11])
    defparam i13904_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_26_lut  (.I0(n68269), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n54538), .O(n27806)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_26  (.CI(n54538), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n54539));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_25_lut  (.I0(n68273), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n54537), .O(n27804)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_25  (.CI(n54537), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n54538));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_24_lut  (.I0(n68278), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n54536), .O(n27802)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_24  (.CI(n54536), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n54537));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_23_lut  (.I0(n68293), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n54535), .O(n27800)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54991 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n72131));
    defparam byte_transmit_counter_0__bdd_4_lut_54991.LUT_INIT = 16'he4aa;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_23  (.CI(n54535), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n54536));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_22_lut  (.I0(n68294), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n54534), .O(n27798)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13899_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [3]), 
            .I3(neopxl_color[3]), .O(n29760));   // verilog/coms.v(130[12] 305[6])
    defparam i13899_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13901_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [1]), 
            .I3(neopxl_color[1]), .O(n29762));   // verilog/coms.v(130[12] 305[6])
    defparam i13901_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_22  (.CI(n54534), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n54535));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_21_lut  (.I0(n68295), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n54533), .O(n27796)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_21  (.CI(n54533), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n54534));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_20_lut  (.I0(n68332), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n54532), .O(n27794)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_20  (.CI(n54532), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n54533));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_19_lut  (.I0(n68337), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n54531), .O(n27792)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut_adj_1303 (.I0(reset), .I1(n39431), .I2(n10_adj_5567), 
            .I3(GND_net), .O(n60769));
    defparam i1_2_lut_3_lut_adj_1303.LUT_INIT = 16'hfbfb;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_19  (.CI(n54531), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n54532));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_18_lut  (.I0(n68342), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n54530), .O(n27790)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1304 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[15] [2]), 
            .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5521));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1304.LUT_INIT = 16'ha088;
    SB_LUT4 i13905_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n29766));   // verilog/coms.v(148[4] 304[11])
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5520));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13906_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n29767));   // verilog/coms.v(148[4] 304[11])
    defparam i13906_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1305 (.I0(n25825), .I1(\data_in_frame[12] [5]), 
            .I2(n56127), .I3(\data_in_frame[10][1] ), .O(n64933));
    defparam i1_2_lut_3_lut_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5519));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5518));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13907_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n29768));   // verilog/coms.v(148[4] 304[11])
    defparam i13907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13908_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n29769));   // verilog/coms.v(148[4] 304[11])
    defparam i13908_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5517));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1306 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26126));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1306.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1307 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [5]), 
            .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5516));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1307.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26447));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1309 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [4]), 
            .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5515));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1309.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5568));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_220_i3_4_lut (.I0(n5_adj_5568), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n63365), .I3(n63147), .O(n3_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_220_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13909_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n29770));   // verilog/coms.v(148[4] 304[11])
    defparam i13909_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n72131_bdd_4_lut (.I0(n72131), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n72134));
    defparam n72131_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_219_i3_4_lut (.I0(n56541), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5569), .I3(n60790), .O(n3_adj_5402));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_219_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i51736_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68380));   // verilog/coms.v(158[12:15])
    defparam i51736_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13910_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n29771));   // verilog/coms.v(148[4] 304[11])
    defparam i13910_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13418_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n29279));   // verilog/coms.v(130[12] 305[6])
    defparam i13418_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[14] [5]), .I1(n26274), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5570));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5512));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13260_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29121));   // verilog/coms.v(130[12] 305[6])
    defparam i13260_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13419_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n29280));   // verilog/coms.v(130[12] 305[6])
    defparam i13419_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13420_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n29281));   // verilog/coms.v(130[12] 305[6])
    defparam i13420_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1312 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1312.LUT_INIT = 16'ha088;
    SB_LUT4 i13421_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n29282));   // verilog/coms.v(130[12] 305[6])
    defparam i13421_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13422_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n29283));   // verilog/coms.v(130[12] 305[6])
    defparam i13422_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1313 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [7]), 
            .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5510));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1313.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n60900), .I3(n61137), .O(n3_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i51727_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68377));   // verilog/coms.v(158[12:15])
    defparam i51727_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13911_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n29772));   // verilog/coms.v(148[4] 304[11])
    defparam i13911_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13423_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n29284));   // verilog/coms.v(130[12] 305[6])
    defparam i13423_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5509));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i52284_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68375));   // verilog/coms.v(158[12:15])
    defparam i52284_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13424_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n29285));   // verilog/coms.v(130[12] 305[6])
    defparam i13424_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1314 (.I0(n55646), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [3]), .I3(\data_out_frame[23] [2]), 
            .O(n63372));
    defparam i3_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1315 (.I0(n61452), .I1(n55517), .I2(n63372), 
            .I3(GND_net), .O(n14_adj_5571));
    defparam i5_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i13425_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n29286));   // verilog/coms.v(130[12] 305[6])
    defparam i13425_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5508));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1316 (.I0(\data_out_frame[21] [1]), .I1(n56573), 
            .I2(n25874), .I3(n55696), .O(n15_adj_5572));
    defparam i6_4_lut_adj_1316.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54986 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n72125));
    defparam byte_transmit_counter_0__bdd_4_lut_54986.LUT_INIT = 16'he4aa;
    SB_LUT4 i8_4_lut_adj_1317 (.I0(n15_adj_5572), .I1(n61378), .I2(n14_adj_5571), 
            .I3(n61195), .O(n63365));
    defparam i8_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i13426_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n29287));   // verilog/coms.v(130[12] 305[6])
    defparam i13426_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n72125_bdd_4_lut (.I0(n72125), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n65364));
    defparam n72125_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13427_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n29288));   // verilog/coms.v(130[12] 305[6])
    defparam i13427_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13428_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n29289));   // verilog/coms.v(130[12] 305[6])
    defparam i13428_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_out_frame[21] [0]), .I1(n24820), 
            .I2(GND_net), .I3(GND_net), .O(n61216));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5507));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13429_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n29290));   // verilog/coms.v(130[12] 305[6])
    defparam i13429_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1319 (.I0(\data_out_frame[22] [7]), .I1(n55893), 
            .I2(n26398), .I3(\data_out_frame[23] [1]), .O(n61378));
    defparam i3_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i13430_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n29291));   // verilog/coms.v(130[12] 305[6])
    defparam i13430_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5506));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1320 (.I0(n61427), .I1(n61009), .I2(n61349), 
            .I3(\data_out_frame[17] [0]), .O(n14_adj_5573));
    defparam i6_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1321 (.I0(n26560), .I1(n61375), .I2(n61307), 
            .I3(n26555), .O(n13_adj_5574));
    defparam i5_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1322 (.I0(\data_out_frame[23] [0]), .I1(n13_adj_5574), 
            .I2(n14_adj_5573), .I3(GND_net), .O(n61137));
    defparam i1_3_lut_adj_1322.LUT_INIT = 16'h6969;
    SB_LUT4 i5_3_lut_adj_1323 (.I0(\data_out_frame[16] [4]), .I1(n61378), 
            .I2(n55519), .I3(GND_net), .O(n14_adj_5575));
    defparam i5_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1324 (.I0(n61137), .I1(n61216), .I2(\data_out_frame[20] [7]), 
            .I3(n60957), .O(n15_adj_5576));
    defparam i6_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i13431_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n29292));   // verilog/coms.v(130[12] 305[6])
    defparam i13431_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13432_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n29293));   // verilog/coms.v(130[12] 305[6])
    defparam i13432_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_4_lut_adj_1325 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [2]), 
            .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1325.LUT_INIT = 16'ha088;
    SB_LUT4 i13433_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n29294));   // verilog/coms.v(130[12] 305[6])
    defparam i13433_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i8_4_lut_adj_1326 (.I0(n15_adj_5576), .I1(n55631), .I2(n14_adj_5575), 
            .I3(\data_out_frame[18] [5]), .O(n63147));
    defparam i8_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1327 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5577));
    defparam i2_2_lut_adj_1327.LUT_INIT = 16'h6666;
    SB_LUT4 i13434_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n29295));   // verilog/coms.v(130[12] 305[6])
    defparam i13434_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1328 (.I0(n7_adj_5577), .I1(n63147), .I2(n61137), 
            .I3(n62513), .O(n60790));
    defparam i4_4_lut_adj_1328.LUT_INIT = 16'h9669;
    SB_LUT4 i18860_1_lut (.I0(PWMLimit[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n34686));   // verilog/coms.v(130[12] 305[6])
    defparam i18860_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13435_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n29296));   // verilog/coms.v(130[12] 305[6])
    defparam i13435_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13436_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n29297));   // verilog/coms.v(130[12] 305[6])
    defparam i13436_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13437_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n29298));   // verilog/coms.v(130[12] 305[6])
    defparam i13437_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13438_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n29299));   // verilog/coms.v(130[12] 305[6])
    defparam i13438_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1329 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [4]), 
            .I2(n56591), .I3(n6_adj_5570), .O(n61102));
    defparam i4_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i13439_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n29300));   // verilog/coms.v(130[12] 305[6])
    defparam i13439_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13440_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n29301));   // verilog/coms.v(130[12] 305[6])
    defparam i13440_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13448_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n29309));   // verilog/coms.v(130[12] 305[6])
    defparam i13448_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i22018_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n29773));   // verilog/coms.v(148[4] 304[11])
    defparam i22018_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13447_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n29308));   // verilog/coms.v(130[12] 305[6])
    defparam i13447_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13446_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n29307));   // verilog/coms.v(130[12] 305[6])
    defparam i13446_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22019_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n29774));   // verilog/coms.v(148[4] 304[11])
    defparam i22019_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13445_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n29306));   // verilog/coms.v(130[12] 305[6])
    defparam i13445_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13914_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n29775));   // verilog/coms.v(148[4] 304[11])
    defparam i13914_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13444_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n29305));   // verilog/coms.v(130[12] 305[6])
    defparam i13444_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13443_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n29304));   // verilog/coms.v(130[12] 305[6])
    defparam i13443_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13442_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n29303));   // verilog/coms.v(130[12] 305[6])
    defparam i13442_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13441_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n29302));   // verilog/coms.v(130[12] 305[6])
    defparam i13441_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1330 (.I0(\data_out_frame[21] [2]), .I1(n26560), 
            .I2(n55598), .I3(\data_out_frame[23] [4]), .O(n61251));
    defparam i2_3_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1331 (.I0(\data_out_frame[23] [6]), .I1(n62642), 
            .I2(\data_out_frame[21] [5]), .I3(\data_out_frame[19] [3]), 
            .O(n61421));
    defparam i1_2_lut_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1332 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[15] [1]), .I3(n4_adj_5578), .O(n61156));
    defparam i1_2_lut_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13915_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n29776));   // verilog/coms.v(148[4] 304[11])
    defparam i13915_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1333 (.I0(n62684), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n56626));
    defparam i1_2_lut_adj_1333.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1334 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[5] [3]), .O(n10_adj_5579));
    defparam i2_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1335 (.I0(n61227), .I1(n56578), .I2(n56626), 
            .I3(n61233), .O(n10_adj_5580));
    defparam i4_4_lut_adj_1335.LUT_INIT = 16'h9669;
    SB_LUT4 i18756_1_lut (.I0(PWMLimit[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n34584));   // verilog/coms.v(130[12] 305[6])
    defparam i18756_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13916_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n29777));   // verilog/coms.v(148[4] 304[11])
    defparam i13916_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_217_i3_4_lut (.I0(n60790), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5580), .I3(n56541), .O(n3_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_18  (.CI(n54530), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n54531));
    SB_LUT4 i6_2_lut_3_lut (.I0(\data_out_frame[6] [1]), .I1(n25461), .I2(\data_out_frame[8][7] ), 
            .I3(GND_net), .O(n18_adj_5581));   // verilog/coms.v(77[16:43])
    defparam i6_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(n56675), .I1(n25927), .I2(GND_net), 
            .I3(GND_net), .O(n61227));
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[25] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5582));
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1338 (.I0(n61188), .I1(n55650), .I2(\data_out_frame[22] [4]), 
            .I3(n6_adj_5582), .O(n60900));
    defparam i4_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n25465));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i13385_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29246));
    defparam i13385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13917_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[15] ), .O(n29778));   // verilog/coms.v(148[4] 304[11])
    defparam i13917_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_216_i3_3_lut (.I0(n60900), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n61227), .I3(GND_net), .O(n3_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 select_787_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13918_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[14] ), .O(n29779));   // verilog/coms.v(148[4] 304[11])
    defparam i13918_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1340 (.I0(n62686), .I1(n56573), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n60957));
    defparam i2_3_lut_adj_1340.LUT_INIT = 16'h6969;
    SB_LUT4 i13382_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29243));
    defparam i13382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_17_lut  (.I0(n68345), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n54529), .O(n27788)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13919_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[13] ), .O(n29780));   // verilog/coms.v(148[4] 304[11])
    defparam i13919_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61385));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i13379_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29240));
    defparam i13379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13371_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29232));
    defparam i13371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n60793));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n61230));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\data_out_frame[22] [5]), .I1(n55644), 
            .I2(GND_net), .I3(GND_net), .O(n61188));
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_17  (.CI(n54529), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n54530));
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n60693));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i13368_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29229));
    defparam i13368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13363_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29224));
    defparam i13363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13920_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[12] ), .O(n29781));   // verilog/coms.v(148[4] 304[11])
    defparam i13920_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5494));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5583));
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1346 (.I0(n24820), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [5]), .I3(n6_adj_5583), .O(n61375));
    defparam i4_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1347 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[20] [7]), 
            .I2(n55639), .I3(n56501), .O(n12_adj_5584));
    defparam i5_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1348 (.I0(\data_out_frame[21] [1]), .I1(n12_adj_5584), 
            .I2(n60957), .I3(n56624), .O(n62684));
    defparam i6_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1349 (.I0(n62684), .I1(n61375), .I2(n55515), 
            .I3(n61089), .O(n20_adj_5585));
    defparam i8_4_lut_adj_1349.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1350 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n60690));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1350.LUT_INIT = 16'h5100;
    SB_LUT4 i7_4_lut_adj_1351 (.I0(n56632), .I1(n55534), .I2(n56492), 
            .I3(n61188), .O(n19_adj_5586));
    defparam i7_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i13359_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29220));
    defparam i13359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13356_3_lut_4_lut (.I0(n8_adj_5327), .I1(n60769), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29217));
    defparam i13356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1352 (.I0(n55598), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[21] [0]), .I3(n62914), .O(n21_adj_5587));
    defparam i9_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_16_lut  (.I0(n68346), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n54528), .O(n27786)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_16  (.CI(n54528), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n54529));
    SB_LUT4 i6_4_lut_adj_1353 (.I0(n21_adj_5587), .I1(\data_out_frame[24] [4]), 
            .I2(n19_adj_5586), .I3(n20_adj_5585), .O(n26_adj_5588));
    defparam i6_4_lut_adj_1353.LUT_INIT = 16'h9669;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_15_lut  (.I0(n68357), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n54527), .O(n27784)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13921_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[11] ), .O(n29782));   // verilog/coms.v(148[4] 304[11])
    defparam i13921_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_15  (.CI(n54527), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n54528));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_14_lut  (.I0(n68358), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n54526), .O(n27782)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_14  (.CI(n54526), .I0(n28031), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n54527));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_13_lut  (.I0(n68359), .I1(n28031), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n54525), .O(n27780)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13922_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[10] ), .O(n29783));   // verilog/coms.v(148[4] 304[11])
    defparam i13922_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14_4_lut_adj_1354 (.I0(\data_out_frame[23] [5]), .I1(\data_out_frame[23] [0]), 
            .I2(n61421), .I3(\data_out_frame[24] [5]), .O(n34));
    defparam i14_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1355 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n60689));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1355.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12_4_lut (.I0(n60819), .I1(\data_out_frame[25] [5]), .I2(\data_out_frame[23] [7]), 
            .I3(n61042), .O(n32));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1356 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n60688));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1356.LUT_INIT = 16'h5100;
    SB_LUT4 i11_4_lut (.I0(n61230), .I1(n60793), .I2(\data_out_frame[24] [6]), 
            .I3(\data_out_frame[25] [6]), .O(n31_adj_5589));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1357 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[23] [1]), .I3(n55731), .O(n35));
    defparam i15_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1358 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n60687));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1358.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i17_4_lut_adj_1359 (.I0(\data_out_frame[24] [7]), .I1(n34), 
            .I2(n26_adj_5588), .I3(n61385), .O(n37_adj_5590));
    defparam i17_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1360 (.I0(n37_adj_5590), .I1(n35), .I2(n31_adj_5589), 
            .I3(n32), .O(n25927));
    defparam i19_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1361 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n60680));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1361.LUT_INIT = 16'h5100;
    SB_LUT4 i2_2_lut_4_lut_adj_1362 (.I0(n61355), .I1(n62822), .I2(n61110), 
            .I3(n61358), .O(n10_adj_5591));   // verilog/coms.v(88[17:63])
    defparam i2_2_lut_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_215_i3_4_lut (.I0(n25927), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n6_adj_5592), .I3(n56675), .O(n3_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_215_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1363 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n60694));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1363.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1364 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n60683));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1364.LUT_INIT = 16'h5100;
    SB_LUT4 i13923_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[9] ), .O(n29784));   // verilog/coms.v(148[4] 304[11])
    defparam i13923_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5489));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1365 (.I0(\data_in_frame[14] [3]), .I1(n56507), 
            .I2(\data_in_frame[16] [4]), .I3(n56563), .O(n25950));
    defparam i2_3_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(\data_in_frame[14] [3]), .I1(n56507), 
            .I2(n56565), .I3(GND_net), .O(n60973));
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1367 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n60691));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1367.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5488));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51677_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68369));   // verilog/coms.v(158[12:15])
    defparam i51677_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i51697_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68367));   // verilog/coms.v(158[12:15])
    defparam i51697_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[14] [3]), .I1(n56507), 
            .I2(n56696), .I3(GND_net), .O(n61185));
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1369 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n60682));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1369.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1370 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n60681));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1370.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1371 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n60685));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1371.LUT_INIT = 16'h5100;
    SB_LUT4 i13305_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29166));
    defparam i13305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1372 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n60686));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1372.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1373 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n60679));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1373.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1374 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n60692));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1374.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5486));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1375 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n60684));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1375.LUT_INIT = 16'h5100;
    SB_LUT4 select_787_Select_213_i3_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n56543), .I3(n61207), .O(n3_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_213_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1376 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61042));
    defparam i1_2_lut_adj_1376.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1377 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n25879));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1378 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[18] [7]), 
            .I2(n25994), .I3(n55945), .O(n14_adj_5593));
    defparam i5_3_lut_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i13302_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29163));
    defparam i13302_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n61006));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 i51696_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68366));   // verilog/coms.v(158[12:15])
    defparam i51696_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1380 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[14] [3]), 
            .I2(n61391), .I3(\data_out_frame[7] [5]), .O(n6_adj_5594));
    defparam i1_2_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i13924_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n29785));   // verilog/coms.v(148[4] 304[11])
    defparam i13924_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13925_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [7]), 
            .I3(\Kp[7] ), .O(n29786));   // verilog/coms.v(148[4] 304[11])
    defparam i13925_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_211_i3_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5595), .I3(n55523), 
            .O(n3_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i13299_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29160));
    defparam i13299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13296_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29157));
    defparam i13296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13293_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29154));
    defparam i13293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1381 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(n4_adj_5596), .I3(GND_net), .O(n55741));   // verilog/coms.v(78[16:27])
    defparam i2_2_lut_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(\data_out_frame[11] [5]), .I1(n55368), 
            .I2(n26185), .I3(GND_net), .O(n61147));
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1383 (.I0(n1168), .I1(n60864), .I2(n10_adj_5597), 
            .I3(n1130), .O(n26185));
    defparam i5_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_210_i3_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5598), .I3(n61181), 
            .O(n3_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_2_lut_3_lut_adj_1384 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n10_adj_5599));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i13290_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29151));
    defparam i13290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13287_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29148));
    defparam i13287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5481));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13926_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [6]), 
            .I3(\Kp[6] ), .O(n29787));   // verilog/coms.v(148[4] 304[11])
    defparam i13926_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1385 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n62824), .I3(GND_net), .O(n62914));
    defparam i2_3_lut_adj_1385.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n61150));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_LUT4 i13284_3_lut_4_lut (.I0(n8_adj_11), .I1(n60769), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29145));
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[12] [0]), .I3(GND_net), .O(n61288));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[8][4] ), 
            .I2(\data_out_frame[11] [0]), .I3(n26405), .O(n14_adj_5600));   // verilog/coms.v(75[16:27])
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1388 (.I0(n61039), .I1(\data_in_frame[19] [2]), 
            .I2(n56565), .I3(GND_net), .O(n61062));
    defparam i2_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1389 (.I0(\data_out_frame[21] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(n61418), .I3(n61291), .O(n10_adj_5601));
    defparam i4_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5480));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_adj_1390 (.I0(n55731), .I1(n10_adj_5601), .I2(n26147), 
            .I3(GND_net), .O(n23471));
    defparam i5_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[4] [1]), 
            .I2(n61000), .I3(n60850), .O(n26215));   // verilog/coms.v(78[16:43])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13551_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29412));
    defparam i13551_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[4] [1]), 
            .I2(n61000), .I3(n60803), .O(n9_adj_5602));   // verilog/coms.v(78[16:43])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1391 (.I0(n55598), .I1(n56632), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n56675));
    defparam i2_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1392 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[14] [7]), .I3(n25658), .O(n61276));
    defparam i2_3_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1393 (.I0(\data_out_frame[18] [1]), .I1(n61159), 
            .I2(n56069), .I3(GND_net), .O(n23430));
    defparam i2_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1394 (.I0(\data_out_frame[20] [5]), .I1(n55644), 
            .I2(n56492), .I3(n55534), .O(n61207));
    defparam i2_3_lut_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1395 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[10] [5]), 
            .I2(n25732), .I3(n26220), .O(n25658));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5478));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13554_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29415));
    defparam i13554_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1396 (.I0(n61273), .I1(n26304), .I2(\data_out_frame[18] [0]), 
            .I3(n61364), .O(n10_adj_5603));
    defparam i4_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(\data_out_frame[20] [2]), .I1(n55499), 
            .I2(n61024), .I3(GND_net), .O(n6_adj_5604));
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'h9696;
    SB_LUT4 i13557_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29418));
    defparam i13557_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_out_frame[21] [7]), .I1(n62513), 
            .I2(n55515), .I3(GND_net), .O(n55534));
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1399 (.I0(\data_out_frame[18] [2]), .I1(n56583), 
            .I2(\data_out_frame[16] [0]), .I3(n6_adj_5605), .O(n61159));
    defparam i4_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i13560_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29421));
    defparam i13560_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13563_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29424));
    defparam i13563_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1400 (.I0(n60828), .I1(n61254), .I2(n26250), 
            .I3(\data_in_frame[9] [2]), .O(n60944));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i13927_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [5]), 
            .I3(\Kp[5] ), .O(n29788));   // verilog/coms.v(148[4] 304[11])
    defparam i13927_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i4_4_lut_adj_1401 (.I0(\data_in_frame[16] [6]), .I1(n60973), 
            .I2(\data_in_frame[19] [1]), .I3(\data_in_frame[16] [5]), .O(n10_adj_5606));
    defparam i4_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1402 (.I0(n60828), .I1(n61254), .I2(n26250), 
            .I3(n55521), .O(n61436));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i13566_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29427));
    defparam i13566_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_out_frame[17] [5]), .I1(n55715), 
            .I2(n25490), .I3(GND_net), .O(n61364));
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(n60779), .I3(GND_net), .O(n6_adj_5607));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1405 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[13] [5]), .I3(n24849), .O(n10_adj_5608));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_out_frame[16] [0]), .I1(n56537), 
            .I2(n61162), .I3(GND_net), .O(n6_adj_5609));
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i13569_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29430));
    defparam i13569_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13928_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n29789));   // verilog/coms.v(148[4] 304[11])
    defparam i13928_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1407 (.I0(n24849), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n61162));
    defparam i1_2_lut_3_lut_adj_1407.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_out_frame[16] [1]), .I1(n55646), 
            .I2(GND_net), .I3(GND_net), .O(n56583));
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(\data_out_frame[11] [6]), .I1(n60867), 
            .I2(GND_net), .I3(GND_net), .O(n61270));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1410 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5610));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1411 (.I0(n7_adj_5610), .I1(n26185), .I2(n62686), 
            .I3(n61270), .O(n56192));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1411.LUT_INIT = 16'h9669;
    SB_LUT4 i13929_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [3]), 
            .I3(\Kp[3] ), .O(n29790));   // verilog/coms.v(148[4] 304[11])
    defparam i13929_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_out_frame[18] [4]), .I1(n55696), 
            .I2(GND_net), .I3(GND_net), .O(n60951));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i13572_3_lut_4_lut (.I0(n39467), .I1(n60769), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29433));
    defparam i13572_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1413 (.I0(n26398), .I1(n61024), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n55893));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i13415_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29276));
    defparam i13415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13930_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [2]), 
            .I3(\Kp[2] ), .O(n29791));   // verilog/coms.v(148[4] 304[11])
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1414 (.I0(\data_out_frame[19] [5]), .I1(n62635), 
            .I2(n62923), .I3(GND_net), .O(n26147));
    defparam i2_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1415 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(n55137), 
            .I2(n25249), .I3(GND_net), .O(n32326));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_adj_1415.LUT_INIT = 16'h2020;
    SB_LUT4 i5_3_lut_adj_1416 (.I0(n61102), .I1(n10_adj_5606), .I2(\data_in_frame[18] [7]), 
            .I3(GND_net), .O(n25923));
    defparam i5_3_lut_adj_1416.LUT_INIT = 16'h6969;
    SB_LUT4 i51740_2_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(n25249), 
            .I2(GND_net), .I3(GND_net), .O(n68385));   // verilog/coms.v(18[27:29])
    defparam i51740_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut_adj_1417 (.I0(n26147), .I1(n55893), .I2(\data_out_frame[20] [0]), 
            .I3(n60951), .O(n55515));
    defparam i3_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1418 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[7] [5]), .I3(n25987), .O(n12_adj_5611));   // verilog/coms.v(73[16:69])
    defparam i5_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i13412_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29273));
    defparam i13412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(n55696), .I1(n55388), .I2(\data_out_frame[18] [3]), 
            .I3(\data_out_frame[18] [4]), .O(n62513));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16479_4_lut (.I0(n32326), .I1(n68385), .I2(Kp_23__N_1748), 
            .I3(n33_adj_5555), .O(n27414));   // verilog/coms.v(18[27:29])
    defparam i16479_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5612));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1421 (.I0(\data_in_frame[5] [4]), .I1(n12_adj_5611), 
            .I2(n61261), .I3(\data_in_frame[5] [3]), .O(n56127));   // verilog/coms.v(73[16:69])
    defparam i6_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i13931_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n29792));   // verilog/coms.v(148[4] 304[11])
    defparam i13931_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13533_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29394));
    defparam i13533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1422 (.I0(\data_out_frame[17] [4]), .I1(n4_adj_5578), 
            .I2(n25490), .I3(n6_adj_5612), .O(n62923));
    defparam i4_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1423 (.I0(n62686), .I1(n55517), .I2(n56192), 
            .I3(n25874), .O(n55696));
    defparam i2_3_lut_4_lut_adj_1423.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1424 (.I0(\data_out_frame[16] [2]), .I1(n56192), 
            .I2(\data_out_frame[16] [1]), .I3(n55646), .O(n55388));
    defparam i2_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\data_out_frame[19] [7]), .I1(n25490), 
            .I2(GND_net), .I3(GND_net), .O(n61273));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1426 (.I0(\data_out_frame[19] [6]), .I1(n62923), 
            .I2(GND_net), .I3(GND_net), .O(n61204));
    defparam i1_2_lut_adj_1426.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1427 (.I0(n61204), .I1(\data_out_frame[22] [2]), 
            .I2(\data_out_frame[20] [0]), .I3(n61273), .O(n10_adj_5613));
    defparam i4_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1428 (.I0(\data_out_frame[11] [6]), .I1(n60867), 
            .I2(n10_adj_5608), .I3(n55578), .O(n55646));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i13932_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n29793));   // verilog/coms.v(148[4] 304[11])
    defparam i13932_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1429 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [3]), .I3(\data_out_frame[20] [2]), 
            .O(n26398));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1430 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(n56192), .I3(n56583), .O(n55631));
    defparam i1_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1431 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n26304));
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'h6666;
    SB_LUT4 i13536_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29397));
    defparam i13536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1432 (.I0(n24849), .I1(n61150), .I2(n10_adj_5603), 
            .I3(\data_out_frame[15] [6]), .O(n62824));
    defparam i5_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1433 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n61147), .I3(n6_adj_5609), .O(n56069));
    defparam i4_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1434 (.I0(n61144), .I1(\data_out_frame[15] [6]), 
            .I2(n56069), .I3(n61165), .O(n10_adj_5614));
    defparam i4_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i13539_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29400));
    defparam i13539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(\data_out_frame[19] [6]), .I1(n62923), 
            .I2(n56728), .I3(\data_out_frame[22] [0]), .O(n61418));
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\data_in_frame[1]_c [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n61012));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h6666;
    SB_LUT4 i13542_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29403));
    defparam i13542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13933_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n29794));   // verilog/coms.v(148[4] 304[11])
    defparam i13933_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13545_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[6]), 
            .I3(\data_in_frame[14][6] ), .O(n29406));
    defparam i13545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13548_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60769), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29409));
    defparam i13548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13934_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n29795));   // verilog/coms.v(148[4] 304[11])
    defparam i13934_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1437 (.I0(n25700), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n61125));
    defparam i1_2_lut_adj_1437.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_adj_1438 (.I0(n55731), .I1(n10_adj_5601), .I2(n26147), 
            .I3(\data_out_frame[24] [2]), .O(n6_adj_5595));
    defparam i2_2_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_212_i3_3_lut_4_lut (.I0(n55523), .I1(n61207), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n61042), .O(n3_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_212_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n26181));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1440 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25604));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1440.LUT_INIT = 16'h6666;
    SB_LUT4 i13703_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29564));
    defparam i13703_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1441 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(GND_net), .I3(GND_net), .O(n61165));
    defparam i1_2_lut_adj_1441.LUT_INIT = 16'h6666;
    SB_LUT4 i13706_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29567));
    defparam i13706_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1442 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[3] [5]), .I3(n6_adj_5607), .O(n25683));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1443 (.I0(n23430), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[22] [5]), .I3(n55644), .O(n56541));
    defparam i1_2_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1444 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[11] [1]), 
            .I2(n61248), .I3(n6_adj_5615), .O(n25490));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1445 (.I0(n55715), .I1(n25490), .I2(GND_net), 
            .I3(GND_net), .O(n55761));
    defparam i1_2_lut_adj_1445.LUT_INIT = 16'h6666;
    SB_LUT4 i13709_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29570));
    defparam i13709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13712_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29573));
    defparam i13712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13715_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29576));
    defparam i13715_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13935_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n29796));   // verilog/coms.v(148[4] 304[11])
    defparam i13935_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1446 (.I0(\data_out_frame[17] [5]), .I1(\data_out_frame[15] [3]), 
            .I2(n61165), .I3(n55761), .O(n56728));
    defparam i1_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i18579_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n29797));   // verilog/coms.v(148[4] 304[11])
    defparam i18579_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1447 (.I0(n26181), .I1(n61125), .I2(n61012), 
            .I3(\data_in_frame[1] [4]), .O(n26621));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i13718_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29579));
    defparam i13718_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1448 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61144));
    defparam i1_2_lut_adj_1448.LUT_INIT = 16'h6666;
    SB_LUT4 i23_4_lut (.I0(\data_out_frame[17] [5]), .I1(n61150), .I2(\data_out_frame[17] [4]), 
            .I3(n61364), .O(n54));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(\data_out_frame[19] [3]), .I1(n56537), .I2(\data_out_frame[19] [7]), 
            .I3(n61424), .O(n52));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1449 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1449.LUT_INIT = 16'ha088;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[17] [7]), .I1(n60982), .I2(\data_out_frame[17] [6]), 
            .I3(\data_out_frame[16] [5]), .O(n53));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[18] [2]), .I3(\data_out_frame[12] [4]), 
            .O(n51));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1450 (.I0(n1516), .I1(n56537), .I2(n61213), 
            .I3(\data_out_frame[14] [3]), .O(n48));
    defparam i17_4_lut_adj_1450.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1451 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[19] [6]), 
            .I2(n61144), .I3(n56728), .O(n50_adj_5616));
    defparam i19_4_lut_adj_1451.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_71_i2_4_lut (.I0(\data_out_frame[8][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(n56127), .I1(\data_in_frame[10][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n60976));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h6666;
    SB_LUT4 i13937_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n29798));   // verilog/coms.v(148[4] 304[11])
    defparam i13937_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18_4_lut_adj_1453 (.I0(n1655), .I1(n56308), .I2(\data_out_frame[18] [7]), 
            .I3(n25604), .O(n49));
    defparam i18_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i13722_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29583));
    defparam i13722_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29_4_lut (.I0(n51), .I1(n53), .I2(n52), .I3(n54), .O(n60));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13725_3_lut_4_lut (.I0(n8_c), .I1(n60740), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29586));
    defparam i13725_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13938_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n29799));   // verilog/coms.v(148[4] 304[11])
    defparam i13938_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 equal_309_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5327));   // verilog/coms.v(157[7:23])
    defparam equal_309_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_308_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_c));   // verilog/coms.v(157[7:23])
    defparam equal_308_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 select_787_Select_70_i2_4_lut (.I0(\data_out_frame[8][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(n4_adj_5578), .I3(GND_net), .O(n61316));
    defparam i2_2_lut_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i24_4_lut_adj_1455 (.I0(n25490), .I1(n48), .I2(\data_out_frame[19] [5]), 
            .I3(n55741), .O(n55));
    defparam i24_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n55), .I1(n60), .I2(n49), .I3(n50_adj_5616), 
            .O(n61452));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_4_lut_adj_1456 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[15] [6]), .I3(\data_out_frame[15] [7]), 
            .O(n21_adj_5617));
    defparam i3_2_lut_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i13939_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n29800));   // verilog/coms.v(148[4] 304[11])
    defparam i13939_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13940_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n29801));   // verilog/coms.v(148[4] 304[11])
    defparam i13940_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1457 (.I0(\data_in_frame[9] [7]), .I1(n60976), 
            .I2(n26621), .I3(n25683), .O(n56591));
    defparam i3_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_69_i2_4_lut (.I0(\data_out_frame[8][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13409_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n29270));
    defparam i13409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13406_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n29267));
    defparam i13406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13941_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n29802));   // verilog/coms.v(148[4] 304[11])
    defparam i13941_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13403_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n29264));
    defparam i13403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1458 (.I0(n62686), .I1(n55517), .I2(GND_net), 
            .I3(GND_net), .O(n56531));
    defparam i1_2_lut_adj_1458.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_68_i2_4_lut (.I0(\data_out_frame[8][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_4_lut_adj_1459 (.I0(\data_out_frame[16] [2]), .I1(n60954), 
            .I2(\data_out_frame[19] [0]), .I3(n56531), .O(n12_adj_5618));
    defparam i5_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_67_i2_4_lut (.I0(\data_out_frame[8][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13400_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n29261));
    defparam i13400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1460 (.I0(n56573), .I1(n12_adj_5618), .I2(n61307), 
            .I3(n56624), .O(n55519));
    defparam i6_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_66_i2_4_lut (.I0(\data_out_frame[8][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13397_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n29258));
    defparam i13397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13394_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n29255));
    defparam i13394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1461 (.I0(\data_out_frame[20] [2]), .I1(n55499), 
            .I2(GND_net), .I3(GND_net), .O(n55650));
    defparam i1_2_lut_adj_1461.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(n62513), .I1(n55515), .I2(GND_net), 
            .I3(GND_net), .O(n56739));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h9999;
    SB_LUT4 i2_2_lut_4_lut_adj_1463 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[20] [5]), .I3(n55644), .O(n6_adj_5569));
    defparam i2_2_lut_4_lut_adj_1463.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13391_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n29252));
    defparam i13391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54976 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n72107));
    defparam byte_transmit_counter_0__bdd_4_lut_54976.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i4_4_lut_adj_1464 (.I0(\data_out_frame[22] [1]), .I1(n26289), 
            .I2(n26293), .I3(n6_adj_5604), .O(n56492));
    defparam i4_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1465 (.I0(\data_out_frame[20] [5]), .I1(n55644), 
            .I2(GND_net), .I3(GND_net), .O(n56578));
    defparam i1_2_lut_adj_1465.LUT_INIT = 16'h6666;
    SB_LUT4 n72107_bdd_4_lut (.I0(n72107), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n72110));
    defparam n72107_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60883));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13388_3_lut_4_lut (.I0(n8_c), .I1(n60769), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n29249));
    defparam i13388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13942_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n29803));   // verilog/coms.v(148[4] 304[11])
    defparam i13942_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1467 (.I0(n62824), .I1(n61089), .I2(n56739), 
            .I3(n23430), .O(n12_adj_5619));
    defparam i5_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_2_lut_3_lut_adj_1468 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n26405));
    defparam i2_2_lut_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1469 (.I0(\data_out_frame[22] [1]), .I1(n12_adj_5619), 
            .I2(n61349), .I3(n55499), .O(n55523));
    defparam i6_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(n1130), .I3(\data_out_frame[4] [6]), .O(n15_adj_5620));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n25461));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1471 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[7] [7]), .I3(\data_out_frame[5] [5]), .O(n61358));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1472 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(n26323), .I3(\data_out_frame[9] [4]), .O(n6_adj_5621));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1472.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(n55523), .I1(n61207), .I2(GND_net), 
            .I3(GND_net), .O(n56006));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_adj_1474 (.I0(\data_out_frame[24] [0]), .I1(n56675), 
            .I2(\data_out_frame[25] [7]), .I3(GND_net), .O(n60819));
    defparam i2_3_lut_adj_1474.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(n1168), .I3(\data_out_frame[6] [7]), .O(n61400));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n61015), .I3(n1191), .O(n1168));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1477 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[4] [7]), .O(n26323));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i27_2_lut (.I0(n23430), .I1(\data_out_frame[20] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n26293));   // verilog/coms.v(100[12:26])
    defparam i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1478 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n61015));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_3_lut_adj_1478.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1479 (.I0(n26293), .I1(n60819), .I2(n56006), 
            .I3(\data_out_frame[22] [4]), .O(n12_adj_5622));
    defparam i5_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i13943_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n29804));   // verilog/coms.v(148[4] 304[11])
    defparam i13943_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_209_i3_4_lut (.I0(n23471), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_5622), .I3(n8_adj_5623), .O(n3_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_209_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_2_lut_3_lut_adj_1480 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n6_adj_5624));   // verilog/coms.v(74[16:62])
    defparam i2_2_lut_3_lut_adj_1480.LUT_INIT = 16'h9696;
    SB_LUT4 i13944_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n29805));   // verilog/coms.v(148[4] 304[11])
    defparam i13944_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(n55525), .I1(n55715), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5625));
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1482 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[15] [2]), .I3(n6_adj_5625), .O(n62635));
    defparam i4_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1483 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[19] [1]), .I3(n61461), .O(n61195));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1484 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n61427));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1484.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1485 (.I0(n60912), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [7]), .I3(\data_out_frame[10] [4]), 
            .O(n14_adj_5626));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1486 (.I0(n37), .I1(\data_out_frame[13] [1]), .I2(n61239), 
            .I3(n25458), .O(n16_adj_5627));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i13945_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n29806));   // verilog/coms.v(148[4] 304[11])
    defparam i13945_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1487 (.I0(\data_out_frame[10] [5]), .I1(n26311), 
            .I2(n55572), .I3(\data_out_frame[10] [6]), .O(n13_adj_5628));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i13946_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n29807));   // verilog/coms.v(148[4] 304[11])
    defparam i13946_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13947_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n29808));   // verilog/coms.v(148[4] 304[11])
    defparam i13947_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11861_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27721));   // verilog/coms.v(109[34:55])
    defparam i11861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48321_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65411));
    defparam i48321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1488 (.I0(n13_adj_5628), .I1(n16_adj_5627), .I2(\data_out_frame[12] [7]), 
            .I3(n14_adj_5626), .O(n18_adj_5629));   // verilog/coms.v(75[16:27])
    defparam i8_4_lut_adj_1488.LUT_INIT = 16'h9669;
    SB_LUT4 i13948_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n29809));   // verilog/coms.v(148[4] 304[11])
    defparam i13948_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(n56545), .I1(n26038), .I2(\data_out_frame[10] [2]), 
            .I3(n31_adj_12), .O(n62886));
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i48322_4_lut (.I0(n65411), .I1(n27721), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n65412));
    defparam i48322_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i9_4_lut_adj_1490 (.I0(n62886), .I1(n18_adj_5629), .I2(n14_adj_5600), 
            .I3(n61394), .O(n55715));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut_adj_1490.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1491 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[8][4] ), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n60799));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1491.LUT_INIT = 16'h9696;
    SB_LUT4 i13949_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n29810));   // verilog/coms.v(148[4] 304[11])
    defparam i13949_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48320_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65410));
    defparam i48320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13950_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n29811));   // verilog/coms.v(148[4] 304[11])
    defparam i13950_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1492 (.I0(n56529), .I1(\data_in_frame[14][6] ), 
            .I2(\data_in_frame[17] [2]), .I3(n25825), .O(n18_adj_5631));
    defparam i7_4_lut_adj_1492.LUT_INIT = 16'h6996;
    SB_LUT4 i13951_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n29812));   // verilog/coms.v(148[4] 304[11])
    defparam i13951_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i3_4_lut_adj_1493 (.I0(n1130), .I1(n60799), .I2(n25461), .I3(\data_out_frame[13] [2]), 
            .O(n61406));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(n61242), .I1(n61406), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5632));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1495 (.I0(n55997), .I1(n18_adj_5631), .I2(n61276), 
            .I3(n60903), .O(n20_adj_5633));
    defparam i9_4_lut_adj_1495.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1496 (.I0(n25465), .I1(n26609), .I2(n61397), 
            .I3(n6_adj_5632), .O(n1720));
    defparam i4_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1497 (.I0(\data_in_frame[15] [1]), .I1(n61381), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5634));
    defparam i4_2_lut_adj_1497.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1498 (.I0(\data_out_frame[14] [2]), .I1(n26308), 
            .I2(n61288), .I3(\data_out_frame[11] [6]), .O(n13_adj_5635));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1499 (.I0(n13_adj_5635), .I1(n4_adj_5596), .I2(\data_out_frame[5] [4]), 
            .I3(\data_out_frame[5] [2]), .O(n55517));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1500 (.I0(\data_out_frame[10] [7]), .I1(n26136), 
            .I2(\data_out_frame[11] [2]), .I3(\data_out_frame[13] [3]), 
            .O(n61242));
    defparam i3_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1501 (.I0(n15_adj_5634), .I1(n20_adj_5633), .I2(n59626), 
            .I3(n61282), .O(n55970));
    defparam i10_4_lut_adj_1501.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1502 (.I0(n61242), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[8][6] ), .I3(n61400), .O(n10_adj_5636));   // verilog/coms.v(100[12:26])
    defparam i4_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1503 (.I0(\data_in_frame[12] [5]), .I1(n61276), 
            .I2(\data_in_frame[16] [7]), .I3(\data_in_frame[12] [3]), .O(n12_adj_5637));
    defparam i5_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1504 (.I0(n56308), .I1(n9_adj_5602), .I2(\data_out_frame[15] [5]), 
            .I3(n10_adj_5636), .O(n56537));
    defparam i2_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25528));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i13952_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n29813));   // verilog/coms.v(148[4] 304[11])
    defparam i13952_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1506 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60803));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1506.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1507 (.I0(n61279), .I1(\data_out_frame[4] [7]), 
            .I2(n60803), .I3(\data_out_frame[7] [0]), .O(n14_adj_5638));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1508 (.I0(\data_out_frame[11] [4]), .I1(n14_adj_5638), 
            .I2(n10_adj_5599), .I3(n26405), .O(n24849));   // verilog/coms.v(88[17:28])
    defparam i7_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(n24849), .I1(n61150), .I2(GND_net), 
            .I3(GND_net), .O(n60874));
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'h6666;
    SB_LUT4 i13953_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n29814));   // verilog/coms.v(148[4] 304[11])
    defparam i13953_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_out_frame[16] [0]), .I1(n56537), 
            .I2(GND_net), .I3(GND_net), .O(n61082));
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n60921));
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1512 (.I0(n60921), .I1(\data_out_frame[4] [7]), 
            .I2(\data_out_frame[6] [7]), .I3(n6_adj_5621), .O(n55368));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(n1168), .I1(n60864), .I2(GND_net), 
            .I3(GND_net), .O(n26136));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1514 (.I0(n26609), .I1(n25879), .I2(\data_out_frame[11] [4]), 
            .I3(n61264), .O(n10_adj_5597));
    defparam i4_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1515 (.I0(n61446), .I1(n61391), .I2(n62942), 
            .I3(n55517), .O(n56501));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[11] [5]), .I1(n55368), 
            .I2(GND_net), .I3(GND_net), .O(n55578));
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26457));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 i13954_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n29815));   // verilog/coms.v(148[4] 304[11])
    defparam i13954_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1518 (.I0(n60864), .I1(n26457), .I2(\data_out_frame[4] [7]), 
            .I3(n37), .O(n14_adj_5639));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i13955_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n29816));   // verilog/coms.v(148[4] 304[11])
    defparam i13955_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1519 (.I0(\data_out_frame[13] [4]), .I1(n14_adj_5639), 
            .I2(n10_adj_5640), .I3(\data_out_frame[9] [2]), .O(n56308));   // verilog/coms.v(88[17:70])
    defparam i7_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1520 (.I0(n61446), .I1(n61391), .I2(n62942), 
            .I3(n61452), .O(n61307));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1521 (.I0(n61147), .I1(\data_out_frame[13] [6]), 
            .I2(n56308), .I3(GND_net), .O(n61403));
    defparam i2_3_lut_adj_1521.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1522 (.I0(n61446), .I1(n61391), .I2(n62942), 
            .I3(\data_out_frame[17] [0]), .O(n61319));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1523 (.I0(\data_out_frame[16] [4]), .I1(n10_adj_5641), 
            .I2(n25712), .I3(n61319), .O(n61424));
    defparam i1_2_lut_4_lut_adj_1523.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1524 (.I0(\data_out_frame[16] [4]), .I1(n10_adj_5641), 
            .I2(n25712), .I3(n61442), .O(n61461));
    defparam i1_2_lut_4_lut_adj_1524.LUT_INIT = 16'h9669;
    SB_LUT4 i13956_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14][6] ), 
            .I3(deadband[22]), .O(n29817));   // verilog/coms.v(148[4] 304[11])
    defparam i13956_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61279));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h6666;
    SB_LUT4 i13957_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n29818));   // verilog/coms.v(148[4] 304[11])
    defparam i13957_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13958_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n29819));   // verilog/coms.v(148[4] 304[11])
    defparam i13958_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1526 (.I0(n25700), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[8][2] ), .I3(\data_in_frame[8] [1]), .O(n6_adj_5566));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1527 (.I0(n31_adj_12), .I1(n26308), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n60867));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i13959_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n29820));   // verilog/coms.v(148[4] 304[11])
    defparam i13959_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_adj_1528 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[7] [7]), 
            .I2(n61027), .I3(\data_in_frame[1]_c [5]), .O(n60779));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i392_2_lut (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1180));   // verilog/coms.v(77[16:27])
    defparam i392_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1529 (.I0(n26323), .I1(n1180), .I2(\data_out_frame[7] [4]), 
            .I3(\data_out_frame[9] [5]), .O(n31_adj_12));
    defparam i3_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1530 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[7] [6]), 
            .I2(n6_adj_5624), .I3(n26311), .O(n4_adj_5596));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26038));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1532 (.I0(\data_out_frame[14] [3]), .I1(n61391), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n61003));
    defparam i2_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i13960_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n29821));   // verilog/coms.v(148[4] 304[11])
    defparam i13960_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_65_i2_4_lut (.I0(\data_out_frame[8][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1533 (.I0(n55741), .I1(\data_out_frame[7] [6]), 
            .I2(n26038), .I3(n6_adj_5594), .O(n56573));
    defparam i4_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1534 (.I0(n60867), .I1(n61236), .I2(n61003), 
            .I3(n60877), .O(n63014));
    defparam i3_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1535 (.I0(n63014), .I1(n61449), .I2(n61245), 
            .I3(n61403), .O(n10_adj_5642));
    defparam i4_4_lut_adj_1535.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1536 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [0]), .I3(n26457), .O(n63376));
    defparam i3_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1537 (.I0(\data_out_frame[11] [7]), .I1(n60782), 
            .I2(\data_out_frame[10] [7]), .I3(n1244), .O(n63283));
    defparam i3_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i13961_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n29822));   // verilog/coms.v(148[4] 304[11])
    defparam i13961_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i10_4_lut_adj_1538 (.I0(n61082), .I1(\data_out_frame[13] [5]), 
            .I2(n26691), .I3(n60874), .O(n28_c));
    defparam i10_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54882 (.I0(byte_transmit_counter[1]), 
            .I1(n65341), .I2(n65342), .I3(byte_transmit_counter[2]), .O(n71957));
    defparam byte_transmit_counter_1__bdd_4_lut_54882.LUT_INIT = 16'he4aa;
    SB_LUT4 i13_4_lut (.I0(n63283), .I1(n55368), .I2(\data_out_frame[12] [7]), 
            .I3(\data_out_frame[13] [7]), .O(n31_adj_5643));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1539 (.I0(\data_out_frame[15] [2]), .I1(n26691), 
            .I2(n10_adj_5642), .I3(\data_out_frame[14] [6]), .O(n22_adj_5644));
    defparam i4_4_lut_adj_1539.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1540 (.I0(n55517), .I1(n1720), .I2(n63376), 
            .I3(\data_out_frame[14] [1]), .O(n30));
    defparam i12_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i13962_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n29823));   // verilog/coms.v(148[4] 304[11])
    defparam i13962_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut_adj_1541 (.I0(n31_adj_5643), .I1(n55715), .I2(n28_c), 
            .I3(n4_adj_5578), .O(n34_adj_5645));
    defparam i16_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1542 (.I0(\data_in_frame[14] [5]), .I1(n12_adj_5637), 
            .I2(\data_in_frame[17] [1]), .I3(n56591), .O(n61039));
    defparam i6_4_lut_adj_1542.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1543 (.I0(\data_out_frame[9] [4]), .I1(n26323), 
            .I2(n25879), .I3(GND_net), .O(n26308));
    defparam i1_2_lut_3_lut_adj_1543.LUT_INIT = 16'h9696;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(n21_adj_5617), .I1(n34_adj_5645), .I2(n30), 
            .I3(n22_adj_5644), .O(n25994));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1545 (.I0(n25994), .I1(n26691), .I2(n56573), 
            .I3(\data_out_frame[16] [6]), .O(n10_adj_5641));
    defparam i4_4_lut_adj_1545.LUT_INIT = 16'h6996;
    SB_LUT4 i13963_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n29824));   // verilog/coms.v(148[4] 304[11])
    defparam i13963_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13964_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n29825));   // verilog/coms.v(148[4] 304[11])
    defparam i13964_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1546 (.I0(\data_out_frame[16] [5]), .I1(n61006), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n25712));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(reset), .I3(GND_net), .O(n22465));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_1547 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n60864));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i13965_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n29826));   // verilog/coms.v(148[4] 304[11])
    defparam i13965_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13966_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n29827));   // verilog/coms.v(148[4] 304[11])
    defparam i13966_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13967_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n29828));   // verilog/coms.v(148[4] 304[11])
    defparam i13967_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1548 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[19] [1]), .I3(n61006), .O(n15_adj_5646));
    defparam i6_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1549 (.I0(n15_adj_5646), .I1(n26555), .I2(n14_adj_5593), 
            .I3(n61424), .O(n26560));
    defparam i8_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1550 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [0]), 
            .I2(n61406), .I3(GND_net), .O(n6_adj_5615));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1550.LUT_INIT = 16'h9696;
    SB_LUT4 n71957_bdd_4_lut (.I0(n71957), .I1(n65435), .I2(n65434), .I3(byte_transmit_counter[2]), 
            .O(n71960));
    defparam n71957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1551 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25874));
    defparam i1_2_lut_adj_1551.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut_adj_1552 (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n10_adj_5640));   // verilog/coms.v(88[17:70])
    defparam i2_2_lut_3_lut_adj_1552.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1553 (.I0(\data_out_frame[16] [1]), .I1(n61195), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n60954));
    defparam i2_3_lut_adj_1553.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1554 (.I0(n55595), .I1(n60954), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5647));
    defparam i1_2_lut_adj_1554.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1555 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n61403), .I3(GND_net), .O(n6_adj_5605));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1555.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1556 (.I0(\data_out_frame[21] [3]), .I1(n25874), 
            .I2(\data_out_frame[17] [1]), .I3(n6_adj_5647), .O(n55598));
    defparam i4_4_lut_adj_1556.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1557 (.I0(\data_out_frame[21] [2]), .I1(n26560), 
            .I2(GND_net), .I3(GND_net), .O(n55639));
    defparam i1_2_lut_adj_1557.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1558 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(n28), .I3(\data_out_frame[12] [2]), .O(n61391));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1559 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n61236));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1559.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1560 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[10] [0]), 
            .I2(n60796), .I3(n61236), .O(n62942));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1560.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1561 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n61449));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1561.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n60666));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61446));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1563 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n60912));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1563.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1564 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5649));   // verilog/coms.v(88[17:70])
    defparam i2_2_lut_adj_1564.LUT_INIT = 16'h6666;
    SB_LUT4 i13968_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n29829));   // verilog/coms.v(148[4] 304[11])
    defparam i13968_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i6_4_lut_adj_1565 (.I0(\data_out_frame[8][1] ), .I1(n61446), 
            .I2(n61355), .I3(n61153), .O(n14_adj_5650));   // verilog/coms.v(88[17:70])
    defparam i6_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1566 (.I0(\data_out_frame[12] [4]), .I1(n14_adj_5650), 
            .I2(n10_adj_5649), .I3(n60912), .O(n1655));   // verilog/coms.v(88[17:70])
    defparam i7_4_lut_adj_1566.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1567 (.I0(n1244), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[4] [0]), .O(n61239));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i13969_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n29830));   // verilog/coms.v(148[4] 304[11])
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i5_4_lut_adj_1568 (.I0(\data_out_frame[12] [6]), .I1(n61358), 
            .I2(n61239), .I3(\data_out_frame[10] [5]), .O(n12_adj_5651));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1568.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1569 (.I0(n60806), .I1(n12_adj_5651), .I2(n61449), 
            .I3(\data_out_frame[8][1] ), .O(n55525));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_1569.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1570 (.I0(\data_out_frame[14] [5]), .I1(n1655), 
            .I2(GND_net), .I3(GND_net), .O(n26691));
    defparam i1_2_lut_adj_1570.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1571 (.I0(n61039), .I1(\data_in_frame[19] [3]), 
            .I2(n55970), .I3(GND_net), .O(n63420));
    defparam i2_3_lut_adj_1571.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1572 (.I0(\data_out_frame[8][1] ), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60796));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1572.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1573 (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n61355));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1574 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60844));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1574.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1575 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[6] [0]), .O(n62822));   // verilog/coms.v(88[17:70])
    defparam i3_4_lut_adj_1575.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61110));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1577 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n61394));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1577.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54842 (.I0(byte_transmit_counter[1]), 
            .I1(n65464), .I2(n65465), .I3(byte_transmit_counter[2]), .O(n71951));
    defparam byte_transmit_counter_1__bdd_4_lut_54842.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1578 (.I0(n61394), .I1(\data_out_frame[12] [5]), 
            .I2(n61110), .I3(\data_out_frame[12] [4]), .O(n14_adj_5652));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i13970_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n29831));   // verilog/coms.v(148[4] 304[11])
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i7_4_lut_adj_1579 (.I0(\data_out_frame[14] [6]), .I1(n14_adj_5652), 
            .I2(n10_adj_5591), .I3(n60796), .O(n26555));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1579.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1580 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60982));
    defparam i1_2_lut_adj_1580.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1581 (.I0(\data_out_frame[15] [0]), .I1(n26691), 
            .I2(n55525), .I3(\data_out_frame[16] [7]), .O(n55595));
    defparam i3_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(n56545), .I1(n26215), .I2(GND_net), 
            .I3(GND_net), .O(n55572));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n60924));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1584 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n60850));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1584.LUT_INIT = 16'h9696;
    SB_LUT4 n71951_bdd_4_lut (.I0(n71951), .I1(n65453), .I2(n65452), .I3(byte_transmit_counter[2]), 
            .O(n71954));
    defparam n71951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1585 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n61264));
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1586 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n55519), .I3(GND_net), .O(n61024));
    defparam i1_2_lut_3_lut_adj_1586.LUT_INIT = 16'h9696;
    SB_LUT4 i13971_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n29832));   // verilog/coms.v(148[4] 304[11])
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61397));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1588 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n61153));
    defparam i1_2_lut_adj_1588.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1589 (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[8][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n61248));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1589.LUT_INIT = 16'h6666;
    SB_LUT4 i13972_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n29833));   // verilog/coms.v(148[4] 304[11])
    defparam i13972_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1590 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(\data_out_frame[18] [6]), .I3(\data_out_frame[16] [5]), 
            .O(n6));
    defparam i1_2_lut_3_lut_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i13973_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n29834));   // verilog/coms.v(148[4] 304[11])
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(\data_out_frame[6] [6]), .I1(n61400), 
            .I2(GND_net), .I3(GND_net), .O(n26609));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'h6666;
    SB_LUT4 i44537_3_lut_4_lut (.I0(n10_adj_5567), .I1(n39431), .I2(n8), 
            .I3(reset), .O(n28096));
    defparam i44537_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i13974_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n29835));   // verilog/coms.v(148[4] 304[11])
    defparam i13974_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i12241_3_lut_4_lut (.I0(n10_adj_5567), .I1(n39431), .I2(reset), 
            .I3(n8_adj_5437), .O(n28102));
    defparam i12241_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i13975_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n29836));   // verilog/coms.v(148[4] 304[11])
    defparam i13975_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(\data_out_frame[6] [1]), .I1(n25461), 
            .I2(GND_net), .I3(GND_net), .O(n25458));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1593 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[4] [6]), .I3(n63330), .O(n12_adj_5654));   // verilog/coms.v(169[9:87])
    defparam i5_4_lut_adj_1593.LUT_INIT = 16'h6996;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13976_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n29837));   // verilog/coms.v(148[4] 304[11])
    defparam i13976_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_adj_1594 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8][1] ), 
            .I2(\data_out_frame[8][4] ), .I3(GND_net), .O(n60782));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1594.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1595 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n60877));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1595.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1596 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61000));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1596.LUT_INIT = 16'h6666;
    SB_LUT4 i52191_2_lut (.I0(n72098), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n68453));
    defparam i52191_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13308_3_lut (.I0(\data_in_frame[10]_c [0]), .I1(rx_data[0]), 
            .I2(n60771), .I3(GND_net), .O(n29169));   // verilog/coms.v(130[12] 305[6])
    defparam i13308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53609_3_lut (.I0(n72182), .I1(n71900), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70699));
    defparam i53609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1597 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(\FRAME_MATCHER.i [0]), .O(n37941));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1597.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1598 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[7] [2]), .I3(n60877), .O(n19_adj_5655));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54857 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n71945));
    defparam byte_transmit_counter_0__bdd_4_lut_54857.LUT_INIT = 16'he4aa;
    SB_LUT4 i11966_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n27827));   // verilog/coms.v(109[34:55])
    defparam i11966_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1599 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n60760), .I3(\FRAME_MATCHER.i [0]), .O(n60766));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1599.LUT_INIT = 16'hfffd;
    SB_LUT4 i48324_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65414));
    defparam i48324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1600 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n60769), .I3(\FRAME_MATCHER.i [0]), .O(n60771));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1600.LUT_INIT = 16'hfffd;
    SB_LUT4 i48325_4_lut (.I0(n65414), .I1(n27827), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n65415));
    defparam i48325_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i48323_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65413));
    defparam i48323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12749_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(LED_c), .I3(n63143), 
            .O(n28610));   // verilog/coms.v(130[12] 305[6])
    defparam i12749_4_lut_4_lut.LUT_INIT = 16'h5444;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1601 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n3483), .I3(\FRAME_MATCHER.i [0]), .O(n8_adj_13));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1601.LUT_INIT = 16'h0020;
    SB_LUT4 i2_2_lut_4_lut_adj_1602 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n32327), .O(n6_adj_5565));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_310_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_5437));   // verilog/coms.v(157[7:23])
    defparam equal_310_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i10_4_lut_adj_1603 (.I0(n19_adj_5655), .I1(n15_adj_5620), .I2(n26609), 
            .I3(n61000), .O(n22_adj_5657));   // verilog/coms.v(77[16:43])
    defparam i10_4_lut_adj_1603.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1604 (.I0(\data_out_frame[6] [4]), .I1(n22_adj_5657), 
            .I2(n18_adj_5581), .I3(\data_out_frame[4] [5]), .O(n63172));   // verilog/coms.v(77[16:43])
    defparam i11_4_lut_adj_1604.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1605 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[7] [0]), 
            .I2(n60782), .I3(n63172), .O(n16_adj_5658));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1605.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1606 (.I0(n61248), .I1(n61409), .I2(\data_out_frame[7] [3]), 
            .I3(n61015), .O(n17_adj_5659));   // verilog/coms.v(77[16:43])
    defparam i7_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i12742_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28603));   // verilog/coms.v(130[12] 305[6])
    defparam i12742_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i6_4_lut_adj_1607 (.I0(n26215), .I1(\data_out_frame[9] [4]), 
            .I2(n61264), .I3(\data_out_frame[9] [5]), .O(n14_adj_5660));
    defparam i6_4_lut_adj_1607.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1608 (.I0(n17_adj_5659), .I1(\data_out_frame[7] [1]), 
            .I2(n16_adj_5658), .I3(\data_out_frame[7] [7]), .O(n63189));   // verilog/coms.v(77[16:43])
    defparam i9_4_lut_adj_1608.LUT_INIT = 16'h6996;
    SB_LUT4 equal_306_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_5567));   // verilog/coms.v(158[12:15])
    defparam equal_306_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1609 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n115), .O(n60760));   // verilog/coms.v(158[12:15])
    defparam i2_3_lut_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1610 (.I0(n63189), .I1(n14_adj_5660), .I2(n10_adj_5579), 
            .I3(n61153), .O(n56545));
    defparam i7_4_lut_adj_1610.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1611 (.I0(\data_out_frame[17] [6]), .I1(n56308), 
            .I2(n25528), .I3(n10_adj_5613), .O(n26289));
    defparam i5_3_lut_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54966 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n72101));
    defparam byte_transmit_counter_0__bdd_4_lut_54966.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1612 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n12_adj_5661));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1612.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_adj_1613 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[8][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n61409));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1613.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1614 (.I0(n60825), .I1(n12_adj_5654), .I2(\data_in_frame[5] [0]), 
            .I3(\data_in_frame[2] [6]), .O(n26250));   // verilog/coms.v(169[9:87])
    defparam i6_4_lut_adj_1614.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1615 (.I0(\data_out_frame[17] [6]), .I1(n56308), 
            .I2(n61162), .I3(n10_adj_5614), .O(n55499));
    defparam i5_3_lut_4_lut_adj_1615.LUT_INIT = 16'h6996;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1616 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(n62914), .I3(n23430), .O(n56553));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut_adj_1616.LUT_INIT = 16'h9669;
    SB_LUT4 n71945_bdd_4_lut (.I0(n71945), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n71948));
    defparam n71945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n72101_bdd_4_lut (.I0(n72101), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n72104));
    defparam n72101_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1617 (.I0(n1191), .I1(n61409), .I2(\data_out_frame[8][4] ), 
            .I3(GND_net), .O(n60806));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1617.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1618 (.I0(n60806), .I1(\data_out_frame[10] [4]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[12] [6]), .O(n14_adj_5662));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1619 (.I0(n61245), .I1(n56545), .I2(n25465), 
            .I3(\data_out_frame[12] [7]), .O(n13_adj_5663));   // verilog/coms.v(88[17:28])
    defparam i5_4_lut_adj_1619.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1620 (.I0(n13_adj_5663), .I1(\data_out_frame[13] [0]), 
            .I2(n14_adj_5662), .I3(GND_net), .O(n4_adj_5578));
    defparam i1_3_lut_adj_1620.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1621 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n61009));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1621.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1622 (.I0(n55631), .I1(n61159), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n55644));
    defparam i1_2_lut_3_lut_adj_1622.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54961 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n72095));
    defparam byte_transmit_counter_0__bdd_4_lut_54961.LUT_INIT = 16'he4aa;
    SB_LUT4 i13977_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n29838));   // verilog/coms.v(148[4] 304[11])
    defparam i13977_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1623 (.I0(n55631), .I1(n61159), .I2(n55893), 
            .I3(GND_net), .O(n61349));
    defparam i1_2_lut_3_lut_adj_1623.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1624 (.I0(\data_out_frame[21] [6]), .I1(n61418), 
            .I2(\data_out_frame[21] [7]), .I3(\data_out_frame[24] [0]), 
            .O(n8_adj_5598));
    defparam i3_3_lut_4_lut_adj_1624.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1625 (.I0(\data_out_frame[21] [6]), .I1(n61418), 
            .I2(n55731), .I3(GND_net), .O(n61089));
    defparam i1_2_lut_3_lut_adj_1625.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1626 (.I0(n55595), .I1(n61316), .I2(n60982), 
            .I3(n26555), .O(n62642));
    defparam i3_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1627 (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(n32330), .I3(GND_net), .O(n5_adj_5547));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1627.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_adj_1628 (.I0(n62642), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[19] [3]), .I3(GND_net), .O(n61291));
    defparam i2_3_lut_adj_1628.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1629 (.I0(n61156), .I1(n61427), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5664));
    defparam i1_2_lut_adj_1629.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1630 (.I0(\data_out_frame[22] [3]), .I1(n26289), 
            .I2(\data_out_frame[24] [4]), .I3(n55650), .O(n56543));
    defparam i2_3_lut_4_lut_adj_1630.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1631 (.I0(\data_out_frame[21] [4]), .I1(\data_out_frame[19] [3]), 
            .I2(n61319), .I3(n6_adj_5664), .O(n56632));
    defparam i4_4_lut_adj_1631.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1632 (.I0(n56632), .I1(n61421), .I2(GND_net), 
            .I3(GND_net), .O(n61181));
    defparam i1_2_lut_adj_1632.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1633 (.I0(\data_out_frame[19] [4]), .I1(n62635), 
            .I2(n61156), .I3(n26555), .O(n55731));
    defparam i3_4_lut_adj_1633.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1634 (.I0(\data_out_frame[22] [3]), .I1(n26289), 
            .I2(n56553), .I3(GND_net), .O(n8_adj_5623));
    defparam i1_2_lut_3_lut_adj_1634.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(\data_out_frame[25] [7]), .I1(n55731), .I2(n61251), 
            .I3(GND_net), .O(n8_adj_5665));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1087_i18_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n4939[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_208_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5665), .I3(n61181), 
            .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_adj_1635 (.I0(\data_in_frame[0] [2]), .I1(ID[4]), .I2(ID[2]), 
            .I3(\data_in_frame[0] [4]), .O(n10_adj_5666));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1635.LUT_INIT = 16'h7bde;
    SB_LUT4 select_787_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1636 (.I0(\data_out_frame[24] [5]), .I1(n56553), 
            .I2(\data_out_frame[25] [0]), .I3(GND_net), .O(n6_adj_5592));
    defparam i2_2_lut_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i12738_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28599));   // verilog/coms.v(130[12] 305[6])
    defparam i12738_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_787_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1637 (.I0(\data_out_frame[24] [5]), .I1(n56553), 
            .I2(n56543), .I3(\FRAME_MATCHER.state[3] ), .O(n3_adj_5395));
    defparam i1_3_lut_4_lut_adj_1637.LUT_INIT = 16'h9600;
    SB_LUT4 i54642_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n39534), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i54642_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 select_787_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1638 (.I0(\data_in_frame[9] [3]), .I1(n60944), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n25765));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1638.LUT_INIT = 16'h9696;
    SB_LUT4 i21704_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1]_c [0]), 
            .I2(n22465), .I3(GND_net), .O(n29109));
    defparam i21704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1639 (.I0(n56127), .I1(Kp_23__N_1080), .I2(n26258), 
            .I3(GND_net), .O(n56581));
    defparam i1_2_lut_3_lut_adj_1639.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1640 (.I0(n55580), .I1(n56075), .I2(n25765), 
            .I3(GND_net), .O(n55511));
    defparam i1_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1641 (.I0(n25746), .I1(n25765), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n25781));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1641.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1087_i19_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1][2] ), .I3(\data_in_frame[17] [2]), .O(n4939[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i19_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i54478_2_lut_3_lut (.I0(n23700), .I1(n23704), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n71568));   // verilog/coms.v(99[12:25])
    defparam i54478_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_198_i2_4_lut (.I0(\data_out_frame[24] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_198_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [5]), 
            .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1087_i20_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1]_c [3]), .I3(\data_in_frame[17] [3]), .O(n4939[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i21_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n4939[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_4_lut_adj_1643 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [4]), 
            .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1643.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1644 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n61119));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1644.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1645 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(ID[6]), .I3(ID[1]), .O(n11_adj_5667));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1645.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_4_lut_adj_1646 (.I0(\data_in_frame[10]_c [0]), .I1(\data_in_frame[9] [6]), 
            .I2(n26262), .I3(\data_in_frame[9] [7]), .O(n25614));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1646.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1647 (.I0(n26057), .I1(\data_in_frame[9] [7]), 
            .I2(n10_adj_5556), .I3(n26258), .O(n61201));
    defparam i5_3_lut_4_lut_adj_1647.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_adj_1648 (.I0(n25781), .I1(n55511), .I2(\data_in_frame[14] [7]), 
            .I3(GND_net), .O(n61381));
    defparam i1_3_lut_adj_1648.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1649 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[4] [2]), .O(n60993));   // verilog/coms.v(76[16:42])
    defparam i1_3_lut_4_lut_adj_1649.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1650 (.I0(n61039), .I1(\data_in_frame[19] [3]), 
            .I2(n55970), .I3(n61062), .O(n55617));
    defparam i1_2_lut_4_lut_adj_1650.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1651 (.I0(n55970), .I1(\data_in_frame[19] [4]), 
            .I2(n62964), .I3(GND_net), .O(n55682));
    defparam i2_3_lut_adj_1651.LUT_INIT = 16'h6969;
    SB_LUT4 mux_1087_i22_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1]_c [5]), .I3(\data_in_frame[17] [5]), .O(n4939[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[16] [5]), 
            .I2(n61185), .I3(GND_net), .O(n61224));
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i23_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1][6] ), .I3(\data_in_frame[17] [6]), .O(n4939[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i13_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n4939[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i14_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n4939[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i15_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n4939[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5668));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'h7bde;
    SB_LUT4 mux_1087_i17_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1]_c [0]), .I3(\data_in_frame[17] [0]), .O(n4939[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54837 (.I0(byte_transmit_counter[1]), 
            .I1(n65392), .I2(n65393), .I3(byte_transmit_counter[2]), .O(n71933));
    defparam byte_transmit_counter_1__bdd_4_lut_54837.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1654 (.I0(n9_adj_5668), .I1(n11_adj_5667), .I2(n10_adj_5666), 
            .I3(n12_adj_5661), .O(n55137));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [4]), 
            .I2(\control_mode[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n8_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode_c[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(n61198), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n64955));
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'h6666;
    SB_LUT4 n71933_bdd_4_lut (.I0(n71933), .I1(n65426), .I2(n65425), .I3(byte_transmit_counter[2]), 
            .O(n71936));
    defparam n71933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\control_mode[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1657 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n26154));   // verilog/coms.v(169[9:87])
    defparam i2_3_lut_adj_1657.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1658 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n25591));   // verilog/coms.v(169[9:87])
    defparam i1_3_lut_adj_1658.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [0]), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'ha088;
    SB_LUT4 i51695_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68365));   // verilog/coms.v(158[12:15])
    defparam i51695_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48218_3_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65308));
    defparam i48218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48219_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65309));
    defparam i48219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48534_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65624));
    defparam i48534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48533_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65623));
    defparam i48533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51694_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68364));   // verilog/coms.v(158[12:15])
    defparam i51694_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1660 (.I0(n56535), .I1(n61381), .I2(n56505), 
            .I3(n64955), .O(n62964));
    defparam i1_4_lut_adj_1660.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1661 (.I0(n26220), .I1(n4_c), .I2(\data_in_frame[8][7] ), 
            .I3(\data_in_frame[8][6] ), .O(n64765));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i16_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n4939[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i6_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n4939[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i5_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n4939[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i5_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i4_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n4939[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i11859_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27719));   // verilog/coms.v(109[34:55])
    defparam i11859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48315_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65405));
    defparam i48315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48316_4_lut (.I0(n65405), .I1(n27719), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n65406));
    defparam i48316_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i48314_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n65404));
    defparam i48314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54822 (.I0(byte_transmit_counter[1]), 
            .I1(n65437), .I2(n65438), .I3(byte_transmit_counter[2]), .O(n71927));
    defparam byte_transmit_counter_1__bdd_4_lut_54822.LUT_INIT = 16'he4aa;
    SB_LUT4 n71927_bdd_4_lut (.I0(n71927), .I1(n65390), .I2(n65389), .I3(byte_transmit_counter[2]), 
            .O(n71930));
    defparam n71927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1662 (.I0(n62964), .I1(n62519), .I2(n55682), 
            .I3(\data_in_frame[19] [5]), .O(n63317));
    defparam i3_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1663 (.I0(n61216), .I1(n61385), .I2(n55639), 
            .I3(n63365), .O(n61233));
    defparam i1_2_lut_4_lut_adj_1663.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_4_lut_adj_1664 (.I0(n61216), .I1(n61385), .I2(n55639), 
            .I3(n61251), .O(n6_adj_5435));
    defparam i2_2_lut_4_lut_adj_1664.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i3_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n4939[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i3_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 n72095_bdd_4_lut (.I0(n72095), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n72098));
    defparam n72095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_54817 (.I0(byte_transmit_counter[1]), 
            .I1(n65455), .I2(n65456), .I3(byte_transmit_counter[2]), .O(n71921));
    defparam byte_transmit_counter_1__bdd_4_lut_54817.LUT_INIT = 16'he4aa;
    SB_LUT4 n71921_bdd_4_lut (.I0(n71921), .I1(n65384), .I2(n65383), .I3(byte_transmit_counter[2]), 
            .O(n71924));
    defparam n71921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1665 (.I0(n63420), .I1(\data_in_frame[21] [5]), 
            .I2(n55682), .I3(GND_net), .O(n61116));
    defparam i2_3_lut_adj_1665.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54956 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n72089));
    defparam byte_transmit_counter_0__bdd_4_lut_54956.LUT_INIT = 16'he4aa;
    SB_LUT4 n72089_bdd_4_lut (.I0(n72089), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n72092));
    defparam n72089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1666 (.I0(\data_in_frame[8][6] ), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8][7] ), .I3(\data_in_frame[11] [3]), .O(n64921));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1666.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1087_i2_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n4939[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i2_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i1_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n4939[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i24_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n4939[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i9_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n4939[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut_adj_1667 (.I0(\data_in_frame[21] [6]), .I1(n61116), 
            .I2(n63317), .I3(GND_net), .O(n60966));
    defparam i2_3_lut_adj_1667.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1087_i10_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n4939[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i11_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n4939[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i12_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n4939[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i1_3_lut_adj_1668 (.I0(\data_in_frame[1][2] ), .I1(\data_in_frame[1]_c [3]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n25700));   // verilog/coms.v(79[16:43])
    defparam i1_3_lut_adj_1668.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1087_i8_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n4939[7]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i7_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n33_adj_5555), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n4939[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54951 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n72083));
    defparam byte_transmit_counter_0__bdd_4_lut_54951.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1669 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n61070));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1669.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1670 (.I0(n25700), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n61036));
    defparam i1_2_lut_adj_1670.LUT_INIT = 16'h6666;
    SB_LUT4 i13653_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29514));
    defparam i13653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13656_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29517));
    defparam i13656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1671 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25260), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n64994));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1671.LUT_INIT = 16'hfff4;
    SB_LUT4 i1_2_lut_adj_1672 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61092));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1672.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(Kp_23__N_799), .I1(n61455), .I2(n61018), 
            .I3(n64693), .O(n56614));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1674 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[0] [7]), 
            .I2(n61036), .I3(n25687), .O(n61027));
    defparam i3_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1675 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n61055));
    defparam i1_2_lut_adj_1675.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1676 (.I0(n25540), .I1(\data_in_frame[7] [6]), 
            .I2(n25700), .I3(GND_net), .O(n23704));
    defparam i2_3_lut_adj_1676.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1677 (.I0(n25683), .I1(n60841), .I2(GND_net), 
            .I3(GND_net), .O(n55700));
    defparam i1_2_lut_adj_1677.LUT_INIT = 16'h6666;
    SB_LUT4 i13660_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29521));
    defparam i13660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13663_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29524));
    defparam i13663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n72083_bdd_4_lut (.I0(n72083), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n72086));
    defparam n72083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13666_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29527));
    defparam i13666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1678 (.I0(n61027), .I1(n56614), .I2(GND_net), 
            .I3(GND_net), .O(n56707));
    defparam i1_2_lut_adj_1678.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1679 (.I0(n25700), .I1(\data_in_frame[3] [3]), 
            .I2(n60993), .I3(GND_net), .O(n64663));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 i13669_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29530));
    defparam i13669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1680 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [3]), 
            .I2(n25614), .I3(GND_net), .O(n61141));
    defparam i2_3_lut_adj_1680.LUT_INIT = 16'h9696;
    SB_LUT4 i53627_3_lut (.I0(n72122), .I1(n71906), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n70717));
    defparam i53627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13672_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29533));
    defparam i13672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13675_3_lut_4_lut (.I0(n8_adj_5437), .I1(n60740), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29536));
    defparam i13675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1681 (.I0(\data_in_frame[0] [3]), .I1(n61092), 
            .I2(n61070), .I3(n60844), .O(Kp_23__N_748));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1681.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1682 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[10][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n64947));
    defparam i1_2_lut_adj_1682.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1683 (.I0(n56563), .I1(\data_in_frame[16] [4]), 
            .I2(n56696), .I3(\data_in_frame[16] [5]), .O(n63034));
    defparam i2_3_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n56707), .I1(n55700), .I2(n23704), 
            .I3(n64947), .O(n56634));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54946 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n72077));
    defparam byte_transmit_counter_0__bdd_4_lut_54946.LUT_INIT = 16'he4aa;
    SB_LUT4 n72077_bdd_4_lut (.I0(n72077), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n72080));
    defparam n72077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i9_4_lut_adj_1685 (.I0(n25598), .I1(\data_in_frame[1] [4]), 
            .I2(Kp_23__N_748), .I3(\data_in_frame[2] [1]), .O(n26_adj_5669));
    defparam i9_4_lut_adj_1685.LUT_INIT = 16'h0440;
    SB_LUT4 select_787_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1686 (.I0(n56634), .I1(n61141), .I2(\data_in_frame[14] [4]), 
            .I3(GND_net), .O(n56696));
    defparam i2_3_lut_adj_1686.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1687 (.I0(n25825), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[12] [4]), .I3(n56634), .O(n56640));
    defparam i2_3_lut_4_lut_adj_1687.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1688 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1]_c [0]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[0] [6]), .O(n24));
    defparam i7_4_lut_adj_1688.LUT_INIT = 16'h8124;
    SB_LUT4 i1_2_lut_4_lut_adj_1689 (.I0(n61439), .I1(\data_in_frame[16] [3]), 
            .I2(n62654), .I3(n26198), .O(n61174));
    defparam i1_2_lut_4_lut_adj_1689.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1690 (.I0(n55617), .I1(\data_in_frame[21] [4]), 
            .I2(n61116), .I3(\data_in_frame[23] [6]), .O(n63036));
    defparam i2_3_lut_4_lut_adj_1690.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1691 (.I0(\data_in_frame[18] [2]), .I1(n56678), 
            .I2(n10_adj_5450), .I3(\data_in_frame[13] [4]), .O(n6_adj_5544));
    defparam i1_2_lut_4_lut_adj_1691.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1692 (.I0(n25825), .I1(\data_in_frame[12] [5]), 
            .I2(n26274), .I3(GND_net), .O(n25817));
    defparam i1_2_lut_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i13879_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [7]), 
            .I3(neopxl_color[23]), .O(n29740));   // verilog/coms.v(130[12] 305[6])
    defparam i13879_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_4_lut_adj_1693 (.I0(n56684), .I1(n56563), .I2(\data_in_frame[16] [3]), 
            .I3(n25950), .O(n56575));
    defparam i1_2_lut_4_lut_adj_1693.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1694 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(n24953), .O(n61198));
    defparam i1_2_lut_4_lut_adj_1694.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1695 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n24953), .I3(GND_net), .O(n55550));
    defparam i1_2_lut_3_lut_adj_1695.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_4_lut_adj_1696 (.I0(n26089), .I1(n26250), .I2(\data_in_frame[9] [2]), 
            .I3(n56614), .O(n10_adj_5448));
    defparam i2_2_lut_4_lut_adj_1696.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_in_frame[10]_c [0]), .I1(\data_in_frame[9] [6]), 
            .I2(n71568), .I3(\data_in_frame[9] [3]), .O(n10_adj_5446));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1697 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_974), .I3(GND_net), .O(n25556));
    defparam i1_2_lut_3_lut_adj_1697.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1698 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [3]), 
            .I2(n61092), .I3(\data_in_frame[2] [1]), .O(n60880));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut_adj_1698.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54941 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n72071));
    defparam byte_transmit_counter_0__bdd_4_lut_54941.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54800 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[1]), .O(n71897));
    defparam byte_transmit_counter_0__bdd_4_lut_54800.LUT_INIT = 16'he4aa;
    SB_LUT4 n71897_bdd_4_lut (.I0(n71897), .I1(\data_out_frame[21] [7]), 
            .I2(\data_out_frame[20] [7]), .I3(byte_transmit_counter[1]), 
            .O(n71900));
    defparam n71897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1699 (.I0(n59688), .I1(n56561), .I2(\data_in_frame[19] [0]), 
            .I3(GND_net), .O(n61310));
    defparam i2_3_lut_adj_1699.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1700 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[6] [7]), .O(n61415));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1700.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1701 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_748), .I3(GND_net), .O(n63255));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1701.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1702 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(n60927), .I3(Kp_23__N_869), .O(n25732));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1702.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1703 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n63380), .I3(\data_in_frame[7] [3]), .O(n55540));
    defparam i2_3_lut_4_lut_adj_1703.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_221_i3_3_lut_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\data_out_frame[25] [4]), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n61233), .O(n3_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_221_i3_3_lut_4_lut.LUT_INIT = 16'h6090;
    SB_LUT4 select_787_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1704 (.I0(n25687), .I1(n61261), .I2(\data_in_frame[1]_c [0]), 
            .I3(n61055), .O(n25987));
    defparam i1_2_lut_4_lut_adj_1704.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_4_lut_adj_1705 (.I0(\data_in_frame[0] [6]), .I1(n26_adj_5669), 
            .I2(n26126), .I3(n61055), .O(n30_adj_5670));
    defparam i13_4_lut_adj_1705.LUT_INIT = 16'h0804;
    SB_LUT4 n72071_bdd_4_lut (.I0(n72071), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8][3] ), .I3(byte_transmit_counter[1]), 
            .O(n65433));
    defparam n72071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1706 (.I0(\data_in_frame[16] [5]), .I1(n61185), 
            .I2(GND_net), .I3(GND_net), .O(n56748));
    defparam i1_2_lut_adj_1706.LUT_INIT = 16'h9999;
    SB_LUT4 i11_4_lut_adj_1707 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1][2] ), 
            .I2(n26447), .I3(\data_in_frame[1]_c [5]), .O(n28_adj_5671));
    defparam i11_4_lut_adj_1707.LUT_INIT = 16'h0800;
    SB_LUT4 select_787_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1708 (.I0(\data_in_frame[6] [7]), .I1(n25591), 
            .I2(n26123), .I3(GND_net), .O(n61254));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1708.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1709 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[4] [7]), .I3(\data_in_frame[7] [1]), .O(n60871));
    defparam i1_2_lut_4_lut_adj_1709.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_173_i2_4_lut (.I0(\data_out_frame[21] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_173_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1710 (.I0(n55617), .I1(\data_in_frame[21] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n55692));
    defparam i1_2_lut_adj_1710.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1711 (.I0(\data_in_frame[5] [0]), .I1(n25598), 
            .I2(\data_in_frame[2] [3]), .I3(n61092), .O(n26120));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1711.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_54795 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n71873));
    defparam byte_transmit_counter_0__bdd_4_lut_54795.LUT_INIT = 16'he4aa;
    SB_LUT4 i32775_3_lut (.I0(control_mode_c[5]), .I1(\data_in_frame[1]_c [5]), 
            .I2(n22465), .I3(GND_net), .O(n29735));
    defparam i32775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1712 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n25598));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1712.LUT_INIT = 16'h9696;
    SB_LUT4 n71873_bdd_4_lut (.I0(n71873), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n71876));
    defparam n71873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1713 (.I0(n56535), .I1(n56678), .I2(\data_in_frame[15] [5]), 
            .I3(\data_in_frame[17] [6]), .O(n61285));
    defparam i1_2_lut_4_lut_adj_1713.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1714 (.I0(\data_in_frame[21] [3]), .I1(n25923), 
            .I2(n61062), .I3(GND_net), .O(n60947));
    defparam i1_3_lut_adj_1714.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut_54897 (.I0(byte_transmit_counter[2]), 
            .I1(n65433), .I2(n65364), .I3(byte_transmit_counter[3]), .O(n71867));
    defparam byte_transmit_counter_2__bdd_4_lut_54897.LUT_INIT = 16'he4aa;
    SB_LUT4 i32774_3_lut (.I0(control_mode_c[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n22465), .I3(GND_net), .O(n29737));
    defparam i32774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71867_bdd_4_lut (.I0(n71867), .I1(n65333), .I2(n65332), .I3(byte_transmit_counter[3]), 
            .O(n71870));
    defparam n71867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1715 (.I0(\data_out_frame[25] [5]), .I1(n62684), 
            .I2(\data_out_frame[23] [3]), .I3(GND_net), .O(n60816));
    defparam i1_2_lut_3_lut_adj_1715.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[20] [2]), .I3(\data_in_frame[17] [0]), .O(n64725));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1717 (.I0(control_mode_c[5]), .I1(\control_mode[6] ), 
            .I2(\control_mode[7] ), .I3(GND_net), .O(n21));
    defparam i1_2_lut_3_lut_adj_1717.LUT_INIT = 16'hfefe;
    SB_LUT4 select_787_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n64725), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[16] [3]), .I3(\data_in_frame[14] [3]), .O(n64727));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5557));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_55016 (.I0(byte_transmit_counter[3]), 
            .I1(n70569), .I2(n68456), .I3(byte_transmit_counter[4]), .O(n72065));
    defparam byte_transmit_counter_3__bdd_4_lut_55016.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_165_i2_4_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_165_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i12_4_lut_adj_1719 (.I0(\data_in_frame[1][6] ), .I1(n24), .I2(Kp_23__N_748), 
            .I3(n60924), .O(n29_c));
    defparam i12_4_lut_adj_1719.LUT_INIT = 16'h0880;
    SB_LUT4 i48100_4_lut (.I0(n25591), .I1(n26154), .I2(n55137), .I3(n63255), 
            .O(n65181));
    defparam i48100_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n60822), .I1(n61134), .I2(n64729), 
            .I3(n64727), .O(n64735));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1721 (.I0(n65181), .I1(n29_c), .I2(n28_adj_5671), 
            .I3(n30_adj_5670), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1721.LUT_INIT = 16'h4000;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n56507), .I1(n61113), .I2(n56640), 
            .I3(n64735), .O(n64741));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n61073), .I1(n56684), .I2(n59626), 
            .I3(n64741), .O(n64747));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n61224), .I1(n55576), .I2(n60960), 
            .I3(n64747), .O(n64753));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n63317), .I1(n55617), .I2(n56555), 
            .I3(n64753), .O(n64759));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1726 (.I0(n1961), .I1(n1958), .I2(n1964), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n62533));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1726.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_1727 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(n64685), .I3(GND_net), .O(n6_adj_5434));
    defparam i1_2_lut_3_lut_adj_1727.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1728 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(n25281), .I3(\FRAME_MATCHER.i [1]), .O(n5));
    defparam i1_3_lut_4_lut_adj_1728.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_3_lut_4_lut_adj_1729 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n39534), .O(n25260));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1729.LUT_INIT = 16'ha8aa;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [2]), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'ha088;
    SB_LUT4 i1_3_lut_adj_1731 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[21] [7]), 
            .I2(n61298), .I3(GND_net), .O(n64679));
    defparam i1_3_lut_adj_1731.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n60906), .I1(n61388), .I2(n56559), 
            .I3(n64759), .O(n63040));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n61301), .I1(n63040), .I2(n60966), 
            .I3(n64679), .O(n61051));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14186_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n30047));
    defparam i14186_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14189_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n30050));
    defparam i14189_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14192_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n30053));
    defparam i14192_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14195_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n30056));
    defparam i14195_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14198_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n30059));
    defparam i14198_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14201_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n30062));
    defparam i14201_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14204_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n30065));
    defparam i14204_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13237_3_lut_4_lut (.I0(n39467), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29098));
    defparam i13237_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13880_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [6]), 
            .I3(neopxl_color[22]), .O(n29741));   // verilog/coms.v(130[12] 305[6])
    defparam i13880_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_787_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i51692_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n68363));   // verilog/coms.v(158[12:15])
    defparam i51692_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n72065_bdd_4_lut (.I0(n72065), .I1(n72026), .I2(n7_adj_5672), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n72065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i4_4_lut_adj_1734 (.I0(n60963), .I1(\data_in_frame[20] [7]), 
            .I2(n56748), .I3(n61310), .O(n10_adj_5673));
    defparam i4_4_lut_adj_1734.LUT_INIT = 16'h9669;
    SB_LUT4 i14021_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29882));
    defparam i14021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1735 (.I0(\data_in_frame[18] [5]), .I1(n10_adj_5673), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n56596));
    defparam i5_3_lut_adj_1735.LUT_INIT = 16'h9696;
    SB_LUT4 i14024_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29885));
    defparam i14024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14027_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29888));
    defparam i14027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1736 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[6] [6]), 
            .I2(n26126), .I3(\data_in_frame[7] [0]), .O(n60828));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1736.LUT_INIT = 16'h6996;
    SB_LUT4 i14030_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29891));
    defparam i14030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32772_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(\data_in_frame[0] [5]), 
            .I3(rx_data[5]), .O(n29894));
    defparam i32772_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i1_2_lut_adj_1737 (.I0(n60828), .I1(n61254), .I2(GND_net), 
            .I3(GND_net), .O(n26089));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1737.LUT_INIT = 16'h6666;
    SB_LUT4 i14036_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29897));
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13892_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [2]), 
            .I3(neopxl_color[10]), .O(n29753));   // verilog/coms.v(130[12] 305[6])
    defparam i13892_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1738 (.I0(\data_in_frame[8][6] ), .I1(n25556), 
            .I2(n26089), .I3(\data_in_frame[11] [2]), .O(n60938));
    defparam i3_4_lut_adj_1738.LUT_INIT = 16'h6996;
    SB_LUT4 i14039_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29900));
    defparam i14039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13819_3_lut_4_lut (.I0(n8), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29680));
    defparam i13819_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1739 (.I0(n17), .I1(n21), .I2(control_mode[0]), 
            .I3(control_mode[1]), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1739.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_1740 (.I0(\data_in_frame[10] [7]), .I1(n60987), 
            .I2(GND_net), .I3(GND_net), .O(n55679));
    defparam i1_2_lut_adj_1740.LUT_INIT = 16'h6666;
    SB_LUT4 i14162_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n30023));
    defparam i14162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14165_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n30026));
    defparam i14165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14168_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n30029));
    defparam i14168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13891_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[5] [3]), 
            .I3(neopxl_color[11]), .O(n29752));   // verilog/coms.v(130[12] 305[6])
    defparam i13891_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1741 (.I0(n26447), .I1(n61412), .I2(n23704), 
            .I3(GND_net), .O(n17_adj_5385));
    defparam i1_2_lut_3_lut_adj_1741.LUT_INIT = 16'h6060;
    SB_LUT4 i14171_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n30032));
    defparam i14171_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14174_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n30035));
    defparam i14174_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1742 (.I0(\data_in_frame[15] [4]), .I1(n60969), 
            .I2(n60940), .I3(\data_in_frame[13] [3]), .O(n56678));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'h6996;
    SB_LUT4 i14177_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n30038));
    defparam i14177_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14180_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n30041));
    defparam i14180_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14183_3_lut_4_lut (.I0(n8_adj_5551), .I1(n60760), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n30044));
    defparam i14183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1743 (.I0(n25687), .I1(n61261), .I2(\data_in_frame[0] [7]), 
            .I3(n60861), .O(n64873));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut_adj_1743.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65349), .I3(n65347), .O(n7_adj_5672));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65403), .I3(n65401), .O(n7_adj_5553));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65412), .I3(n65410), .O(n7_adj_5451));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65415), .I3(n65413), .O(n7));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_14));   // verilog/TinyFPGA_B.v(242[22:30])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1744 (.I0(\data_in_frame[13] [4]), .I1(n59626), 
            .I2(\data_in_frame[13] [3]), .I3(GND_net), .O(n56535));
    defparam i1_3_lut_adj_1744.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1745 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n61098));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1745.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1][6] ), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_772));   // verilog/coms.v(81[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65355), .I3(n65353), .O(n7_adj_5405));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n65406), .I3(n65404), .O(n7_adj_5442));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_3_lut_4_lut_adj_1746 (.I0(\data_in_frame[13] [4]), .I1(n60996), 
            .I2(\data_in_frame[13] [2]), .I3(n55550), .O(n60903));   // verilog/coms.v(88[17:63])
    defparam i1_3_lut_4_lut_adj_1746.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1747 (.I0(\data_in_frame[13] [4]), .I1(n60996), 
            .I2(n61129), .I3(n25746), .O(n55705));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_4_lut_adj_1747.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1748 (.I0(\data_in_frame[0] [0]), .I1(n61352), 
            .I2(Kp_23__N_772), .I3(\data_in_frame[1]_c [5]), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1748.LUT_INIT = 16'h6996;
    SB_LUT4 i13900_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[6] [2]), 
            .I3(neopxl_color[2]), .O(n29761));   // verilog/coms.v(130[12] 305[6])
    defparam i13900_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1749 (.I0(control_mode[0]), .I1(n17), 
            .I2(n21), .I3(control_mode[1]), .O(n15_adj_15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1749.LUT_INIT = 16'hfeff;
    SB_LUT4 i4_4_lut_adj_1750 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8][5] ), 
            .I2(\data_in_frame[6] [3]), .I3(n6_adj_5550), .O(n25647));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1750.LUT_INIT = 16'h6996;
    SB_LUT4 i12170_1_lut (.I0(n3483), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28031));   // verilog/coms.v(148[4] 304[11])
    defparam i12170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1751 (.I0(control_mode[0]), .I1(n17), 
            .I2(n21), .I3(control_mode[1]), .O(n15_adj_16));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1752 (.I0(\data_in_frame[3] [5]), .I1(n55544), 
            .I2(n61267), .I3(n60837), .O(n16));   // verilog/coms.v(81[16:27])
    defparam i6_4_lut_adj_1752.LUT_INIT = 16'h6996;
    SB_LUT4 i13885_3_lut_4_lut_4_lut (.I0(reset), .I1(n32326), .I2(\data_in_frame[4] [1]), 
            .I3(neopxl_color[17]), .O(n29746));   // verilog/coms.v(130[12] 305[6])
    defparam i13885_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1753 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(n60855));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_3_lut_adj_1753.LUT_INIT = 16'h9696;
    uart_tx tx (.r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3536[1] (\r_SM_Main_2__N_3536[1] ), 
            .n1(n1), .tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data[7:1], 
            \tx_data[0] }), .n5227(n5227), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .GND_net(GND_net), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n29(n29), .n23(n23), .n62322(n62322), .n27(n27), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n60413(n60413), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n63831(n63831), .r_Clock_Count({r_Clock_Count}), .n27514(n27514), 
            .n29671(n29671), .n61481(n61481), .n29123(n29123), .tx_active(tx_active), 
            .n72442(n72442), .VCC_net(VCC_net), .n63819(n63819), .n6(n6_adj_17), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.GND_net(GND_net), .baudrate({baudrate}), .r_Rx_Data(r_Rx_Data), 
            .n29(n29), .n23(n23), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .r_SM_Main({r_SM_Main_adj_31}), .n27(n27), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), .n5224(n5224), 
            .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .clk16MHz(clk16MHz), 
            .RX_N_2(RX_N_2), .n25296(n25296), .VCC_net(VCC_net), .r_Clock_Count({r_Clock_Count_adj_32}), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_29 ), 
            .n60415(n60415), .n63843(n63843), .n27507(n27507), .n27511(n27511), 
            .n29674(n29674), .n56754(n56754), .rx_data_ready(rx_data_ready), 
            .n29679(n29679), .rx_data({rx_data}), .n29646(n29646), .n29645(n29645), 
            .n29644(n29644), .n29642(n29642), .n29641(n29641), .n29640(n29640), 
            .n29639(n29639), .n61483(n61483), .n6(n6_adj_30), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n64131(n64131), .n64079(n64079), .n64167(n64167), .n64205(n64205), 
            .n64169(n64169), .n64151(n64151), .n64133(n64133), .n64097(n64097), 
            .n4(n4), .n63821(n63821)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_SM_Main, \r_SM_Main_2__N_3536[1] , n1, tx_o, clk16MHz, 
            tx_data, n5227, \o_Rx_DV_N_3488[12] , GND_net, \o_Rx_DV_N_3488[24] , 
            n29, n23, n62322, n27, \r_Bit_Index[0] , n60413, \r_SM_Main_2__N_3545[0] , 
            n63831, r_Clock_Count, n27514, n29671, n61481, n29123, 
            tx_active, n72442, VCC_net, n63819, n6, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_SM_Main;
    input \r_SM_Main_2__N_3536[1] ;
    output n1;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    input n5227;
    input \o_Rx_DV_N_3488[12] ;
    input GND_net;
    input \o_Rx_DV_N_3488[24] ;
    input n29;
    input n23;
    input n62322;
    input n27;
    output \r_Bit_Index[0] ;
    output n60413;
    input \r_SM_Main_2__N_3545[0] ;
    input n63831;
    output [8:0]r_Clock_Count;
    output n27514;
    input n29671;
    output n61481;
    input n29123;
    output tx_active;
    input n72442;
    input VCC_net;
    output n63819;
    output n6;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n28833, n3, n22515;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n21335, n68413, n68410, n3_adj_5296;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n21334, n61591, o_Tx_Serial_N_3598;
    wire [8:0]n41;
    wire [2:0]n460;
    
    wire n28597, n63799, n63805, n65359, n65360, n65366, n65365, 
        n54624, n54623, n54622, n54621, n54620, n54619, n54618, 
        n54617, n71909;
    
    SB_LUT4 i54627_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3536[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28833));
    defparam i54627_4_lut.LUT_INIT = 16'h1115;
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n21335), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i52232_3_lut (.I0(n5227), .I1(\o_Rx_DV_N_3488[12] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n68413));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i52232_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i52223_4_lut (.I0(n68413), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n68410));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i52223_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n68410), .I1(n62322), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5296));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'hc0ca;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5296), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n22515), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n60413));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i5819_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n63831), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n21334));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i5819_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i5820_3_lut (.I0(n21334), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21335));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i5820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44553_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n61591));
    defparam i44553_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3598), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_2056__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n28833));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27514), 
            .D(n460[1]), .R(n28597));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27514), 
            .D(n460[2]), .R(n28597));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29671));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2336_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2336_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i44451_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n61481));
    defparam i44451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5227), .I2(n60413), 
            .I3(GND_net), .O(n63799));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), .I3(n63799), 
            .O(n63805));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(n63805), .I1(n61591), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n28597));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'h0323;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29123));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2329_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2329_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n72442));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i48269_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n65359));
    defparam i48269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48270_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n65360));
    defparam i48270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48276_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n65366));
    defparam i48276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48275_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n65365));
    defparam i48275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2056_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n54624), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2056_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n54623), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_9 (.CI(n54623), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n54624));
    SB_LUT4 r_Clock_Count_2056_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n54622), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_8 (.CI(n54622), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n54623));
    SB_LUT4 r_Clock_Count_2056_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n54621), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_7 (.CI(n54621), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n54622));
    SB_LUT4 r_Clock_Count_2056_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n54620), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_6 (.CI(n54620), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n54621));
    SB_LUT4 r_Clock_Count_2056_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n54619), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_5 (.CI(n54619), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n54620));
    SB_LUT4 r_Clock_Count_2056_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n54618), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_4 (.CI(n54618), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n54619));
    SB_LUT4 r_Clock_Count_2056_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n54617), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_3 (.CI(n54617), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n54618));
    SB_LUT4 r_Clock_Count_2056_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n54617));
    SB_LUT4 i54732_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n27514));
    defparam i54732_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n65365), 
            .I2(n65366), .I3(r_Bit_Index[2]), .O(n71909));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n71909_bdd_4_lut (.I0(n71909), .I1(n65360), .I2(n65359), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3598));
    defparam n71909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut (.I0(n60413), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n63819));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n22515));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n62322), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (GND_net, baudrate, r_Rx_Data, n29, n23, \o_Rx_DV_N_3488[12] , 
            r_SM_Main, n27, \o_Rx_DV_N_3488[24] , \r_SM_Main_2__N_3446[1] , 
            n5224, \o_Rx_DV_N_3488[8] , clk16MHz, RX_N_2, n25296, 
            VCC_net, r_Clock_Count, \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , 
            \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[7] , \r_Bit_Index[0] , 
            n60415, n63843, n27507, n27511, n29674, n56754, rx_data_ready, 
            n29679, rx_data, n29646, n29645, n29644, n29642, n29641, 
            n29640, n29639, n61483, n6, \o_Rx_DV_N_3488[0] , n64131, 
            n64079, n64167, n64205, n64169, n64151, n64133, n64097, 
            n4, n63821) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [31:0]baudrate;
    output r_Rx_Data;
    output n29;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    output [2:0]r_SM_Main;
    output n27;
    output \o_Rx_DV_N_3488[24] ;
    input \r_SM_Main_2__N_3446[1] ;
    input n5224;
    output \o_Rx_DV_N_3488[8] ;
    input clk16MHz;
    input RX_N_2;
    output n25296;
    input VCC_net;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[7] ;
    output \r_Bit_Index[0] ;
    output n60415;
    input n63843;
    output n27507;
    output n27511;
    input n29674;
    input n56754;
    output rx_data_ready;
    input n29679;
    output [7:0]rx_data;
    input n29646;
    input n29645;
    input n29644;
    input n29642;
    input n29641;
    input n29640;
    input n29639;
    output n61483;
    output n6;
    output \o_Rx_DV_N_3488[0] ;
    input n64131;
    output n64079;
    input n64167;
    output n64205;
    output n64169;
    output n64151;
    output n64133;
    output n64097;
    output n4;
    output n63821;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2945;
    wire [23:0]n8261;
    wire [23:0]n294;
    
    wire n3053, n33, n2943, n3051, n37, n2949, n3057, n2950, 
        n3058, n23_c, n25, n2956, n3064, n2957, n3065, n60447, 
        n68310, n68307, n68304, n28831, n63775, n63781, n27630, 
        n11, n2947, n3055, n2948, n3056, n27_adj_5024, n29_adj_5025, 
        n2951, n3059, n2955, n3063, n13, n21, n2952, n3060, 
        n2953, n3061, n2954, n3062, n15, n17, n19, n538, n3054, 
        n31, n69120, n858, n698, n70105, n70609, n70601, n69122, 
        n2240;
    wire [23:0]n8105;
    
    wire n2366, n856, n2239, n2365, n3066, n8, n1011, n2238, 
        n2364, n1460, n70804, n2237, n2363, n70805, n16, n39, 
        n34, n35, n69112, n1459, n2236, n2362, n14, n69109, 
        n71303, n69822, n1602, n10, n70810, n70811, n69141, n70085, 
        n12, n20, n69820, n2235, n2361, n70984, n71506, n70886, 
        n71546, n3049, n71547, n68398, n68404, n68395, n3048, 
        n71062, n68401, n3, n3047, n71063, n1742, n2234, n2360, 
        n2829;
    wire [23:0]n8235;
    
    wire n2940, n2828, n2939, n2830, n2941, n41, n2832, n37_adj_5026, 
        n2833, n2944, n35_adj_5027, n2713;
    wire [23:0]n8209;
    
    wire n2827, n1879, n2714, n2233, n2359, n2719, n2831, n39_adj_5028, 
        n2718, n37_adj_5029, n2715, n43, n2716, n41_adj_5030, n2835, 
        n31_adj_5031;
    wire [23:0]n8131;
    
    wire n2353, n2638, n54066, n2354, n2519, n54065, n2834, n33_adj_5032, 
        n2838, n25_adj_5033, n2837, n27_adj_5034, n2836, n29_adj_5035, 
        n3_adj_5036, n2843, n15_adj_5037, n2842, n17_adj_5038, n2841, 
        n19_adj_5039, n2840, n21_adj_5040, n2839, n23_adj_5041, r_Rx_Data_R, 
        n35_adj_5042, n69297, n2844, n70254, n70677, n70673, n69304, 
        n2845, n12_adj_5043, n70826, n2355, n2397, n54064, n2013, 
        n2232, n2358, n20_adj_5044, n38, n70827, n69279, n18, 
        n69271, n71277, n2356, n2272, n54063, n69804, n16_adj_5045, 
        n24, n14_adj_5046, n69329, n71295, n71296, n71135, n71012, 
        n71498, n69802, n2357, n2144, n54062, n71548, n71549, 
        n2231, n2721, n2722, n2946, n29_adj_5047, n31_adj_5048, 
        n2723, n2724, n2725, n23_adj_5049, n25_adj_5050, n27_adj_5051, 
        n2717, n2942, n39_adj_5052, n2729, n2730, n54061, n13_adj_5053, 
        n15_adj_5054, n2720, n33_adj_5055, n2728, n2726, n2230, 
        n2604;
    wire [23:0]n8183;
    
    wire n2596, n2599, n54060, n41_adj_5056, n2597, n45, n2600, 
        n39_adj_5057, n54059, n2602, n54058, n2603, n54057, n33_adj_5058, 
        n54056, n35_adj_5059, n2598, n54055, n43_adj_5060, n2611, 
        n54054, n54053, n2612, n17_adj_5061, n2727, n19_adj_5062, 
        n2607, n2608, n2601, n2609, n21_adj_5063, n23_adj_5064, 
        n25_adj_5065, n2367, n54052, n37_adj_5066, n2229, n25388, 
        n63707, n61824, n2605, n2606, n27_adj_5067, n29_adj_5068, 
        n31_adj_5069, n69378, n70295, n70701, n64425, n3_adj_5070, 
        n64429, n5, n64433, n8_adj_5071;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n2227, n54045, n2228, n54044, n70697;
    wire [7:0]n1;
    
    wire n69383, n65165, n65275, n2, n10006, n54043, n14_adj_5073, 
        n54042, n54041, n70838, n70839, n54040, n54039, n54038, 
        n22, n40, n54037, n54036, n69369, n54035, n54034, n2099;
    wire [23:0]n8079;
    
    wire n20_adj_5074, n69363, n70882, n2100, n43_adj_5075, n2101, 
        n54033, n41_adj_5076, n69798, n2102, n39_adj_5077, n2103, 
        n37_adj_5078, n25411, n48, n2104, n54032, n2106, n2105, 
        n31_adj_5079, n33_adj_5080, n35_adj_5081, n2108, n18_adj_5082, 
        n26, n16_adj_5083, n69395, n71289, n71290, n63705, n61828, 
        n71143, n2109, n2107, n25_adj_5084, n27_adj_5085, n29_adj_5086, 
        n2110, n23_adj_5087, n68564, n68560, n71024, n22_adj_5088, 
        n28, n30, n71353, n26_adj_5089, n34_adj_5090, n24_adj_5091, 
        n68556, n71409, n69796, n71410, n71286, n71355, n70743, 
        n68562, n71082, n42, n71339, n2476;
    wire [23:0]n8157;
    
    wire n71340, n2487, n2477, n2481, n1967;
    wire [23:0]n8053;
    
    wire n1971, n37_adj_5092, n37_adj_5093, n1968, n60695, n2478, 
        n43_adj_5094, n68315, n68312, n2479, n1972, n41_adj_5095, 
        n35_adj_5096, n1977, n1969, n2480, n39_adj_5097, n2486, 
        n2485, n41_adj_5098, n1970, n39_adj_5099, n1973, n1975, 
        n1974, n29_adj_5100, n31_adj_5101, n27_adj_5102, n29_adj_5103, 
        n33_adj_5104, n1831;
    wire [23:0]n8027;
    
    wire n1966, n1833, n2489, n2610, n19_adj_5105, n21_adj_5106, 
        n1838, n1832, n1837, n35_adj_5107, n2483, n1836, n37_adj_5108, 
        n1834, n41_adj_5109, n2482, n1835, n39_adj_5110, n1840, 
        n2484, n31_adj_5111, n33_adj_5112, n35_adj_5113, n1693;
    wire [23:0]n8001;
    
    wire n2491, n1694, n1697, n39_adj_5114, n1698, n37_adj_5121, 
        n39_adj_5122, n25437, n48_adj_5123, n1841, n1695, n43_adj_5124, 
        n45_adj_5125, n43_adj_5126, n2098, n54021, n41_adj_5127, n54020, 
        n54019, n54018, n33_adj_5128, n35_adj_5129, n37_adj_5130, 
        n54017, n54016, n29_adj_5131, n1696, n54015;
    wire [2:0]n479;
    
    wire n28600, n31_adj_5132, n41_adj_5133, n1700, n54014, n1699, 
        n48_adj_5134, n1839, n31_adj_5135, n33_adj_5136, n35_adj_5137, 
        n1702, n29_adj_5138, n68648, n54013, n21_adj_5139, n54012, 
        n2488, n23_adj_5140, n41_adj_5141, n54011, n32, n40_adj_5142, 
        n37_adj_5143, n54010, n28_adj_5144, n71096, n71097, n68642, 
        n30_adj_5145, n68637, n71094, n70849, n71394, n71395, n1553;
    wire [23:0]n7975;
    
    wire n39_adj_5146, n1552, n1554, n43_adj_5147, n1556, n39_adj_5148, 
        n1557, n37_adj_5149, n1555, n41_adj_5150, n1558, n1414;
    wire [23:0]n7949;
    
    wire n1409, n1410, n43_adj_5151, n1408, n63701, n48_adj_5152, 
        n1560, n1411, n1413, n37_adj_5153, n41_adj_5154, n1261;
    wire [23:0]n7923;
    
    wire n1262, n45_adj_5155, n35_adj_5156, n1266, n1264, n41_adj_5157, 
        n1412, n39_adj_5158, n1263, n43_adj_5159, n1115;
    wire [23:0]n7897;
    
    wire n1265, n1112, n1111, n1113, n29_adj_5160, n31_adj_5161, 
        n1116, n1114, n41_adj_5162, n38_adj_5163, n40_adj_5164, n36, 
        n68729, n71403, n71404, n71294, n961, n40_adj_5165, n959, 
        n62259, n44_adj_5166, n46, n61512, n960, n9783, n21502, 
        n21504, n962, n42_adj_5167, n43_adj_5168, n25353, n48_adj_5169, 
        n803, n62307, n44_adj_5170, n46_adj_5171, n61510, n804, 
        n42_adj_5172, n64625, n64627, n64537, n64533, n64535, n64531, 
        n64517, n64447, n64529, n64437, n25376, n61508, n805, 
        n42_adj_5173, n71116, n71117, n48_adj_5174, n68723, n48_adj_5175, 
        n64383, n33_adj_5176, n64543, n64487, n64483, n25429, n64241, 
        n64261, n64489, n25426, n25423, n65018, n64465, n63715, 
        n64467, n64405, n64473, n39219, n64331, n62319, n62748, 
        n68324, n61539, n64475, n68325, n23_adj_5177, n25_adj_5178, 
        n64461, n65132, n64409, n64463, n65271, n27_adj_5179, n64623, 
        n65067, n21_adj_5180, n68544, n63625, n63623, n64271, n64267, 
        n64269, n64265, n65235, n68540, n64277, n63665, n65116, 
        n39221, n63983, n64001, n65219, n65120, n65069, n65291, 
        n20_adj_5181, n26_adj_5182, n28_adj_5183, n64039, n65213, 
        n64067, n65289, n68718, n71576, n24_adj_5184, n32_adj_5185, 
        n22_adj_5186, n68538, n71411, n71412, n71284, n64275, n70739, 
        n68542, n71413, n71151, n71514, n71515, n71419, n64273, 
        n72443, n25_adj_5187, n63811, n27_adj_5188, n63817, n2490, 
        n64287, n19_adj_5189, n68516, n68512, n70737, n18_adj_5190, 
        n70902, n70903, n68514, n70341, n24_adj_5191, n26_adj_5192, 
        n69780, n64289, n68374, n46_adj_5193, n48_adj_5194, n64417, 
        n64545, n25391, n22_adj_5195, n30_adj_5196, n20_adj_5197, 
        n68508, n71415, n71416, n64629, n64485, n61796, n71280, 
        n69494, n70878, n71157, n71351, n21488, n21490;
    wire [23:0]n8313;
    
    wire n3151, n3186, n54340, n3152, n3082, n54339, n3153, n3188, 
        n54338, n3154, n3084, n54337, n3155, n2977, n54336, n44_adj_5198, 
        n3156, n2867, n54335, n3157, n2754, n54334, n3158, n54333, 
        n23_adj_5199, n3159, n54332, n3160, n54331, n3161, n54330, 
        n3162, n54329, n3163, n54328, n3164, n54327, n54000, n3165, 
        n54326, n53999, n3166, n54325, n53998, n3167, n54324, 
        n3168, n54323, n53997, n3169, n54322, n53996, n3170, n54321, 
        n53995, n3171, n54320, n53994, n3172, n54319, n63721, 
        n54318, n53993, n25_adj_5200, n53992, n53991, n1976, n53990, 
        n53989, n53988, n53987, n53986, n61816, n53985, n61857, 
        n42_adj_5201, n71114, n53984, n53983, n71115, n53982, n65267;
    wire [23:0]n8287;
    
    wire n3046, n54299, n53981, n54298, n54297, n53980, n54296, 
        n53979, n3050, n54295, n54294, n53978, n3052, n54293, 
        n54292, n54291, n17_adj_5202, n63703, n61837, n54290, n54289, 
        n54288, n54287, n54286, n69457, n54285, n54284, n54283, 
        n54282, n54281, n54280, n54279, n63719, n61800, n38_adj_5203, 
        n40_adj_5204, n42_adj_5205, n68741, n71112, n71113, n61812, 
        n48_adj_5206, n69451, n61808, n63697, n1267, n1415, n34_adj_5207, 
        n71108, n65263, n61804, n71030, n16_adj_5208, n71109, n68709, 
        n69721, n36_adj_5209, n38_adj_5210, n44_adj_5211, n70449, 
        n70896, n39_adj_5212, n2938, n54261, n54260, n70897, n53943, 
        n53942, n53941, n53940, n53939, n53938, n69453, n70303, 
        n22_adj_5213, n70880, n53937, n53936, n1701, n53935, n69786, 
        n54259, n54258, n54257, n32_adj_5214, n71106, n71107, n68696, 
        n69713, n53908, n53907, n53906, n53905, n34_adj_5215, n70451, 
        n53904, n53903, n70841, n53902, n1559, n53901, n53900, 
        n71104, n53899, n41_adj_5216, n53898, n39_adj_5217, n53723, 
        n53897, n53722, n63607, n29_adj_5218, n65297, n53721, n63751, 
        n53896, n53720;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n71105, n53719, n63749, n53895, n53718, n63747, n31_adj_5219, 
        n53894, n53893, n33_adj_5220, n35_adj_5221, n53717, n53892, 
        n53716, n63745, n53715, n63743, n61846, n53714, n63605, 
        n37_adj_5222, n53891, n53890, n23_adj_5223, n53889, n25_adj_5224, 
        n7, n45_adj_5225, n53713, n63741, n53888, n53712, n53887, 
        n48_adj_5226, n53886, n9, n17_adj_5227, n53885, n21_adj_5228, 
        n53711, n53710, n63699, n61850, n11_adj_5229, n53709, n53708, 
        n53707, n13_adj_5230, n53706, n15_adj_5231, n27_adj_5232, 
        n53705, n53704, n53703, n53702, n19_adj_5233, n53701, n43_adj_5234, 
        n53700, n69005, n62613, n20_adj_5235, n28_adj_5236, n69015, 
        n16_adj_5237, n68979, n8_adj_5238, n53866, n53865, n24_adj_5239, 
        n53864, n53863, n53862, n3274, n69038, n53861, n61854, 
        n69989, n69979, n71190, n70533, n71366, n12_adj_5240, n48_adj_5241, 
        n4_c, n70790, n70791, n68999, n10_adj_5242, n30_adj_5243, 
        n69001, n18_adj_5244, n69446, n71275, n71311, n69848, n71510, 
        n71511, n6_adj_5245, n64515, n64505, n70792, n70793, n68981, 
        n70892, n54256, n69846, n54255, n54254, n71425, n54253, 
        n68989, n71356, n54252, n54251, n69854, n63677, n54250, 
        n71276, n54249, n3253, n54248, n54247, n71358, n54246, 
        n54245, n71163, n63685, n54244, n54243, n33_adj_5246, n54242, 
        n63717, n31_adj_5247, n37_adj_5248, n35_adj_5249, n25_adj_5250, 
        n61840, n27_adj_5251, n54232, n54231, n54230, n9_adj_5252, 
        n54229, n54228, n21_adj_5253, n32_adj_5254, n71102, n23_adj_5255, 
        n54227, n11_adj_5256, n54226, n19_adj_5257, n13_adj_5258, 
        n71103, n54225, n54224, n15_adj_5259, n68673, n69633, n54223, 
        n54222, n54221, n54220, n54219, n54218, n70307, n54217, 
        n54216, n17_adj_5260, n54215, n54214, n29_adj_5261, n34_adj_5262, 
        n70453, n69074, n70845, n71100, n70047, n70577, n70575, 
        n69078, n6_adj_5263, n70894, n54197, n54196, n54195, n70798, 
        n54194, n54193, n71101, n54192, n54191, n54190, n54189, 
        n54188, n54187, n54186, n14_adj_5264, n32_adj_5265, n54185, 
        n69784, n70799, n54184, n71440, n54183, n71441, n69060, 
        n54182, n12_adj_5266, n69056, n71305, n54181, n54585, n69834, 
        n54180, n54584, n63713, n8_adj_5267, n70800, n54583, n54582, 
        n70801, n54581, n54580, n54579, n69086, n70035, n10_adj_5268, 
        n70890, n69832, n70976, n71508, n71090, n71556, n71557, 
        n71553, n71341, n71342, n29_adj_5269, n31_adj_5270, n54156, 
        n54155, n54154, n54153, n54152, n54151, n54150, n54149, 
        n33_adj_5271, n54148, n54147, n54146, n54145, n27_adj_5272, 
        n54144, n54143, n54142, n54141, n68627, n54140, n63711, 
        n30_adj_5273, n38_adj_5274, n26_adj_5275, n65022, n71092, 
        n71093, n54112, n54111, n54110, n54109, n54108, n54107, 
        n54106, n54105, n54104, n68621, n54103, n54102, n54101, 
        n28_adj_5276, n68619, n71405, n54100, n54099, n54098, n54097, 
        n70853, n63709, n61820, n71542, n71543, n71503, n48_adj_5277, 
        n65185, n65259, n64539, n17_adj_5278, n19_adj_5279, n64547, 
        n27_adj_5280, n65287, n68587, n30_adj_5281, n38_adj_5282, 
        n61831, n26_adj_5283, n21_adj_5284, n71144, n71145, n68575, 
        n28_adj_5285, n68573, n71407, n70857, n71544, n71545, n71501, 
        n65187, n65231, n69193, n70175, n70635, n70629, n69197, 
        n10_adj_5286, n70818, n70819, n18_adj_5287, n36_adj_5288, 
        n69186, n16_adj_5289, n69182, n71299, n69810, n14_adj_5290, 
        n22_adj_5291, n12_adj_5292, n69207, n71297, n71298, n71133, 
        n70996, n71504, n69808, n71558, n71559, n71555, n25379, 
        n14_adj_5293, n15_adj_5294;
    
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8261[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8261[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8261[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8261[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8261[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8261[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52335_2_lut (.I0(n60447), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n68310));
    defparam i52335_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i52327_4_lut (.I0(n68310), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n68307));
    defparam i52327_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51602_4_lut (.I0(n68307), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n68304));
    defparam i51602_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i54617_4_lut (.I0(r_SM_Main[2]), .I1(n68304), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(r_SM_Main[1]), .O(n28831));
    defparam i54617_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut (.I0(n60447), .I1(r_SM_Main[1]), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n63775));
    defparam i1_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_988 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n63775), .O(n63781));
    defparam i1_4_lut_adj_988.LUT_INIT = 16'h0100;
    SB_LUT4 i54533_4_lut (.I0(r_SM_Main[2]), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n63781), .O(n27630));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i54533_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8261[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8261[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8261[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8261[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8261[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8261[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8261[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52030_4_lut (.I0(n31), .I1(n19), .I2(n17), .I3(n15), .O(n69120));
    defparam i52030_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53015_4_lut (.I0(n13), .I1(n11), .I2(n3065), .I3(baudrate[2]), 
            .O(n70105));
    defparam i53015_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53519_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n70105), 
            .O(n70609));
    defparam i53519_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53511_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n70609), 
            .O(n70601));
    defparam i53511_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52032_4_lut (.I0(n31), .I1(n29_adj_5025), .I2(n27_adj_5024), 
            .I3(n70601), .O(n69122));
    defparam i52032_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8105[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8105[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8105[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53714_3_lut (.I0(n8), .I1(baudrate[13]), .I2(n31), .I3(GND_net), 
            .O(n70804));   // verilog/uart_rx.v(119[33:55])
    defparam i53714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8105[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53715_3_lut (.I0(n70804), .I1(baudrate[14]), .I2(n33), .I3(GND_net), 
            .O(n70805));   // verilog/uart_rx.v(119[33:55])
    defparam i53715_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16), .I1(baudrate[17]), 
            .I2(n39), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52022_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69120), 
            .O(n69112));
    defparam i52022_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8105[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54213_4_lut (.I0(n34), .I1(n14), .I2(n39), .I3(n69109), 
            .O(n71303));   // verilog/uart_rx.v(119[33:55])
    defparam i54213_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52732_3_lut (.I0(n70805), .I1(baudrate[15]), .I2(n35), .I3(GND_net), 
            .O(n69822));   // verilog/uart_rx.v(119[33:55])
    defparam i52732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53720_3_lut (.I0(n10), .I1(baudrate[10]), .I2(n25), .I3(GND_net), 
            .O(n70810));   // verilog/uart_rx.v(119[33:55])
    defparam i53720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53721_3_lut (.I0(n70810), .I1(baudrate[11]), .I2(n27_adj_5024), 
            .I3(GND_net), .O(n70811));   // verilog/uart_rx.v(119[33:55])
    defparam i53721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52995_4_lut (.I0(n27_adj_5024), .I1(n25), .I2(n23_c), .I3(n69141), 
            .O(n70085));
    defparam i52995_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12), .I1(baudrate[9]), 
            .I2(n23_c), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52730_3_lut (.I0(n70811), .I1(baudrate[12]), .I2(n29_adj_5025), 
            .I3(GND_net), .O(n69820));   // verilog/uart_rx.v(119[33:55])
    defparam i52730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8105[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53894_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n69122), 
            .O(n70984));
    defparam i53894_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54416_4_lut (.I0(n69822), .I1(n71303), .I2(n39), .I3(n69112), 
            .O(n71506));   // verilog/uart_rx.v(119[33:55])
    defparam i54416_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53796_4_lut (.I0(n69820), .I1(n20), .I2(n29_adj_5025), .I3(n70085), 
            .O(n70886));   // verilog/uart_rx.v(119[33:55])
    defparam i53796_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54456_4_lut (.I0(n70886), .I1(n71506), .I2(n39), .I3(n70984), 
            .O(n71546));   // verilog/uart_rx.v(119[33:55])
    defparam i54456_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54457_3_lut (.I0(n71546), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n71547));   // verilog/uart_rx.v(119[33:55])
    defparam i54457_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52084_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5224), .I3(\o_Rx_DV_N_3488[8] ), .O(n68398));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52084_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i52217_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n60447), 
            .I3(r_SM_Main[0]), .O(n68404));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52217_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i52079_4_lut (.I0(n68398), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n68395));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52079_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53972_3_lut (.I0(n71547), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n71062));   // verilog/uart_rx.v(119[33:55])
    defparam i53972_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52089_4_lut (.I0(n68404), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n68401));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52089_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n68401), .I1(n68395), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i53973_3_lut (.I0(n71062), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n71063));   // verilog/uart_rx.v(119[33:55])
    defparam i53973_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8105[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8235[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8235[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8235[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8235[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8235[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8209[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8209[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8105[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8209[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8209[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8209[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8209[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n54066), 
            .O(n8131[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2751_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n54065), 
            .O(n8131[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3_adj_5036), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52207_4_lut (.I0(n35_adj_5042), .I1(n23_adj_5041), .I2(n21_adj_5040), 
            .I3(n19_adj_5039), .O(n69297));
    defparam i52207_4_lut.LUT_INIT = 16'haaab;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 i53164_4_lut (.I0(n17_adj_5038), .I1(n15_adj_5037), .I2(n2844), 
            .I3(baudrate[2]), .O(n70254));
    defparam i53164_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53587_4_lut (.I0(n23_adj_5041), .I1(n21_adj_5040), .I2(n19_adj_5039), 
            .I3(n70254), .O(n70677));
    defparam i53587_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53583_4_lut (.I0(n29_adj_5035), .I1(n27_adj_5034), .I2(n25_adj_5033), 
            .I3(n70677), .O(n70673));
    defparam i53583_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52214_4_lut (.I0(n35_adj_5042), .I1(n33_adj_5032), .I2(n31_adj_5031), 
            .I3(n70673), .O(n69304));
    defparam i52214_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2751_16 (.CI(n54065), .I0(n2354), .I1(n2519), .CO(n54066));
    SB_LUT4 i53736_3_lut (.I0(n12_adj_5043), .I1(baudrate[13]), .I2(n35_adj_5042), 
            .I3(GND_net), .O(n70826));   // verilog/uart_rx.v(119[33:55])
    defparam i53736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n54064), 
            .O(n8131[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8105[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5044), .I1(baudrate[17]), 
            .I2(n43), .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53737_3_lut (.I0(n70826), .I1(baudrate[14]), .I2(n37_adj_5029), 
            .I3(GND_net), .O(n70827));   // verilog/uart_rx.v(119[33:55])
    defparam i53737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52189_4_lut (.I0(n41_adj_5030), .I1(n39_adj_5028), .I2(n37_adj_5029), 
            .I3(n69297), .O(n69279));
    defparam i52189_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54187_4_lut (.I0(n38), .I1(n18), .I2(n43), .I3(n69271), 
            .O(n71277));   // verilog/uart_rx.v(119[33:55])
    defparam i54187_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2751_15 (.CI(n54064), .I0(n2355), .I1(n2397), .CO(n54065));
    SB_LUT4 add_2751_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n54063), 
            .O(n8131[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52714_3_lut (.I0(n70827), .I1(baudrate[15]), .I2(n39_adj_5028), 
            .I3(GND_net), .O(n69804));   // verilog/uart_rx.v(119[33:55])
    defparam i52714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5045), .I1(baudrate[9]), 
            .I2(n27_adj_5034), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54205_4_lut (.I0(n24), .I1(n14_adj_5046), .I2(n27_adj_5034), 
            .I3(n69329), .O(n71295));   // verilog/uart_rx.v(119[33:55])
    defparam i54205_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54206_3_lut (.I0(n71295), .I1(baudrate[10]), .I2(n29_adj_5035), 
            .I3(GND_net), .O(n71296));   // verilog/uart_rx.v(119[33:55])
    defparam i54206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54045_3_lut (.I0(n71296), .I1(baudrate[11]), .I2(n31_adj_5031), 
            .I3(GND_net), .O(n71135));   // verilog/uart_rx.v(119[33:55])
    defparam i54045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53922_4_lut (.I0(n41_adj_5030), .I1(n39_adj_5028), .I2(n37_adj_5029), 
            .I3(n69304), .O(n71012));
    defparam i53922_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54408_4_lut (.I0(n69804), .I1(n71277), .I2(n43), .I3(n69279), 
            .O(n71498));   // verilog/uart_rx.v(119[33:55])
    defparam i54408_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52712_3_lut (.I0(n71135), .I1(baudrate[12]), .I2(n33_adj_5032), 
            .I3(GND_net), .O(n69802));   // verilog/uart_rx.v(119[33:55])
    defparam i52712_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_14 (.CI(n54063), .I0(n2356), .I1(n2272), .CO(n54064));
    SB_LUT4 add_2751_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n54062), 
            .O(n8131[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54458_4_lut (.I0(n69802), .I1(n71498), .I2(n43), .I3(n71012), 
            .O(n71548));   // verilog/uart_rx.v(119[33:55])
    defparam i54458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54459_3_lut (.I0(n71548), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n71549));   // verilog/uart_rx.v(119[33:55])
    defparam i54459_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8105[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8209[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8209[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8235[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8235[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8209[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8209[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8235[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8209[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8235[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8235[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_13 (.CI(n54062), .I0(n2357), .I1(n2144), .CO(n54063));
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8209[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8235[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8209[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8209[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8235[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8235[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n54061), 
            .O(n8131[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8235[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_12 (.CI(n54061), .I0(n2358), .I1(n2013), .CO(n54062));
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8209[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8235[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8209[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8209[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8235[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8105[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8183[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8183[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8183[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n54060), 
            .O(n8131[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8183[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8183[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_11 (.CI(n54060), .I0(n2359), .I1(n1879), .CO(n54061));
    SB_LUT4 add_2751_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n54059), 
            .O(n8131[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8183[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_10 (.CI(n54059), .I0(n2360), .I1(n1742), .CO(n54060));
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2751_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n54058), 
            .O(n8131[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_9 (.CI(n54058), .I0(n2361), .I1(n1602), .CO(n54059));
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8183[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n54057), 
            .O(n8131[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_8 (.CI(n54057), .I0(n2362), .I1(n1459), .CO(n54058));
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n54056), 
            .O(n8131[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8183[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_7 (.CI(n54056), .I0(n2363), .I1(n1460), .CO(n54057));
    SB_LUT4 add_2751_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n54055), 
            .O(n8131[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_6 (.CI(n54055), .I0(n2364), .I1(n1011), .CO(n54056));
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8183[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n54054), 
            .O(n8131[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_5 (.CI(n54054), .I0(n2365), .I1(n856), .CO(n54055));
    SB_LUT4 add_2751_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n54053), 
            .O(n8131[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8183[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8183[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_4 (.CI(n54053), .I0(n2366), .I1(n698), .CO(n54054));
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8183[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8183[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8183[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n54052), 
            .O(n8131[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_3 (.CI(n54052), .I0(n2367), .I1(n858), .CO(n54053));
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8105[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54624_3_lut (.I0(n25388), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25296));   // verilog/uart_rx.v(119[33:55])
    defparam i54624_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_2751_2_lut (.I0(n61824), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2751_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54052));
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8183[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8183[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52288_4_lut (.I0(n37_adj_5066), .I1(n25_adj_5065), .I2(n23_adj_5064), 
            .I3(n21_adj_5063), .O(n69378));
    defparam i52288_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53205_4_lut (.I0(n19_adj_5062), .I1(n17_adj_5061), .I2(n2729), 
            .I3(baudrate[2]), .O(n70295));
    defparam i53205_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53611_4_lut (.I0(n25_adj_5065), .I1(n23_adj_5064), .I2(n21_adj_5063), 
            .I3(n70295), .O(n70701));
    defparam i53611_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_989 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n64425));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_989.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5070));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_990 (.I0(r_Clock_Count[3]), .I1(n3_adj_5070), .I2(\o_Rx_DV_N_3488[4] ), 
            .I3(n64425), .O(n64429));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_991 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n64429), .O(n64433));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_991.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5071));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_992 (.I0(r_Clock_Count[6]), .I1(n8_adj_5071), .I2(n64433), 
            .I3(\o_Rx_DV_N_3488[7] ), .O(n60447));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfdfe;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n60415));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_2750_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n54045), 
            .O(n8105[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2750_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n54044), 
            .O(n8105[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53607_4_lut (.I0(n31_adj_5069), .I1(n29_adj_5068), .I2(n27_adj_5067), 
            .I3(n70701), .O(n70697));
    defparam i53607_4_lut.LUT_INIT = 16'hfeff;
    SB_DFFESR r_Clock_Count_2053__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27630), .D(n1[0]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_CARRY add_2750_15 (.CI(n54044), .I0(n2228), .I1(n2397), .CO(n54045));
    SB_LUT4 i52293_4_lut (.I0(n37_adj_5066), .I1(n35_adj_5059), .I2(n33_adj_5058), 
            .I3(n70697), .O(n69383));
    defparam i52293_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48084_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n60447), .I2(GND_net), 
            .I3(GND_net), .O(n65165));
    defparam i48084_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48194_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n65165), .O(n65275));
    defparam i48194_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n63843), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n65275), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n10006));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 add_2750_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n54043), 
            .O(n8105[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_14 (.CI(n54043), .I0(n2229), .I1(n2272), .CO(n54044));
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n10006), .I1(n2), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3_adj_5036));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_2750_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n54042), 
            .O(n8105[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_13 (.CI(n54042), .I0(n2230), .I1(n2144), .CO(n54043));
    SB_LUT4 add_2750_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n54041), 
            .O(n8105[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53748_3_lut (.I0(n14_adj_5073), .I1(baudrate[13]), .I2(n37_adj_5066), 
            .I3(GND_net), .O(n70838));   // verilog/uart_rx.v(119[33:55])
    defparam i53748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2750_12 (.CI(n54041), .I0(n2231), .I1(n2013), .CO(n54042));
    SB_LUT4 i53749_3_lut (.I0(n70838), .I1(baudrate[14]), .I2(n39_adj_5057), 
            .I3(GND_net), .O(n70839));   // verilog/uart_rx.v(119[33:55])
    defparam i53749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n54040), 
            .O(n8105[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_11 (.CI(n54040), .I0(n2232), .I1(n1879), .CO(n54041));
    SB_LUT4 add_2750_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n54039), 
            .O(n8105[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_10 (.CI(n54039), .I0(n2233), .I1(n1742), .CO(n54040));
    SB_LUT4 add_2750_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n54038), 
            .O(n8105[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_9 (.CI(n54038), .I0(n2234), .I1(n1602), .CO(n54039));
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n54037), 
            .O(n8105[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_8 (.CI(n54037), .I0(n2235), .I1(n1459), .CO(n54038));
    SB_LUT4 add_2750_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n54036), 
            .O(n8105[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52279_4_lut (.I0(n43_adj_5060), .I1(n41_adj_5056), .I2(n39_adj_5057), 
            .I3(n69378), .O(n69369));
    defparam i52279_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8105[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2750_7 (.CI(n54036), .I0(n2236), .I1(n1460), .CO(n54037));
    SB_LUT4 add_2750_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n54035), 
            .O(n8105[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_6 (.CI(n54035), .I0(n2237), .I1(n1011), .CO(n54036));
    SB_LUT4 add_2750_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n54034), 
            .O(n8105[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_5 (.CI(n54034), .I0(n2238), .I1(n856), .CO(n54035));
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8079[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53792_4_lut (.I0(n40), .I1(n20_adj_5074), .I2(n45), .I3(n69363), 
            .O(n70882));   // verilog/uart_rx.v(119[33:55])
    defparam i53792_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8079[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8079[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n54033), 
            .O(n8105[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52708_3_lut (.I0(n70839), .I1(baudrate[15]), .I2(n41_adj_5056), 
            .I3(GND_net), .O(n69798));   // verilog/uart_rx.v(119[33:55])
    defparam i52708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8079[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2750_4 (.CI(n54033), .I0(n2239), .I1(n698), .CO(n54034));
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8079[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(n25411), .I1(n48), .I2(baudrate[0]), .I3(GND_net), 
            .O(n2240));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8079[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n54032), 
            .O(n8105[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8079[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8079[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2750_3 (.CI(n54032), .I0(n2240), .I1(n858), .CO(n54033));
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8079[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_5082), .I1(baudrate[9]), 
            .I2(n29_adj_5068), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54199_4_lut (.I0(n26), .I1(n16_adj_5083), .I2(n29_adj_5068), 
            .I3(n69395), .O(n71289));   // verilog/uart_rx.v(119[33:55])
    defparam i54199_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54200_3_lut (.I0(n71289), .I1(baudrate[10]), .I2(n31_adj_5069), 
            .I3(GND_net), .O(n71290));   // verilog/uart_rx.v(119[33:55])
    defparam i54200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_2_lut (.I0(n61828), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2750_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54032));
    SB_LUT4 i54053_3_lut (.I0(n71290), .I1(baudrate[11]), .I2(n33_adj_5058), 
            .I3(GND_net), .O(n71143));   // verilog/uart_rx.v(119[33:55])
    defparam i54053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8079[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8079[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8079[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51474_4_lut (.I0(n29_adj_5086), .I1(n27_adj_5085), .I2(n25_adj_5084), 
            .I3(n23_adj_5087), .O(n68564));
    defparam i51474_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51470_4_lut (.I0(n35_adj_5081), .I1(n33_adj_5080), .I2(n31_adj_5079), 
            .I3(n68564), .O(n68560));
    defparam i51470_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53934_4_lut (.I0(n43_adj_5060), .I1(n41_adj_5056), .I2(n39_adj_5057), 
            .I3(n69383), .O(n71024));
    defparam i53934_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28), .I1(baudrate[7]), 
            .I2(n33_adj_5080), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54263_4_lut (.I0(n69798), .I1(n70882), .I2(n45), .I3(n69369), 
            .O(n71353));   // verilog/uart_rx.v(119[33:55])
    defparam i54263_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5089), .I1(baudrate[9]), 
            .I2(n37_adj_5078), .I3(GND_net), .O(n34_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54319_4_lut (.I0(n34_adj_5090), .I1(n24_adj_5091), .I2(n37_adj_5078), 
            .I3(n68556), .O(n71409));   // verilog/uart_rx.v(119[33:55])
    defparam i54319_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52706_3_lut (.I0(n71143), .I1(baudrate[12]), .I2(n35_adj_5059), 
            .I3(GND_net), .O(n69796));   // verilog/uart_rx.v(119[33:55])
    defparam i52706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54320_3_lut (.I0(n71409), .I1(baudrate[10]), .I2(n39_adj_5077), 
            .I3(GND_net), .O(n71410));   // verilog/uart_rx.v(119[33:55])
    defparam i54320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54196_3_lut (.I0(n71410), .I1(baudrate[11]), .I2(n41_adj_5076), 
            .I3(GND_net), .O(n71286));   // verilog/uart_rx.v(119[33:55])
    defparam i54196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54265_4_lut (.I0(n69796), .I1(n71353), .I2(n45), .I3(n71024), 
            .O(n71355));   // verilog/uart_rx.v(119[33:55])
    defparam i54265_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53653_4_lut (.I0(n41_adj_5076), .I1(n39_adj_5077), .I2(n37_adj_5078), 
            .I3(n68560), .O(n70743));
    defparam i53653_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53992_4_lut (.I0(n30), .I1(n22_adj_5088), .I2(n33_adj_5080), 
            .I3(n68562), .O(n71082));   // verilog/uart_rx.v(119[33:55])
    defparam i53992_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54059_3_lut (.I0(n71286), .I1(baudrate[12]), .I2(n43_adj_5075), 
            .I3(GND_net), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam i54059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54249_4_lut (.I0(n42), .I1(n71082), .I2(n43_adj_5075), .I3(n70743), 
            .O(n71339));   // verilog/uart_rx.v(119[33:55])
    defparam i54249_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8157[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54250_3_lut (.I0(n71339), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n71340));   // verilog/uart_rx.v(119[33:55])
    defparam i54250_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8157[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8157[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8157[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8053[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8053[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8053[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n60695));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8157[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52311_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5224), .I3(n60695), .O(n68315));
    defparam i52311_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i52304_4_lut (.I0(n68315), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n68312));
    defparam i52304_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8157[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8053[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(r_SM_Main[1]), .I1(n68312), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27507));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8053[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8053[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8157[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8157[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8157[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8053[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8053[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8053[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8053[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8027[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8027[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8157[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8027[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8027[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8027[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8157[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8027[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8027[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8157[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8027[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8027[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8157[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8001[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8157[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8131[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8001[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8131[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8001[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Clock_Count_2053__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27630), .D(n1[7]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27630), .D(n1[6]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27630), .D(n1[5]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27630), .D(n1[4]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27630), .D(n1[3]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27630), .D(n1[2]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27630), .D(n1[1]), .R(n28831));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8001[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_993 (.I0(n25437), .I1(n48_adj_5123), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_993.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8131[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8001[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8131[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8131[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n54021), 
            .O(n8079[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2749_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n54020), 
            .O(n8079[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_13 (.CI(n54020), .I0(n2099), .I1(n2272), .CO(n54021));
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8131[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n54019), 
            .O(n8079[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_12 (.CI(n54019), .I0(n2100), .I1(n2144), .CO(n54020));
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8131[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n54018), 
            .O(n8079[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8131[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2749_11 (.CI(n54018), .I0(n2101), .I1(n2013), .CO(n54019));
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2749_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n54017), 
            .O(n8079[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8131[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2749_10 (.CI(n54017), .I0(n2102), .I1(n1879), .CO(n54018));
    SB_LUT4 add_2749_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n54016), 
            .O(n8079[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8131[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8001[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2749_9 (.CI(n54016), .I0(n2103), .I1(n1742), .CO(n54017));
    SB_LUT4 add_2749_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n54015), 
            .O(n8079[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27511), 
            .D(n479[1]), .R(n28600));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27511), 
            .D(n479[2]), .R(n28600));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2749_8 (.CI(n54015), .I0(n2104), .I1(n1602), .CO(n54016));
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8001[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n54014), 
            .O(n8079[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8001[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_994 (.I0(n63707), .I1(n48_adj_5134), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2749_7 (.CI(n54014), .I0(n2105), .I1(n1459), .CO(n54015));
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8001[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51558_4_lut (.I0(n35_adj_5137), .I1(n33_adj_5136), .I2(n31_adj_5135), 
            .I3(n29_adj_5138), .O(n68648));
    defparam i51558_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8131[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n54013), 
            .O(n8079[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_6 (.CI(n54013), .I0(n2106), .I1(n1460), .CO(n54014));
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2749_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n54012), 
            .O(n8079[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_5 (.CI(n54012), .I0(n2107), .I1(n1011), .CO(n54013));
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2749_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n54011), 
            .O(n8079[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_4 (.CI(n54011), .I0(n2108), .I1(n856), .CO(n54012));
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32), .I1(baudrate[9]), 
            .I2(n43_adj_5124), .I3(GND_net), .O(n40_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2749_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n54010), 
            .O(n8079[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_3 (.CI(n54010), .I0(n2109), .I1(n698), .CO(n54011));
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54006_3_lut (.I0(n28_adj_5144), .I1(baudrate[5]), .I2(n35_adj_5137), 
            .I3(GND_net), .O(n71096));   // verilog/uart_rx.v(119[33:55])
    defparam i54006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54007_3_lut (.I0(n71096), .I1(baudrate[6]), .I2(n37_adj_5121), 
            .I3(GND_net), .O(n71097));   // verilog/uart_rx.v(119[33:55])
    defparam i54007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51552_4_lut (.I0(n41_adj_5133), .I1(n39_adj_5114), .I2(n37_adj_5121), 
            .I3(n68648), .O(n68642));
    defparam i51552_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54004_4_lut (.I0(n40_adj_5142), .I1(n30_adj_5145), .I2(n43_adj_5124), 
            .I3(n68637), .O(n71094));   // verilog/uart_rx.v(119[33:55])
    defparam i54004_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2749_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8079[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n54010));
    SB_LUT4 i53759_3_lut (.I0(n71097), .I1(baudrate[7]), .I2(n39_adj_5114), 
            .I3(GND_net), .O(n70849));   // verilog/uart_rx.v(119[33:55])
    defparam i53759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54304_4_lut (.I0(n70849), .I1(n71094), .I2(n43_adj_5124), 
            .I3(n68642), .O(n71394));   // verilog/uart_rx.v(119[33:55])
    defparam i54304_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54305_3_lut (.I0(n71394), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n71395));   // verilog/uart_rx.v(119[33:55])
    defparam i54305_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7975[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7975[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7975[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7975[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5148));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7975[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7975[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7975[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7949[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7949[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7949[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7949[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_995 (.I0(n63701), .I1(n48_adj_5152), .I2(GND_net), 
            .I3(GND_net), .O(n1560));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7949[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7949[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7923[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7923[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7923[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7923[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7923[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7897[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7897[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7897[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7897[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7897[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7897[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5163), .I1(baudrate[4]), 
            .I2(n41_adj_5162), .I3(GND_net), .O(n40_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54313_4_lut (.I0(n40_adj_5164), .I1(n36), .I2(n41_adj_5162), 
            .I3(n68729), .O(n71403));   // verilog/uart_rx.v(119[33:55])
    defparam i54313_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54314_3_lut (.I0(n71403), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n71404));   // verilog/uart_rx.v(119[33:55])
    defparam i54314_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54204_3_lut (.I0(n71404), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n71294));   // verilog/uart_rx.v(119[33:55])
    defparam i54204_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5165), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i4216_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n62259), .I3(n44_adj_5166), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i4216_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i742_4_lut (.I0(n61512), .I1(n294[18]), .I2(n46), .I3(baudrate[5]), 
            .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 i5983_4_lut (.I0(n960), .I1(n9783), .I2(n21502), .I3(baudrate[3]), 
            .O(n21504));   // verilog/uart_rx.v(119[33:55])
    defparam i5983_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5166), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i4194_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam i4194_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5982_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21502));   // verilog/uart_rx.v(119[33:55])
    defparam i5982_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5167), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_996 (.I0(n25353), .I1(n48_adj_5169), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_996.LUT_INIT = 16'hefef;
    SB_LUT4 i4045_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n62307), .I3(n44_adj_5170), 
            .O(n46_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam i4045_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i639_4_lut (.I0(n61510), .I1(n294[19]), .I2(n46_adj_5171), 
            .I3(baudrate[4]), .O(n61512));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5172), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_2_lut_adj_997 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n64625));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n64627));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_999 (.I0(n64537), .I1(n64533), .I2(n64535), .I3(n64531), 
            .O(n64517));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(n64625), .I1(n64447), .I2(n64529), 
            .I3(n64437), .O(n25376));
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i534_3_lut (.I0(n61508), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n61510));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54026_3_lut (.I0(n42_adj_5173), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n71116));   // verilog/uart_rx.v(119[33:55])
    defparam i54026_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54027_3_lut (.I0(n71116), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n71117));   // verilog/uart_rx.v(119[33:55])
    defparam i54027_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53735_3_lut (.I0(n71117), .I1(baudrate[4]), .I2(n61510), 
            .I3(GND_net), .O(n48_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam i53735_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i51633_2_lut (.I0(baudrate[1]), .I1(n294[20]), .I2(GND_net), 
            .I3(GND_net), .O(n68723));   // verilog/uart_rx.v(119[33:55])
    defparam i51633_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52292_4_lut (.I0(n25388), .I1(n68723), .I2(n48_adj_5175), 
            .I3(baudrate[0]), .O(n804));
    defparam i52292_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n64383));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1002 (.I0(n64383), .I1(n64543), .I2(n64487), 
            .I3(n64483), .O(n25429));
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n64437));
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(n64529), .I1(n64437), .I2(n64241), 
            .I3(baudrate[19]), .O(n64261));
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1005 (.I0(n64261), .I1(n64489), .I2(n64531), 
            .I3(n64487), .O(n25426));
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'hfffe;
    SB_LUT4 i47944_2_lut (.I0(baudrate[17]), .I1(n25423), .I2(GND_net), 
            .I3(GND_net), .O(n65018));
    defparam i47944_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n64465));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut (.I0(n71549), .I1(baudrate[19]), .I2(n2827), 
            .I3(n63715), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n64467));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n64405));
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'heeee;
    SB_LUT4 i54620_2_lut_4_lut (.I0(n71549), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25429), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i54620_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(n64473), .I1(n64537), .I2(baudrate[16]), 
            .I3(n39219), .O(n64331));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'h0100;
    SB_LUT4 i52403_3_lut (.I0(n62319), .I1(n62748), .I2(baudrate[2]), 
            .I3(GND_net), .O(n68324));   // verilog/uart_rx.v(119[33:55])
    defparam i52403_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i52211_4_lut (.I0(n61539), .I1(n64331), .I2(n64475), .I3(n64405), 
            .O(n68325));   // verilog/uart_rx.v(119[33:55])
    defparam i52211_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n68325), .I1(n68324), .I2(n294[21]), 
            .I3(n65018), .O(n61508));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n64461));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'heeee;
    SB_LUT4 i48053_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n65132));
    defparam i48053_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48190_4_lut (.I0(n65132), .I1(n64409), .I2(n64463), .I3(baudrate[9]), 
            .O(n65271));
    defparam i48190_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54745_2_lut (.I0(n48_adj_5175), .I1(n25388), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i54745_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n64623));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'heeee;
    SB_LUT4 i44501_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n61539));
    defparam i44501_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47990_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n65067));
    defparam i47990_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5180));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51454_4_lut (.I0(n27_adj_5179), .I1(n25_adj_5178), .I2(n23_adj_5177), 
            .I3(n21_adj_5180), .O(n68544));
    defparam i51454_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(n64543), .I1(n63625), .I2(n63623), 
            .I3(n64533), .O(n25423));
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i48154_4_lut (.I0(n64271), .I1(n64267), .I2(n64269), .I3(n64265), 
            .O(n65235));
    defparam i48154_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51450_4_lut (.I0(n33_adj_5176), .I1(n31_adj_5161), .I2(n29_adj_5160), 
            .I3(n68544), .O(n68540));
    defparam i51450_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(baudrate[17]), .I1(n64277), .I2(baudrate[2]), 
            .I3(n39219), .O(n63665));
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n65235), .I1(n63665), .I2(n25423), 
            .I3(n65116), .O(n62748));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n39221), .O(n63983));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(n63983), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n64001));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h0002;
    SB_LUT4 i48210_4_lut (.I0(n65219), .I1(n65116), .I2(n65120), .I3(n65069), 
            .O(n65291));
    defparam i48210_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(n65271), .I1(n65291), .I2(n61539), 
            .I3(n64001), .O(n62319));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n62319), .I1(baudrate[2]), 
            .I2(n62748), .I3(GND_net), .O(n48_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_5181));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5182), .I1(baudrate[7]), 
            .I2(n31_adj_5161), .I3(GND_net), .O(n28_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n64039));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h0100;
    SB_LUT4 i48132_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n65213));
    defparam i48132_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1019 (.I0(n61539), .I1(n64039), .I2(n64623), 
            .I3(baudrate[16]), .O(n64067));
    defparam i1_4_lut_adj_1019.LUT_INIT = 16'h0004;
    SB_LUT4 i48208_4_lut (.I0(n65213), .I1(n65116), .I2(n65120), .I3(n65069), 
            .O(n65289));
    defparam i48208_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54486_4_lut (.I0(n65271), .I1(n68718), .I2(n65289), .I3(n64067), 
            .O(n71576));
    defparam i54486_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5184), .I1(baudrate[9]), 
            .I2(n35_adj_5156), .I3(GND_net), .O(n32_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29674));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .D(n56754));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i54321_4_lut (.I0(n32_adj_5185), .I1(n22_adj_5186), .I2(n35_adj_5156), 
            .I3(n68538), .O(n71411));   // verilog/uart_rx.v(119[33:55])
    defparam i54321_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54322_3_lut (.I0(n71411), .I1(baudrate[10]), .I2(n37_adj_5143), 
            .I3(GND_net), .O(n71412));   // verilog/uart_rx.v(119[33:55])
    defparam i54322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54194_3_lut (.I0(n71412), .I1(baudrate[11]), .I2(n39_adj_5146), 
            .I3(GND_net), .O(n71284));   // verilog/uart_rx.v(119[33:55])
    defparam i54194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n64271));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n64275));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'heeee;
    SB_LUT4 i53649_4_lut (.I0(n39_adj_5146), .I1(n37_adj_5143), .I2(n35_adj_5156), 
            .I3(n68540), .O(n70739));
    defparam i53649_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54323_4_lut (.I0(n28_adj_5183), .I1(n20_adj_5181), .I2(n31_adj_5161), 
            .I3(n68542), .O(n71413));   // verilog/uart_rx.v(119[33:55])
    defparam i54323_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54061_3_lut (.I0(n71284), .I1(baudrate[12]), .I2(n41_adj_5141), 
            .I3(GND_net), .O(n71151));   // verilog/uart_rx.v(119[33:55])
    defparam i54061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54424_4_lut (.I0(n71151), .I1(n71413), .I2(n41_adj_5141), 
            .I3(n70739), .O(n71514));   // verilog/uart_rx.v(119[33:55])
    defparam i54424_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54425_3_lut (.I0(n71514), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n71515));   // verilog/uart_rx.v(119[33:55])
    defparam i54425_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54329_3_lut (.I0(n71515), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n71419));   // verilog/uart_rx.v(119[33:55])
    defparam i54329_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54065_3_lut (.I0(n71419), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam i54065_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n64273));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n64277));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n65069));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n29679));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29646));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29645));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29644));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29642));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29641));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29640));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29639));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n72443));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8131[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n64267));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8131[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2314_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2314_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i44453_2_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n61483));
    defparam i44453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i44551_2_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i44551_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5224), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60415), .O(n63811));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1027 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n63811), .O(n63817));
    defparam i1_4_lut_adj_1027.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(n63817), .I1(n6), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n28600));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'h0323;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n64265));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8131[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n64269));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(n64269), .I1(n64265), .I2(n64267), 
            .I3(n65069), .O(n64287));
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5189));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51426_4_lut (.I0(n25_adj_5187), .I1(n23_adj_5140), .I2(n21_adj_5139), 
            .I3(n19_adj_5189), .O(n68516));
    defparam i51426_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51422_4_lut (.I0(n31_adj_5132), .I1(n29_adj_5131), .I2(n27_adj_5188), 
            .I3(n68516), .O(n68512));
    defparam i51422_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53647_4_lut (.I0(n37_adj_5130), .I1(n35_adj_5129), .I2(n33_adj_5128), 
            .I3(n68512), .O(n70737));
    defparam i53647_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53812_3_lut (.I0(n18_adj_5190), .I1(baudrate[13]), .I2(n41_adj_5127), 
            .I3(GND_net), .O(n70902));   // verilog/uart_rx.v(119[33:55])
    defparam i53812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53813_3_lut (.I0(n70902), .I1(baudrate[14]), .I2(n43_adj_5126), 
            .I3(GND_net), .O(n70903));   // verilog/uart_rx.v(119[33:55])
    defparam i53813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2307_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2307_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53251_4_lut (.I0(n43_adj_5126), .I1(n41_adj_5127), .I2(n29_adj_5131), 
            .I3(n68514), .O(n70341));
    defparam i53251_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_5191), .I1(baudrate[7]), 
            .I2(n29_adj_5131), .I3(GND_net), .O(n26_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52690_3_lut (.I0(n70903), .I1(baudrate[15]), .I2(n45_adj_5125), 
            .I3(GND_net), .O(n69780));   // verilog/uart_rx.v(119[33:55])
    defparam i52690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(n64277), .I1(n64273), .I2(n64275), 
            .I3(n64271), .O(n64289));
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(n64289), .I1(n25426), .I2(n64287), 
            .I3(GND_net), .O(n25388));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n68374), .I1(baudrate[2]), 
            .I2(n71576), .I3(n48_adj_5175), .O(n46_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5193), .I1(baudrate[3]), 
            .I2(n61508), .I3(GND_net), .O(n48_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n64405), .I1(n64465), .I2(n64467), 
            .I3(n64463), .O(n64417));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n64417), .I1(n25429), .I2(n64409), 
            .I3(n64545), .O(n25391));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 i23457_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n39221));
    defparam i23457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1036 (.I0(n25391), .I1(n48_adj_5194), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1036.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5195), .I1(baudrate[9]), 
            .I2(n33_adj_5128), .I3(GND_net), .O(n30_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54325_4_lut (.I0(n30_adj_5196), .I1(n20_adj_5197), .I2(n33_adj_5128), 
            .I3(n68508), .O(n71415));   // verilog/uart_rx.v(119[33:55])
    defparam i54325_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i23455_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n39219));
    defparam i23455_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i54326_3_lut (.I0(n71415), .I1(baudrate[10]), .I2(n35_adj_5129), 
            .I3(GND_net), .O(n71416));   // verilog/uart_rx.v(119[33:55])
    defparam i54326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44756_1_lut_4_lut (.I0(n64627), .I1(n64629), .I2(n64485), 
            .I3(n64625), .O(n61796));
    defparam i44756_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54190_3_lut (.I0(n71416), .I1(baudrate[11]), .I2(n37_adj_5130), 
            .I3(GND_net), .O(n71280));   // verilog/uart_rx.v(119[33:55])
    defparam i54190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52404_4_lut (.I0(n43_adj_5126), .I1(n41_adj_5127), .I2(n39_adj_5122), 
            .I3(n70737), .O(n69494));
    defparam i52404_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53788_4_lut (.I0(n69780), .I1(n26_adj_5192), .I2(n45_adj_5125), 
            .I3(n70341), .O(n70878));   // verilog/uart_rx.v(119[33:55])
    defparam i53788_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54067_3_lut (.I0(n71280), .I1(baudrate[12]), .I2(n39_adj_5122), 
            .I3(GND_net), .O(n71157));   // verilog/uart_rx.v(119[33:55])
    defparam i54067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54261_4_lut (.I0(n71157), .I1(n70878), .I2(n45_adj_5125), 
            .I3(n69494), .O(n71351));   // verilog/uart_rx.v(119[33:55])
    defparam i54261_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8131[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5972_4_lut (.I0(n804), .I1(n39219), .I2(n21488), .I3(baudrate[2]), 
            .O(n21490));   // verilog/uart_rx.v(119[33:55])
    defparam i5972_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8157[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n54340), 
            .O(n8313[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n54339), 
            .O(n8313[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_24 (.CI(n54339), .I0(n3152), .I1(n3082), .CO(n54340));
    SB_LUT4 add_2758_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n54338), 
            .O(n8313[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_23 (.CI(n54338), .I0(n3153), .I1(n3188), .CO(n54339));
    SB_LUT4 add_2758_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n54337), 
            .O(n8313[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_22 (.CI(n54337), .I0(n3154), .I1(n3084), .CO(n54338));
    SB_LUT4 add_2758_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n54336), 
            .O(n8313[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_21 (.CI(n54336), .I0(n3155), .I1(n2977), .CO(n54337));
    SB_LUT4 div_37_i535_4_lut (.I0(n71576), .I1(n44_adj_5198), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 add_2758_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n54335), 
            .O(n8313[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_20 (.CI(n54335), .I0(n3156), .I1(n2867), .CO(n54336));
    SB_LUT4 add_2758_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n54334), 
            .O(n8313[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_19 (.CI(n54334), .I0(n3157), .I1(n2754), .CO(n54335));
    SB_LUT4 add_2758_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n54333), 
            .O(n8313[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_18 (.CI(n54333), .I0(n3158), .I1(n2638), .CO(n54334));
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2758_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n54332), 
            .O(n8313[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_17 (.CI(n54332), .I0(n3159), .I1(n2519), .CO(n54333));
    SB_LUT4 add_2758_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n54331), 
            .O(n8313[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_16 (.CI(n54331), .I0(n3160), .I1(n2397), .CO(n54332));
    SB_LUT4 add_2758_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n54330), 
            .O(n8313[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_15 (.CI(n54330), .I0(n3161), .I1(n2272), .CO(n54331));
    SB_LUT4 add_2758_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n54329), 
            .O(n8313[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_14 (.CI(n54329), .I0(n3162), .I1(n2144), .CO(n54330));
    SB_LUT4 add_2758_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n54328), 
            .O(n8313[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_13 (.CI(n54328), .I0(n3163), .I1(n2013), .CO(n54329));
    SB_LUT4 add_2758_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n54327), 
            .O(n8313[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_12 (.CI(n54327), .I0(n3164), .I1(n1879), .CO(n54328));
    SB_LUT4 add_2748_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n54000), 
            .O(n8053[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n54326), 
            .O(n8313[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_11 (.CI(n54326), .I0(n3165), .I1(n1742), .CO(n54327));
    SB_LUT4 add_2748_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n53999), 
            .O(n8053[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n54325), 
            .O(n8313[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_10 (.CI(n54325), .I0(n3166), .I1(n1602), .CO(n54326));
    SB_CARRY add_2748_13 (.CI(n53999), .I0(n1967), .I1(n2144), .CO(n54000));
    SB_LUT4 add_2748_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n53998), 
            .O(n8053[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n54324), 
            .O(n8313[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_9 (.CI(n54324), .I0(n3167), .I1(n1459), .CO(n54325));
    SB_CARRY add_2748_12 (.CI(n53998), .I0(n1968), .I1(n2013), .CO(n53999));
    SB_LUT4 add_2758_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n54323), 
            .O(n8313[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_8 (.CI(n54323), .I0(n3168), .I1(n1460), .CO(n54324));
    SB_LUT4 add_2748_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n53997), 
            .O(n8053[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_11 (.CI(n53997), .I0(n1969), .I1(n1879), .CO(n53998));
    SB_LUT4 add_2758_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n54322), 
            .O(n8313[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_7 (.CI(n54322), .I0(n3169), .I1(n1011), .CO(n54323));
    SB_LUT4 add_2748_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n53996), 
            .O(n8053[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_10 (.CI(n53996), .I0(n1970), .I1(n1742), .CO(n53997));
    SB_LUT4 add_2758_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n54321), 
            .O(n8313[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_6 (.CI(n54321), .I0(n3170), .I1(n856), .CO(n54322));
    SB_LUT4 add_2748_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n53995), 
            .O(n8053[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_9 (.CI(n53995), .I0(n1971), .I1(n1602), .CO(n53996));
    SB_LUT4 add_2758_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n54320), 
            .O(n8313[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_5 (.CI(n54320), .I0(n3171), .I1(n698), .CO(n54321));
    SB_LUT4 add_2748_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n53994), 
            .O(n8053[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_8 (.CI(n53994), .I0(n1972), .I1(n1459), .CO(n53995));
    SB_LUT4 add_2758_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n54319), 
            .O(n8313[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_4 (.CI(n54319), .I0(n3172), .I1(n858), .CO(n54320));
    SB_LUT4 add_2758_3_lut (.I0(n61796), .I1(GND_net), .I2(n538), .I3(n54318), 
            .O(n63721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2748_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n53993), 
            .O(n8053[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_7 (.CI(n53993), .I0(n1973), .I1(n1460), .CO(n53994));
    SB_CARRY add_2758_3 (.CI(n54318), .I0(GND_net), .I1(n538), .CO(n54319));
    SB_CARRY add_2758_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n54318));
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2748_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n53992), 
            .O(n8053[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_6 (.CI(n53992), .I0(n1974), .I1(n1011), .CO(n53993));
    SB_LUT4 add_2748_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n53991), 
            .O(n8053[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_5 (.CI(n53991), .I0(n1975), .I1(n856), .CO(n53992));
    SB_LUT4 add_2748_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n53990), 
            .O(n8053[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_4 (.CI(n53990), .I0(n1976), .I1(n698), .CO(n53991));
    SB_LUT4 add_2748_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n53989), 
            .O(n8053[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_3 (.CI(n53989), .I0(n1977), .I1(n858), .CO(n53990));
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_5170), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 add_2748_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53989));
    SB_LUT4 add_2747_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n53988), 
            .O(n8027[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n53987), 
            .O(n8027[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_12 (.CI(n53987), .I0(n1832), .I1(n2013), .CO(n53988));
    SB_LUT4 add_2747_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n53986), 
            .O(n8027[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_11 (.CI(n53986), .I0(n1833), .I1(n1879), .CO(n53987));
    SB_LUT4 i44776_1_lut (.I0(n25423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61816));
    defparam i44776_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 add_2747_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n53985), 
            .O(n8027[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(n64475), .I1(n25376), .I2(n64517), 
            .I3(n64473), .O(n25353));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'hfffe;
    SB_CARRY add_2747_10 (.CI(n53985), .I0(n1834), .I1(n1742), .CO(n53986));
    SB_LUT4 i23463_rep_5_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n61857));   // verilog/uart_rx.v(119[33:55])
    defparam i23463_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n61857), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i54024_3_lut (.I0(n42_adj_5201), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n71114));   // verilog/uart_rx.v(119[33:55])
    defparam i54024_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2747_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n53984), 
            .O(n8027[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_9 (.CI(n53984), .I0(n1835), .I1(n1602), .CO(n53985));
    SB_LUT4 add_2747_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n53983), 
            .O(n8027[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_8 (.CI(n53983), .I0(n1836), .I1(n1459), .CO(n53984));
    SB_LUT4 i54025_3_lut (.I0(n71114), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n71115));   // verilog/uart_rx.v(119[33:55])
    defparam i54025_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53739_3_lut (.I0(n71115), .I1(baudrate[5]), .I2(n61512), 
            .I3(GND_net), .O(n48_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam i53739_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 add_2747_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n53982), 
            .O(n8027[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_7 (.CI(n53982), .I0(n1837), .I1(n1460), .CO(n53983));
    SB_LUT4 i1_3_lut_adj_1038 (.I0(n65267), .I1(n48_adj_5174), .I2(baudrate[0]), 
            .I3(GND_net), .O(n962));
    defparam i1_3_lut_adj_1038.LUT_INIT = 16'h1010;
    SB_LUT4 add_2757_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n54299), 
            .O(n8287[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2747_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n53981), 
            .O(n8027[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n54298), 
            .O(n8287[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_22 (.CI(n54298), .I0(n3047), .I1(n3188), .CO(n54299));
    SB_CARRY add_2747_6 (.CI(n53981), .I0(n1838), .I1(n1011), .CO(n53982));
    SB_LUT4 add_2757_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n54297), 
            .O(n8287[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_21 (.CI(n54297), .I0(n3048), .I1(n3084), .CO(n54298));
    SB_LUT4 add_2747_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n53980), 
            .O(n8027[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n54296), 
            .O(n8287[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_20 (.CI(n54296), .I0(n3049), .I1(n2977), .CO(n54297));
    SB_CARRY add_2747_5 (.CI(n53980), .I0(n1839), .I1(n856), .CO(n53981));
    SB_LUT4 add_2747_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n53979), 
            .O(n8027[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n54295), 
            .O(n8287[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_19 (.CI(n54295), .I0(n3050), .I1(n2867), .CO(n54296));
    SB_CARRY add_2747_4 (.CI(n53979), .I0(n1840), .I1(n698), .CO(n53980));
    SB_LUT4 add_2757_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n54294), 
            .O(n8287[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_18 (.CI(n54294), .I0(n3051), .I1(n2754), .CO(n54295));
    SB_LUT4 add_2747_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n53978), 
            .O(n8027[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_3 (.CI(n53978), .I0(n1841), .I1(n858), .CO(n53979));
    SB_LUT4 i52287_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i52287_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 add_2757_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n54293), 
            .O(n8287[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_17 (.CI(n54293), .I0(n3052), .I1(n2638), .CO(n54294));
    SB_LUT4 add_2757_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n54292), 
            .O(n8287[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_16 (.CI(n54292), .I0(n3053), .I1(n2519), .CO(n54293));
    SB_LUT4 add_2757_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n54291), 
            .O(n8287[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2747_2_lut (.I0(n61837), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2757_15 (.CI(n54291), .I0(n3054), .I1(n2397), .CO(n54292));
    SB_LUT4 add_2757_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n54290), 
            .O(n8287[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53978));
    SB_CARRY add_2757_14 (.CI(n54290), .I0(n3055), .I1(n2272), .CO(n54291));
    SB_LUT4 add_2757_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n54289), 
            .O(n8287[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_13 (.CI(n54289), .I0(n3056), .I1(n2144), .CO(n54290));
    SB_LUT4 add_2757_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n54288), 
            .O(n8287[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_12 (.CI(n54288), .I0(n3057), .I1(n2013), .CO(n54289));
    SB_LUT4 add_2757_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n54287), 
            .O(n8287[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_11 (.CI(n54287), .I0(n3058), .I1(n1879), .CO(n54288));
    SB_LUT4 add_2757_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n54286), 
            .O(n8287[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_10 (.CI(n54286), .I0(n3059), .I1(n1742), .CO(n54287));
    SB_LUT4 i52367_4_lut (.I0(n23_adj_5199), .I1(n21_adj_5106), .I2(n19_adj_5105), 
            .I3(n17_adj_5202), .O(n69457));
    defparam i52367_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2757_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n54285), 
            .O(n8287[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_9 (.CI(n54285), .I0(n3060), .I1(n1602), .CO(n54286));
    SB_LUT4 add_2757_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n54284), 
            .O(n8287[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_8 (.CI(n54284), .I0(n3061), .I1(n1459), .CO(n54285));
    SB_LUT4 add_2757_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n54283), 
            .O(n8287[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_7 (.CI(n54283), .I0(n3062), .I1(n1460), .CO(n54284));
    SB_LUT4 add_2757_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n54282), 
            .O(n8287[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_6 (.CI(n54282), .I0(n3063), .I1(n1011), .CO(n54283));
    SB_LUT4 add_2757_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n54281), 
            .O(n8287[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_5 (.CI(n54281), .I0(n3064), .I1(n856), .CO(n54282));
    SB_LUT4 add_2757_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n54280), 
            .O(n8287[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_4 (.CI(n54280), .I0(n3065), .I1(n698), .CO(n54281));
    SB_LUT4 add_2757_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n54279), 
            .O(n8287[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_3 (.CI(n54279), .I0(n3066), .I1(n858), .CO(n54280));
    SB_LUT4 add_2757_2_lut (.I0(n61800), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63719)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2757_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54279));
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5204), .I1(baudrate[4]), 
            .I2(n43_adj_5168), .I3(GND_net), .O(n42_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54022_4_lut (.I0(n42_adj_5205), .I1(n38_adj_5203), .I2(n43_adj_5168), 
            .I3(n68741), .O(n71112));   // verilog/uart_rx.v(119[33:55])
    defparam i54022_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54023_3_lut (.I0(n71112), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n71113));   // verilog/uart_rx.v(119[33:55])
    defparam i54023_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i44772_1_lut (.I0(n25426), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61812));
    defparam i44772_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53741_3_lut (.I0(n71113), .I1(baudrate[6]), .I2(n1111), .I3(GND_net), 
            .O(n48_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam i53741_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52361_4_lut (.I0(n29_adj_5103), .I1(n27_adj_5102), .I2(n25_adj_5200), 
            .I3(n69457), .O(n69451));
    defparam i52361_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i44768_1_lut (.I0(n25429), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61808));
    defparam i44768_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(n63697), .I1(n48_adj_5206), .I2(GND_net), 
            .I3(GND_net), .O(n1267));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7923[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54018_3_lut (.I0(n34_adj_5207), .I1(baudrate[5]), .I2(n41_adj_5157), 
            .I3(GND_net), .O(n71108));   // verilog/uart_rx.v(119[33:55])
    defparam i54018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48183_1_lut (.I0(n65263), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61804));
    defparam i48183_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53940_4_lut (.I0(n35_adj_5113), .I1(n33_adj_5112), .I2(n31_adj_5111), 
            .I3(n69451), .O(n71030));
    defparam i53940_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54019_3_lut (.I0(n71108), .I1(baudrate[6]), .I2(n43_adj_5159), 
            .I3(GND_net), .O(n71109));   // verilog/uart_rx.v(119[33:55])
    defparam i54019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52631_4_lut (.I0(n43_adj_5159), .I1(n41_adj_5157), .I2(n39_adj_5158), 
            .I3(n68709), .O(n69721));
    defparam i52631_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36_adj_5209), .I1(baudrate[4]), 
            .I2(n39_adj_5158), .I3(GND_net), .O(n38_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53747_3_lut (.I0(n71109), .I1(baudrate[7]), .I2(n45_adj_5155), 
            .I3(GND_net), .O(n44_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam i53747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53359_4_lut (.I0(n44_adj_5211), .I1(n38_adj_5210), .I2(n45_adj_5155), 
            .I3(n69721), .O(n70449));   // verilog/uart_rx.v(119[33:55])
    defparam i53359_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53806_3_lut (.I0(n16_adj_5208), .I1(baudrate[13]), .I2(n39_adj_5097), 
            .I3(GND_net), .O(n70896));   // verilog/uart_rx.v(119[33:55])
    defparam i53806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53360_3_lut (.I0(n70449), .I1(baudrate[8]), .I2(n1408), .I3(GND_net), 
            .O(n48_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam i53360_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7923[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7949[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2756_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n54261), 
            .O(n8261[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2756_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n54260), 
            .O(n8261[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53807_3_lut (.I0(n70896), .I1(baudrate[14]), .I2(n41_adj_5095), 
            .I3(GND_net), .O(n70897));   // verilog/uart_rx.v(119[33:55])
    defparam i53807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2746_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n53943), 
            .O(n8001[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2746_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n53942), 
            .O(n8001[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_10 (.CI(n53942), .I0(n1694), .I1(n1879), .CO(n53943));
    SB_LUT4 i1_2_lut_adj_1040 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n64463));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'heeee;
    SB_LUT4 add_2746_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n53941), 
            .O(n8001[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_9 (.CI(n53941), .I0(n1695), .I1(n1742), .CO(n53942));
    SB_LUT4 add_2746_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n53940), 
            .O(n8001[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_8 (.CI(n53940), .I0(n1696), .I1(n1602), .CO(n53941));
    SB_LUT4 add_2746_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n53939), 
            .O(n8001[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_7 (.CI(n53939), .I0(n1697), .I1(n1459), .CO(n53940));
    SB_LUT4 add_2746_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n53938), 
            .O(n8001[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_6 (.CI(n53938), .I0(n1698), .I1(n1460), .CO(n53939));
    SB_LUT4 i53213_4_lut (.I0(n41_adj_5095), .I1(n39_adj_5097), .I2(n27_adj_5102), 
            .I3(n69453), .O(n70303));
    defparam i53213_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53790_3_lut (.I0(n22_adj_5213), .I1(baudrate[7]), .I2(n27_adj_5102), 
            .I3(GND_net), .O(n70880));   // verilog/uart_rx.v(119[33:55])
    defparam i53790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2746_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n53937), 
            .O(n8001[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_21 (.CI(n54260), .I0(n2939), .I1(n3084), .CO(n54261));
    SB_CARRY add_2746_5 (.CI(n53937), .I0(n1699), .I1(n1011), .CO(n53938));
    SB_LUT4 add_2746_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n53936), 
            .O(n8001[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_4 (.CI(n53936), .I0(n1700), .I1(n856), .CO(n53937));
    SB_LUT4 add_2746_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n53935), 
            .O(n8001[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_3 (.CI(n53935), .I0(n1701), .I1(n698), .CO(n53936));
    SB_LUT4 add_2746_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8001[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52696_3_lut (.I0(n70897), .I1(baudrate[15]), .I2(n43_adj_5094), 
            .I3(GND_net), .O(n69786));   // verilog/uart_rx.v(119[33:55])
    defparam i52696_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2746_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n53935));
    SB_LUT4 add_2756_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n54259), 
            .O(n8261[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_20 (.CI(n54259), .I0(n2940), .I1(n2977), .CO(n54260));
    SB_LUT4 add_2756_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n54258), 
            .O(n8261[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_19 (.CI(n54258), .I0(n2941), .I1(n2867), .CO(n54259));
    SB_LUT4 add_2756_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n54257), 
            .O(n8261[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54016_3_lut (.I0(n32_adj_5214), .I1(baudrate[5]), .I2(n39_adj_5212), 
            .I3(GND_net), .O(n71106));   // verilog/uart_rx.v(119[33:55])
    defparam i54016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54017_3_lut (.I0(n71106), .I1(baudrate[6]), .I2(n41_adj_5154), 
            .I3(GND_net), .O(n71107));   // verilog/uart_rx.v(119[33:55])
    defparam i54017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52623_4_lut (.I0(n41_adj_5154), .I1(n39_adj_5212), .I2(n37_adj_5153), 
            .I3(n68696), .O(n69713));
    defparam i52623_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2745_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n53908), 
            .O(n7975[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n53907), 
            .O(n7975[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_10 (.CI(n53907), .I0(n1553), .I1(n1742), .CO(n53908));
    SB_LUT4 add_2745_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n53906), 
            .O(n7975[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_9 (.CI(n53906), .I0(n1554), .I1(n1602), .CO(n53907));
    SB_LUT4 add_2745_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n53905), 
            .O(n7975[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53361_3_lut (.I0(n34_adj_5215), .I1(baudrate[4]), .I2(n37_adj_5153), 
            .I3(GND_net), .O(n70451));   // verilog/uart_rx.v(119[33:55])
    defparam i53361_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2745_8 (.CI(n53905), .I0(n1555), .I1(n1459), .CO(n53906));
    SB_LUT4 add_2745_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n53904), 
            .O(n7975[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_7 (.CI(n53904), .I0(n1556), .I1(n1460), .CO(n53905));
    SB_LUT4 add_2745_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n53903), 
            .O(n7975[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53751_3_lut (.I0(n71107), .I1(baudrate[7]), .I2(n43_adj_5151), 
            .I3(GND_net), .O(n70841));   // verilog/uart_rx.v(119[33:55])
    defparam i53751_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2745_6 (.CI(n53903), .I0(n1557), .I1(n1011), .CO(n53904));
    SB_LUT4 add_2745_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n53902), 
            .O(n7975[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_5 (.CI(n53902), .I0(n1558), .I1(n856), .CO(n53903));
    SB_LUT4 add_2745_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n53901), 
            .O(n7975[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_4 (.CI(n53901), .I0(n1559), .I1(n698), .CO(n53902));
    SB_LUT4 add_2745_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n53900), 
            .O(n7975[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54014_4_lut (.I0(n70841), .I1(n70451), .I2(n43_adj_5151), 
            .I3(n69713), .O(n71104));   // verilog/uart_rx.v(119[33:55])
    defparam i54014_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2745_3 (.CI(n53900), .I0(n1560), .I1(n858), .CO(n53901));
    SB_LUT4 add_2745_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7975[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53900));
    SB_LUT4 add_2744_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n53899), 
            .O(n7949[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8313[20]), .I3(n294[1]), .O(n41_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2744_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n53898), 
            .O(n7949[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_9 (.CI(n53898), .I0(n1409), .I1(n1602), .CO(n53899));
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8313[19]), .I3(n294[1]), .O(n39_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n53723), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2744_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n53897), 
            .O(n7949[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n63607), .I1(n25296), .I2(VCC_net), 
            .I3(n53722), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_8 (.CI(n53897), .I0(n1410), .I1(n1459), .CO(n53898));
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8313[14]), .I3(n294[1]), .O(n29_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_25 (.CI(n53722), .I0(n25296), .I1(VCC_net), 
            .CO(n53723));
    SB_LUT4 sub_38_add_2_24_lut (.I0(n63751), .I1(n65297), .I2(VCC_net), 
            .I3(n53721), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2744_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n53896), 
            .O(n7949[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_24 (.CI(n53721), .I0(n65297), .I1(VCC_net), 
            .CO(n53722));
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n53720), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_7 (.CI(n53896), .I0(n1411), .I1(n1460), .CO(n53897));
    SB_LUT4 i54015_3_lut (.I0(n71104), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n71105));   // verilog/uart_rx.v(119[33:55])
    defparam i54015_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY sub_38_add_2_23 (.CI(n53720), .I0(n294[21]), .I1(VCC_net), 
            .CO(n53721));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n63749), .I1(n294[20]), .I2(VCC_net), 
            .I3(n53719), .O(n63751)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2744_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n53895), 
            .O(n7949[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_22 (.CI(n53719), .I0(n294[20]), .I1(VCC_net), 
            .CO(n53720));
    SB_LUT4 sub_38_add_2_21_lut (.I0(n63747), .I1(n294[19]), .I2(VCC_net), 
            .I3(n53718), .O(n63749)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_6 (.CI(n53895), .I0(n1412), .I1(n1011), .CO(n53896));
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8313[15]), .I3(n294[1]), .O(n31_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2744_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n53894), 
            .O(n7949[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_5 (.CI(n53894), .I0(n1413), .I1(n856), .CO(n53895));
    SB_LUT4 add_2744_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n53893), 
            .O(n7949[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_4 (.CI(n53893), .I0(n1414), .I1(n698), .CO(n53894));
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8313[16]), .I3(n294[1]), .O(n33_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8313[17]), .I3(n294[1]), .O(n35_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_21 (.CI(n53718), .I0(n294[19]), .I1(VCC_net), 
            .CO(n53719));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n53717), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2744_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n53892), 
            .O(n7949[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n53717), .I0(n294[18]), .I1(VCC_net), 
            .CO(n53718));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n63745), .I1(n294[17]), .I2(VCC_net), 
            .I3(n53716), .O(n63747)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_3 (.CI(n53892), .I0(n1415), .I1(n858), .CO(n53893));
    SB_CARRY sub_38_add_2_19 (.CI(n53716), .I0(n294[17]), .I1(VCC_net), 
            .CO(n53717));
    SB_LUT4 sub_38_add_2_18_lut (.I0(n63743), .I1(n294[16]), .I2(VCC_net), 
            .I3(n53715), .O(n63745)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2744_2_lut (.I0(n61846), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_38_add_2_18 (.CI(n53715), .I0(n294[16]), .I1(VCC_net), 
            .CO(n53716));
    SB_LUT4 sub_38_add_2_17_lut (.I0(n63605), .I1(n294[15]), .I2(VCC_net), 
            .I3(n53714), .O(n63607)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53892));
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8313[18]), .I3(n294[1]), .O(n37_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 add_2743_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n53891), 
            .O(n7923[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n53890), 
            .O(n7923[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8313[11]), .I3(n294[1]), .O(n23_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2743_8 (.CI(n53890), .I0(n1262), .I1(n1459), .CO(n53891));
    SB_LUT4 add_2743_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n53889), 
            .O(n7923[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8313[12]), .I3(n294[1]), .O(n25_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8313[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8313[22]), .I3(n294[1]), .O(n45_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_17 (.CI(n53714), .I0(n294[15]), .I1(VCC_net), 
            .CO(n53715));
    SB_CARRY add_2743_7 (.CI(n53889), .I0(n1263), .I1(n1460), .CO(n53890));
    SB_LUT4 sub_38_add_2_16_lut (.I0(n63741), .I1(n294[14]), .I2(VCC_net), 
            .I3(n53713), .O(n63743)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2743_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n53888), 
            .O(n7923[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_16 (.CI(n53713), .I0(n294[14]), .I1(VCC_net), 
            .CO(n53714));
    SB_CARRY add_2743_6 (.CI(n53888), .I0(n1264), .I1(n1011), .CO(n53889));
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n53712), .O(n63741)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2743_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n53887), 
            .O(n7923[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53753_3_lut (.I0(n71105), .I1(baudrate[9]), .I2(n1552), .I3(GND_net), 
            .O(n48_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam i53753_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2743_5 (.CI(n53887), .I0(n1265), .I1(n856), .CO(n53888));
    SB_LUT4 add_2743_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n53886), 
            .O(n7923[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8313[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8313[8]), .I3(n294[1]), .O(n17_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY add_2743_4 (.CI(n53886), .I0(n1266), .I1(n698), .CO(n53887));
    SB_LUT4 add_2743_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n53885), 
            .O(n7923[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7949[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8313[10]), .I3(n294[1]), .O(n21_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_15 (.CI(n53712), .I0(n294[13]), .I1(VCC_net), 
            .CO(n53713));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n53711), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_3 (.CI(n53885), .I0(n1267), .I1(n858), .CO(n53886));
    SB_CARRY sub_38_add_2_14 (.CI(n53711), .I0(n294[12]), .I1(VCC_net), 
            .CO(n53712));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n53710), .O(n63605)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_2743_2_lut (.I0(n61850), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7975[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8313[5]), .I3(n294[1]), .O(n11_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_13 (.CI(n53710), .I0(n294[11]), .I1(VCC_net), 
            .CO(n53711));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n53709), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53885));
    SB_CARRY sub_38_add_2_12 (.CI(n53709), .I0(n294[10]), .I1(VCC_net), 
            .CO(n53710));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n53708), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n53708), .I0(n294[9]), .I1(VCC_net), 
            .CO(n53709));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n53707), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8313[6]), .I3(n294[1]), .O(n13_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_10 (.CI(n53707), .I0(n294[8]), .I1(VCC_net), 
            .CO(n53708));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n53706), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n64487));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8313[7]), .I3(n294[1]), .O(n15_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8313[13]), .I3(n294[1]), .O(n27_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_9 (.CI(n53706), .I0(n294[7]), .I1(VCC_net), 
            .CO(n53707));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n53705), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n53705), .I0(n294[6]), .I1(VCC_net), 
            .CO(n53706));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n53704), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n53704), .I0(n294[5]), .I1(VCC_net), 
            .CO(n53705));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n53703), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n53703), .I0(n294[4]), .I1(VCC_net), 
            .CO(n53704));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n53702), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8313[9]), .I3(n294[1]), .O(n19_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_5 (.CI(n53702), .I0(n294[3]), .I1(VCC_net), 
            .CO(n53703));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n53701), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8313[21]), .I3(n294[1]), .O(n43_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_CARRY sub_38_add_2_4 (.CI(n53701), .I0(n294[2]), .I1(VCC_net), 
            .CO(n53702));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n53700), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51915_4_lut (.I0(n27_adj_5232), .I1(n15_adj_5231), .I2(n13_adj_5230), 
            .I3(n11_adj_5229), .O(n69005));
    defparam i51915_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY sub_38_add_2_3 (.CI(n53700), .I0(n294[1]), .I1(VCC_net), 
            .CO(n53701));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n62613), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n62613), .I1(GND_net), 
            .CO(n53700));
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5235), .I1(baudrate[9]), 
            .I2(n31_adj_5111), .I3(GND_net), .O(n28_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51925_4_lut (.I0(n21_adj_5228), .I1(n19_adj_5233), .I2(n17_adj_5227), 
            .I3(n9), .O(n69015));
    defparam i51925_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5234), .I3(GND_net), .O(n16_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n64485));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'heeee;
    SB_LUT4 i51889_2_lut (.I0(n43_adj_5234), .I1(n19_adj_5233), .I2(GND_net), 
            .I3(GND_net), .O(n68979));
    defparam i51889_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5227), .I3(GND_net), .O(n8_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2742_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n53866), 
            .O(n7897[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2742_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n53865), 
            .O(n7897[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5237), .I1(baudrate[22]), 
            .I2(n45_adj_5225), .I3(GND_net), .O(n24_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2742_7 (.CI(n53865), .I0(n1112), .I1(n1460), .CO(n53866));
    SB_LUT4 add_2742_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n53864), 
            .O(n7897[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n64483));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'heeee;
    SB_CARRY add_2742_6 (.CI(n53864), .I0(n1113), .I1(n1011), .CO(n53865));
    SB_LUT4 add_2742_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n53863), 
            .O(n7897[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_5 (.CI(n53863), .I0(n1114), .I1(n856), .CO(n53864));
    SB_LUT4 add_2742_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n53862), 
            .O(n7897[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8313[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51948_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n69038));
    defparam i51948_3_lut.LUT_INIT = 16'hbebe;
    SB_CARRY add_2742_4 (.CI(n53862), .I0(n1115), .I1(n698), .CO(n53863));
    SB_LUT4 add_2742_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n53861), 
            .O(n7897[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_3 (.CI(n53861), .I0(n1116), .I1(n858), .CO(n53862));
    SB_LUT4 add_2742_2_lut (.I0(n61854), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2742_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n53861));
    SB_LUT4 i52899_4_lut (.I0(n13_adj_5230), .I1(n11_adj_5229), .I2(n9), 
            .I3(n69038), .O(n69989));
    defparam i52899_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52889_4_lut (.I0(n19_adj_5233), .I1(n17_adj_5227), .I2(n15_adj_5231), 
            .I3(n69989), .O(n69979));
    defparam i52889_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i54100_4_lut (.I0(n25_adj_5224), .I1(n23_adj_5223), .I2(n21_adj_5228), 
            .I3(n69979), .O(n71190));
    defparam i54100_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53443_4_lut (.I0(n31_adj_5219), .I1(n29_adj_5218), .I2(n27_adj_5232), 
            .I3(n71190), .O(n70533));
    defparam i53443_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54276_4_lut (.I0(n37_adj_5222), .I1(n35_adj_5221), .I2(n33_adj_5220), 
            .I3(n70533), .O(n71366));
    defparam i54276_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5220), .I3(GND_net), .O(n12_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63721), .I3(n48_adj_5241), .O(n4_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i53700_3_lut (.I0(n4_c), .I1(baudrate[13]), .I2(n27_adj_5232), 
            .I3(GND_net), .O(n70790));   // verilog/uart_rx.v(119[33:55])
    defparam i53700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53701_3_lut (.I0(n70790), .I1(baudrate[14]), .I2(n29_adj_5218), 
            .I3(GND_net), .O(n70791));   // verilog/uart_rx.v(119[33:55])
    defparam i53701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51909_2_lut (.I0(n33_adj_5220), .I1(n15_adj_5231), .I2(GND_net), 
            .I3(GND_net), .O(n68999));
    defparam i51909_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13_adj_5230), .I3(GND_net), .O(n10_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12_adj_5240), .I1(baudrate[17]), 
            .I2(n35_adj_5221), .I3(GND_net), .O(n30_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51911_4_lut (.I0(n33_adj_5220), .I1(n31_adj_5219), .I2(n29_adj_5218), 
            .I3(n69005), .O(n69001));
    defparam i51911_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54185_4_lut (.I0(n28_adj_5236), .I1(n18_adj_5244), .I2(n31_adj_5111), 
            .I3(n69446), .O(n71275));   // verilog/uart_rx.v(119[33:55])
    defparam i54185_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54221_4_lut (.I0(n30_adj_5243), .I1(n10_adj_5242), .I2(n35_adj_5221), 
            .I3(n68999), .O(n71311));   // verilog/uart_rx.v(119[33:55])
    defparam i54221_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52758_3_lut (.I0(n70791), .I1(baudrate[15]), .I2(n31_adj_5219), 
            .I3(GND_net), .O(n69848));   // verilog/uart_rx.v(119[33:55])
    defparam i52758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54420_4_lut (.I0(n69848), .I1(n71311), .I2(n35_adj_5221), 
            .I3(n69001), .O(n71510));   // verilog/uart_rx.v(119[33:55])
    defparam i54420_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54421_3_lut (.I0(n71510), .I1(baudrate[18]), .I2(n37_adj_5222), 
            .I3(GND_net), .O(n71511));   // verilog/uart_rx.v(119[33:55])
    defparam i54421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(n64529), .I1(n64485), .I2(n64487), 
            .I3(baudrate[11]), .O(n64515));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(n64515), .I1(n64517), .I2(n64505), 
            .I3(n64461), .O(n25437));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'hfffe;
    SB_LUT4 i53702_3_lut (.I0(n6_adj_5245), .I1(baudrate[10]), .I2(n21_adj_5228), 
            .I3(GND_net), .O(n70792));   // verilog/uart_rx.v(119[33:55])
    defparam i53702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53703_3_lut (.I0(n70792), .I1(baudrate[11]), .I2(n23_adj_5223), 
            .I3(GND_net), .O(n70793));   // verilog/uart_rx.v(119[33:55])
    defparam i53703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51891_4_lut (.I0(n43_adj_5234), .I1(n25_adj_5224), .I2(n23_adj_5223), 
            .I3(n69015), .O(n68981));
    defparam i51891_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53802_4_lut (.I0(n24_adj_5239), .I1(n8_adj_5238), .I2(n45_adj_5225), 
            .I3(n68979), .O(n70892));   // verilog/uart_rx.v(119[33:55])
    defparam i53802_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2756_18 (.CI(n54257), .I0(n2942), .I1(n2754), .CO(n54258));
    SB_LUT4 add_2756_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n54256), 
            .O(n8261[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52756_3_lut (.I0(n70793), .I1(baudrate[12]), .I2(n25_adj_5224), 
            .I3(GND_net), .O(n69846));   // verilog/uart_rx.v(119[33:55])
    defparam i52756_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_17 (.CI(n54256), .I0(n2943), .I1(n2638), .CO(n54257));
    SB_LUT4 add_2756_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n54255), 
            .O(n8261[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_16 (.CI(n54255), .I0(n2944), .I1(n2519), .CO(n54256));
    SB_LUT4 add_2756_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n54254), 
            .O(n8261[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54335_3_lut (.I0(n71511), .I1(baudrate[19]), .I2(n39_adj_5217), 
            .I3(GND_net), .O(n71425));   // verilog/uart_rx.v(119[33:55])
    defparam i54335_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_15 (.CI(n54254), .I0(n2945), .I1(n2397), .CO(n54255));
    SB_LUT4 add_2756_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n54253), 
            .O(n8261[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51899_4_lut (.I0(n43_adj_5234), .I1(n41_adj_5216), .I2(n39_adj_5217), 
            .I3(n71366), .O(n68989));
    defparam i51899_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54266_4_lut (.I0(n69846), .I1(n70892), .I2(n45_adj_5225), 
            .I3(n68981), .O(n71356));   // verilog/uart_rx.v(119[33:55])
    defparam i54266_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2756_14 (.CI(n54253), .I0(n2946), .I1(n2272), .CO(n54254));
    SB_LUT4 add_2756_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n54252), 
            .O(n8261[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_13 (.CI(n54252), .I0(n2947), .I1(n2144), .CO(n54253));
    SB_LUT4 add_2756_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n54251), 
            .O(n8261[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52764_3_lut (.I0(n71425), .I1(baudrate[20]), .I2(n41_adj_5216), 
            .I3(GND_net), .O(n69854));   // verilog/uart_rx.v(119[33:55])
    defparam i52764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n63677));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'heeee;
    SB_CARRY add_2756_12 (.CI(n54251), .I0(n2948), .I1(n2013), .CO(n54252));
    SB_LUT4 add_2756_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n54250), 
            .O(n8261[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54186_3_lut (.I0(n71275), .I1(baudrate[10]), .I2(n33_adj_5112), 
            .I3(GND_net), .O(n71276));   // verilog/uart_rx.v(119[33:55])
    defparam i54186_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_11 (.CI(n54250), .I0(n2949), .I1(n1879), .CO(n54251));
    SB_LUT4 add_2756_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n54249), 
            .O(n8261[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8313[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2756_10 (.CI(n54249), .I0(n2950), .I1(n1742), .CO(n54250));
    SB_LUT4 add_2756_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n54248), 
            .O(n8261[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_9 (.CI(n54248), .I0(n2951), .I1(n1602), .CO(n54249));
    SB_LUT4 add_2756_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n54247), 
            .O(n8261[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54268_4_lut (.I0(n69854), .I1(n71356), .I2(n45_adj_5225), 
            .I3(n68989), .O(n71358));   // verilog/uart_rx.v(119[33:55])
    defparam i54268_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2756_8 (.CI(n54247), .I0(n2952), .I1(n1459), .CO(n54248));
    SB_LUT4 add_2756_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n54246), 
            .O(n8261[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_7 (.CI(n54246), .I0(n2953), .I1(n1460), .CO(n54247));
    SB_LUT4 add_2756_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n54245), 
            .O(n8261[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54073_3_lut (.I0(n71276), .I1(baudrate[11]), .I2(n35_adj_5113), 
            .I3(GND_net), .O(n71163));   // verilog/uart_rx.v(119[33:55])
    defparam i54073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(n64623), .I1(n64487), .I2(n63677), 
            .I3(n64485), .O(n63685));
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'hfffe;
    SB_CARRY add_2756_6 (.CI(n54245), .I0(n2954), .I1(n1011), .CO(n54246));
    SB_LUT4 add_2756_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n54244), 
            .O(n8261[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_5 (.CI(n54244), .I0(n2955), .I1(n856), .CO(n54245));
    SB_LUT4 add_2756_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n54243), 
            .O(n8261[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54648_4_lut (.I0(n63685), .I1(n71358), .I2(baudrate[23]), 
            .I3(n3253), .O(n62613));   // verilog/uart_rx.v(119[33:55])
    defparam i54648_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2756_4 (.CI(n54243), .I0(n2956), .I1(n698), .CO(n54244));
    SB_LUT4 add_2756_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n54242), 
            .O(n8261[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_3 (.CI(n54242), .I0(n2957), .I1(n858), .CO(n54243));
    SB_LUT4 add_2756_2_lut (.I0(n61804), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2756_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54242));
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23475_rep_4_2_lut (.I0(n7975[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n61840));   // verilog/uart_rx.v(119[33:55])
    defparam i23475_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2755_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n54232), 
            .O(n8235[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2755_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n54231), 
            .O(n8235[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_20 (.CI(n54231), .I0(n2828), .I1(n2977), .CO(n54232));
    SB_LUT4 add_2755_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n54230), 
            .O(n8235[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_19 (.CI(n54230), .I0(n2829), .I1(n2867), .CO(n54231));
    SB_LUT4 add_2755_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n54229), 
            .O(n8235[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_18 (.CI(n54229), .I0(n2830), .I1(n2754), .CO(n54230));
    SB_LUT4 add_2755_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n54228), 
            .O(n8235[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n61840), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i54012_3_lut (.I0(n32_adj_5254), .I1(baudrate[6]), .I2(n39_adj_5148), 
            .I3(GND_net), .O(n71102));   // verilog/uart_rx.v(119[33:55])
    defparam i54012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_17 (.CI(n54228), .I0(n2831), .I1(n2638), .CO(n54229));
    SB_LUT4 add_2755_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n54227), 
            .O(n8235[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_16 (.CI(n54227), .I0(n2832), .I1(n2519), .CO(n54228));
    SB_LUT4 add_2755_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n54226), 
            .O(n8235[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54013_3_lut (.I0(n71102), .I1(baudrate[7]), .I2(n41_adj_5150), 
            .I3(GND_net), .O(n71103));   // verilog/uart_rx.v(119[33:55])
    defparam i54013_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2755_15 (.CI(n54226), .I0(n2833), .I1(n2397), .CO(n54227));
    SB_LUT4 add_2755_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n54225), 
            .O(n8235[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_14 (.CI(n54225), .I0(n2834), .I1(n2272), .CO(n54226));
    SB_LUT4 add_2755_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n54224), 
            .O(n8235[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52543_4_lut (.I0(n41_adj_5150), .I1(n39_adj_5148), .I2(n37_adj_5149), 
            .I3(n68673), .O(n69633));
    defparam i52543_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2755_13 (.CI(n54224), .I0(n2835), .I1(n2144), .CO(n54225));
    SB_LUT4 add_2755_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n54223), 
            .O(n8235[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_12 (.CI(n54223), .I0(n2836), .I1(n2013), .CO(n54224));
    SB_LUT4 add_2755_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n54222), 
            .O(n8235[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_11 (.CI(n54222), .I0(n2837), .I1(n1879), .CO(n54223));
    SB_LUT4 add_2755_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n54221), 
            .O(n8235[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_10 (.CI(n54221), .I0(n2838), .I1(n1742), .CO(n54222));
    SB_LUT4 add_2755_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n54220), 
            .O(n8235[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_9 (.CI(n54220), .I0(n2839), .I1(n1602), .CO(n54221));
    SB_LUT4 add_2755_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n54219), 
            .O(n8235[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_8 (.CI(n54219), .I0(n2840), .I1(n1459), .CO(n54220));
    SB_LUT4 add_2755_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n54218), 
            .O(n8235[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53217_4_lut (.I0(n41_adj_5095), .I1(n39_adj_5097), .I2(n37_adj_5093), 
            .I3(n71030), .O(n70307));
    defparam i53217_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2755_7 (.CI(n54218), .I0(n2841), .I1(n1460), .CO(n54219));
    SB_LUT4 add_2755_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n54217), 
            .O(n8235[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_6 (.CI(n54217), .I0(n2842), .I1(n1011), .CO(n54218));
    SB_LUT4 add_2755_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n54216), 
            .O(n8235[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_5 (.CI(n54216), .I0(n2843), .I1(n856), .CO(n54217));
    SB_LUT4 add_2755_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n54215), 
            .O(n8235[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_4 (.CI(n54215), .I0(n2844), .I1(n698), .CO(n54216));
    SB_LUT4 add_2755_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n54214), 
            .O(n8235[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2755_3 (.CI(n54214), .I0(n2845), .I1(n858), .CO(n54215));
    SB_LUT4 add_2755_2_lut (.I0(n61808), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63715)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2755_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54214));
    SB_LUT4 i53363_3_lut (.I0(n34_adj_5262), .I1(baudrate[5]), .I2(n37_adj_5149), 
            .I3(GND_net), .O(n70453));   // verilog/uart_rx.v(119[33:55])
    defparam i53363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51984_4_lut (.I0(n29_adj_5261), .I1(n17_adj_5260), .I2(n15_adj_5259), 
            .I3(n13_adj_5258), .O(n69074));
    defparam i51984_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53755_3_lut (.I0(n71103), .I1(baudrate[8]), .I2(n43_adj_5147), 
            .I3(GND_net), .O(n70845));   // verilog/uart_rx.v(119[33:55])
    defparam i53755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54010_4_lut (.I0(n70845), .I1(n70453), .I2(n43_adj_5147), 
            .I3(n69633), .O(n71100));   // verilog/uart_rx.v(119[33:55])
    defparam i54010_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52957_4_lut (.I0(n11_adj_5256), .I1(n9_adj_5252), .I2(n3171), 
            .I3(baudrate[2]), .O(n70047));
    defparam i52957_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i53487_4_lut (.I0(n17_adj_5260), .I1(n15_adj_5259), .I2(n13_adj_5258), 
            .I3(n70047), .O(n70577));
    defparam i53487_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53485_4_lut (.I0(n23_adj_5255), .I1(n21_adj_5253), .I2(n19_adj_5257), 
            .I3(n70577), .O(n70575));
    defparam i53485_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51988_4_lut (.I0(n29_adj_5261), .I1(n27_adj_5251), .I2(n25_adj_5250), 
            .I3(n70575), .O(n69078));
    defparam i51988_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53804_4_lut (.I0(n69786), .I1(n70880), .I2(n43_adj_5094), 
            .I3(n70303), .O(n70894));   // verilog/uart_rx.v(119[33:55])
    defparam i53804_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2754_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n54197), 
            .O(n8209[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2754_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n54196), 
            .O(n8209[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_19 (.CI(n54196), .I0(n2714), .I1(n2867), .CO(n54197));
    SB_LUT4 add_2754_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n54195), 
            .O(n8209[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53708_3_lut (.I0(n6_adj_5263), .I1(baudrate[13]), .I2(n29_adj_5261), 
            .I3(GND_net), .O(n70798));   // verilog/uart_rx.v(119[33:55])
    defparam i53708_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_18 (.CI(n54195), .I0(n2715), .I1(n2754), .CO(n54196));
    SB_LUT4 add_2754_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n54194), 
            .O(n8209[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_17 (.CI(n54194), .I0(n2716), .I1(n2638), .CO(n54195));
    SB_LUT4 add_2754_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n54193), 
            .O(n8209[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54011_3_lut (.I0(n71100), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n71101));   // verilog/uart_rx.v(119[33:55])
    defparam i54011_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2754_16 (.CI(n54193), .I0(n2717), .I1(n2519), .CO(n54194));
    SB_LUT4 add_2754_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n54192), 
            .O(n8209[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_15 (.CI(n54192), .I0(n2718), .I1(n2397), .CO(n54193));
    SB_LUT4 add_2754_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n54191), 
            .O(n8209[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_14 (.CI(n54191), .I0(n2719), .I1(n2272), .CO(n54192));
    SB_LUT4 add_2754_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n54190), 
            .O(n8209[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_13 (.CI(n54190), .I0(n2720), .I1(n2144), .CO(n54191));
    SB_LUT4 add_2754_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n54189), 
            .O(n8209[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_12 (.CI(n54189), .I0(n2721), .I1(n2013), .CO(n54190));
    SB_LUT4 add_2754_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n54188), 
            .O(n8209[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_11 (.CI(n54188), .I0(n2722), .I1(n1879), .CO(n54189));
    SB_LUT4 add_2754_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n54187), 
            .O(n8209[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53757_3_lut (.I0(n71101), .I1(baudrate[10]), .I2(n1693), 
            .I3(GND_net), .O(n48_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam i53757_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2754_10 (.CI(n54187), .I0(n2723), .I1(n1742), .CO(n54188));
    SB_LUT4 add_2754_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n54186), 
            .O(n8209[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5264), .I1(baudrate[17]), 
            .I2(n37_adj_5248), .I3(GND_net), .O(n32_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_9 (.CI(n54186), .I0(n2724), .I1(n1602), .CO(n54187));
    SB_LUT4 add_2754_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n54185), 
            .O(n8209[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52694_3_lut (.I0(n71163), .I1(baudrate[12]), .I2(n37_adj_5093), 
            .I3(GND_net), .O(n69784));   // verilog/uart_rx.v(119[33:55])
    defparam i52694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53709_3_lut (.I0(n70798), .I1(baudrate[14]), .I2(n31_adj_5247), 
            .I3(GND_net), .O(n70799));   // verilog/uart_rx.v(119[33:55])
    defparam i53709_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_8 (.CI(n54185), .I0(n2725), .I1(n1459), .CO(n54186));
    SB_LUT4 add_2754_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n54184), 
            .O(n8209[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54350_4_lut (.I0(n69784), .I1(n70894), .I2(n43_adj_5094), 
            .I3(n70307), .O(n71440));   // verilog/uart_rx.v(119[33:55])
    defparam i54350_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2754_7 (.CI(n54184), .I0(n2726), .I1(n1460), .CO(n54185));
    SB_LUT4 add_2754_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n54183), 
            .O(n8209[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54351_3_lut (.I0(n71440), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n71441));   // verilog/uart_rx.v(119[33:55])
    defparam i54351_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51970_4_lut (.I0(n35_adj_5249), .I1(n33_adj_5246), .I2(n31_adj_5247), 
            .I3(n69074), .O(n69060));
    defparam i51970_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2754_6 (.CI(n54183), .I0(n2727), .I1(n1011), .CO(n54184));
    SB_LUT4 add_2754_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n54182), 
            .O(n8209[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54215_4_lut (.I0(n32_adj_5265), .I1(n12_adj_5266), .I2(n37_adj_5248), 
            .I3(n69056), .O(n71305));   // verilog/uart_rx.v(119[33:55])
    defparam i54215_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2754_5 (.CI(n54182), .I0(n2728), .I1(n856), .CO(n54183));
    SB_LUT4 add_2754_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n54181), 
            .O(n8209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n54585), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52744_3_lut (.I0(n70799), .I1(baudrate[15]), .I2(n33_adj_5246), 
            .I3(GND_net), .O(n69834));   // verilog/uart_rx.v(119[33:55])
    defparam i52744_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_4 (.CI(n54181), .I0(n2729), .I1(n698), .CO(n54182));
    SB_LUT4 add_2754_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n54180), 
            .O(n8209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n54584), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_3 (.CI(n54180), .I0(n2730), .I1(n858), .CO(n54181));
    SB_LUT4 add_2754_2_lut (.I0(n61812), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY r_Clock_Count_2053_add_4_8 (.CI(n54584), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n54585));
    SB_LUT4 i53710_3_lut (.I0(n8_adj_5267), .I1(baudrate[10]), .I2(n23_adj_5255), 
            .I3(GND_net), .O(n70800));   // verilog/uart_rx.v(119[33:55])
    defparam i53710_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54180));
    SB_LUT4 r_Clock_Count_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n54583), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_7 (.CI(n54583), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n54584));
    SB_LUT4 r_Clock_Count_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n54582), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_6 (.CI(n54582), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n54583));
    SB_LUT4 i53711_3_lut (.I0(n70800), .I1(baudrate[11]), .I2(n25_adj_5250), 
            .I3(GND_net), .O(n70801));   // verilog/uart_rx.v(119[33:55])
    defparam i53711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n54581), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_5 (.CI(n54581), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n54582));
    SB_LUT4 r_Clock_Count_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n54580), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_4 (.CI(n54580), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n54581));
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7975[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n54579), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_3 (.CI(n54579), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n54580));
    SB_LUT4 r_Clock_Count_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n54579));
    SB_LUT4 i52945_4_lut (.I0(n25_adj_5250), .I1(n23_adj_5255), .I2(n21_adj_5253), 
            .I3(n69086), .O(n70035));
    defparam i52945_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53800_3_lut (.I0(n10_adj_5268), .I1(baudrate[9]), .I2(n21_adj_5253), 
            .I3(GND_net), .O(n70890));   // verilog/uart_rx.v(119[33:55])
    defparam i53800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52742_3_lut (.I0(n70801), .I1(baudrate[12]), .I2(n27_adj_5251), 
            .I3(GND_net), .O(n69832));   // verilog/uart_rx.v(119[33:55])
    defparam i52742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53886_4_lut (.I0(n35_adj_5249), .I1(n33_adj_5246), .I2(n31_adj_5247), 
            .I3(n69078), .O(n70976));
    defparam i53886_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54418_4_lut (.I0(n69834), .I1(n71305), .I2(n37_adj_5248), 
            .I3(n69060), .O(n71508));   // verilog/uart_rx.v(119[33:55])
    defparam i54418_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54000_4_lut (.I0(n69832), .I1(n70890), .I2(n27_adj_5251), 
            .I3(n70035), .O(n71090));   // verilog/uart_rx.v(119[33:55])
    defparam i54000_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54466_4_lut (.I0(n71090), .I1(n71508), .I2(n37_adj_5248), 
            .I3(n70976), .O(n71556));   // verilog/uart_rx.v(119[33:55])
    defparam i54466_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8001[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54467_3_lut (.I0(n71556), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n71557));   // verilog/uart_rx.v(119[33:55])
    defparam i54467_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8027[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54463_3_lut (.I0(n71557), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n71553));   // verilog/uart_rx.v(119[33:55])
    defparam i54463_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54251_3_lut (.I0(n71553), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n71341));   // verilog/uart_rx.v(119[33:55])
    defparam i54251_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54252_3_lut (.I0(n71341), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n71342));   // verilog/uart_rx.v(119[33:55])
    defparam i54252_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52754_3_lut (.I0(n71342), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam i52754_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2753_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n54156), 
            .O(n8183[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2753_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n54155), 
            .O(n8183[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_18 (.CI(n54155), .I0(n2597), .I1(n2754), .CO(n54156));
    SB_LUT4 add_2753_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n54154), 
            .O(n8183[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_17 (.CI(n54154), .I0(n2598), .I1(n2638), .CO(n54155));
    SB_LUT4 add_2753_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n54153), 
            .O(n8183[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_16 (.CI(n54153), .I0(n2599), .I1(n2519), .CO(n54154));
    SB_LUT4 add_2753_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n54152), 
            .O(n8183[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_15 (.CI(n54152), .I0(n2600), .I1(n2397), .CO(n54153));
    SB_LUT4 add_2753_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n54151), 
            .O(n8183[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_14 (.CI(n54151), .I0(n2601), .I1(n2272), .CO(n54152));
    SB_LUT4 add_2753_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n54150), 
            .O(n8183[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_13 (.CI(n54150), .I0(n2602), .I1(n2144), .CO(n54151));
    SB_LUT4 add_2753_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n54149), 
            .O(n8183[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_12 (.CI(n54149), .I0(n2603), .I1(n2013), .CO(n54150));
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n54148), 
            .O(n8183[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_11 (.CI(n54148), .I0(n2604), .I1(n1879), .CO(n54149));
    SB_LUT4 add_2753_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n54147), 
            .O(n8183[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_10 (.CI(n54147), .I0(n2605), .I1(n1742), .CO(n54148));
    SB_LUT4 add_2753_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n54146), 
            .O(n8183[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_9 (.CI(n54146), .I0(n2606), .I1(n1602), .CO(n54147));
    SB_LUT4 add_2753_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n54145), 
            .O(n8183[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_8 (.CI(n54145), .I0(n2607), .I1(n1459), .CO(n54146));
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n54144), 
            .O(n8183[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_7 (.CI(n54144), .I0(n2608), .I1(n1460), .CO(n54145));
    SB_LUT4 add_2753_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n54143), 
            .O(n8183[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_6 (.CI(n54143), .I0(n2609), .I1(n1011), .CO(n54144));
    SB_LUT4 add_2753_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n54142), 
            .O(n8183[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_5 (.CI(n54142), .I0(n2610), .I1(n856), .CO(n54143));
    SB_LUT4 add_2753_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n54141), 
            .O(n8183[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_4 (.CI(n54141), .I0(n2611), .I1(n698), .CO(n54142));
    SB_LUT4 i51537_4_lut (.I0(n33_adj_5271), .I1(n31_adj_5270), .I2(n29_adj_5269), 
            .I3(n27_adj_5272), .O(n68627));
    defparam i51537_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2753_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n54140), 
            .O(n8183[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_3 (.CI(n54140), .I0(n2612), .I1(n858), .CO(n54141));
    SB_LUT4 add_2753_2_lut (.I0(n61816), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2753_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54140));
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5273), .I1(baudrate[9]), 
            .I2(n41_adj_5109), .I3(GND_net), .O(n38_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8157[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47948_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25423), .I3(baudrate[15]), .O(n65022));
    defparam i47948_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47947_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25423), .I3(GND_net), .O(n61824));
    defparam i47947_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i54002_3_lut (.I0(n26_adj_5275), .I1(baudrate[5]), .I2(n33_adj_5271), 
            .I3(GND_net), .O(n71092));   // verilog/uart_rx.v(119[33:55])
    defparam i54002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54003_3_lut (.I0(n71092), .I1(baudrate[6]), .I2(n35_adj_5107), 
            .I3(GND_net), .O(n71093));   // verilog/uart_rx.v(119[33:55])
    defparam i54003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54558_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25423), .I3(n48_adj_5134), .O(n294[8]));
    defparam i54558_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8183[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n54112), 
            .O(n8157[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2752_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n54111), 
            .O(n8157[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_17 (.CI(n54111), .I0(n2477), .I1(n2638), .CO(n54112));
    SB_LUT4 add_2752_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n54110), 
            .O(n8157[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_16 (.CI(n54110), .I0(n2478), .I1(n2519), .CO(n54111));
    SB_LUT4 add_2752_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n54109), 
            .O(n8157[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_15 (.CI(n54109), .I0(n2479), .I1(n2397), .CO(n54110));
    SB_LUT4 add_2752_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n54108), 
            .O(n8157[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_14 (.CI(n54108), .I0(n2480), .I1(n2272), .CO(n54109));
    SB_LUT4 add_2752_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n54107), 
            .O(n8157[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_13 (.CI(n54107), .I0(n2481), .I1(n2144), .CO(n54108));
    SB_LUT4 add_2752_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n54106), 
            .O(n8157[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_12 (.CI(n54106), .I0(n2482), .I1(n2013), .CO(n54107));
    SB_LUT4 add_2752_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n54105), 
            .O(n8157[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_11 (.CI(n54105), .I0(n2483), .I1(n1879), .CO(n54106));
    SB_LUT4 add_2752_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n54104), 
            .O(n8157[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51531_4_lut (.I0(n39_adj_5110), .I1(n37_adj_5108), .I2(n35_adj_5107), 
            .I3(n68627), .O(n68621));
    defparam i51531_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2752_10 (.CI(n54104), .I0(n2484), .I1(n1742), .CO(n54105));
    SB_LUT4 add_2752_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n54103), 
            .O(n8157[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_9 (.CI(n54103), .I0(n2485), .I1(n1602), .CO(n54104));
    SB_LUT4 add_2752_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n54102), 
            .O(n8157[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_8 (.CI(n54102), .I0(n2486), .I1(n1459), .CO(n54103));
    SB_LUT4 add_2752_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n54101), 
            .O(n8157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_7 (.CI(n54101), .I0(n2487), .I1(n1460), .CO(n54102));
    SB_LUT4 i54315_4_lut (.I0(n38_adj_5274), .I1(n28_adj_5276), .I2(n41_adj_5109), 
            .I3(n68619), .O(n71405));   // verilog/uart_rx.v(119[33:55])
    defparam i54315_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2752_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n54100), 
            .O(n8157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_6 (.CI(n54100), .I0(n2488), .I1(n1011), .CO(n54101));
    SB_LUT4 add_2752_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n54099), 
            .O(n8157[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_5 (.CI(n54099), .I0(n2489), .I1(n856), .CO(n54100));
    SB_LUT4 add_2752_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n54098), 
            .O(n8157[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_4 (.CI(n54098), .I0(n2490), .I1(n698), .CO(n54099));
    SB_LUT4 add_2752_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n54097), 
            .O(n8157[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_3 (.CI(n54097), .I0(n2491), .I1(n858), .CO(n54098));
    SB_LUT4 i53763_3_lut (.I0(n71093), .I1(baudrate[7]), .I2(n37_adj_5108), 
            .I3(GND_net), .O(n70853));   // verilog/uart_rx.v(119[33:55])
    defparam i53763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_2_lut (.I0(n61820), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n63709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2752_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n54097));
    SB_LUT4 i54452_4_lut (.I0(n70853), .I1(n71405), .I2(n41_adj_5109), 
            .I3(n68621), .O(n71542));   // verilog/uart_rx.v(119[33:55])
    defparam i54452_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54453_3_lut (.I0(n71542), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n71543));   // verilog/uart_rx.v(119[33:55])
    defparam i54453_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54413_3_lut (.I0(n71543), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n71503));   // verilog/uart_rx.v(119[33:55])
    defparam i54413_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54347_3_lut (.I0(n71503), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam i54347_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8027[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8053[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8209[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48104_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n65185));
    defparam i48104_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n64447));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48186_2_lut_3_lut_4_lut (.I0(baudrate[7]), .I1(n65259), .I2(baudrate[5]), 
            .I3(baudrate[6]), .O(n65267));
    defparam i48186_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n64533));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n64535));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n64529));
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n64531));
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8235[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n64241));
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n64537));
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n64489));
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8235[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1055 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n64539));
    defparam i1_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 i48179_1_lut (.I0(n65259), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61850));
    defparam i48179_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1056 (.I0(n64489), .I1(n64537), .I2(n64241), 
            .I3(GND_net), .O(n64547));
    defparam i1_3_lut_adj_1056.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1057 (.I0(n64547), .I1(n64543), .I2(n64545), 
            .I3(n64539), .O(n25411));
    defparam i1_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48206_4_lut (.I0(n65263), .I1(n65116), .I2(n61539), .I3(baudrate[4]), 
            .O(n65287));
    defparam i48206_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54725_4_lut (.I0(n65235), .I1(n65069), .I2(n65287), .I3(n65067), 
            .O(n65297));
    defparam i54725_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51497_4_lut (.I0(n33_adj_5104), .I1(n31_adj_5101), .I2(n29_adj_5100), 
            .I3(n27_adj_5280), .O(n68587));
    defparam i51497_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5281), .I1(baudrate[10]), 
            .I2(n41_adj_5098), .I3(GND_net), .O(n38_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23484_rep_3_2_lut (.I0(n8053[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n61831));   // verilog/uart_rx.v(119[33:55])
    defparam i23484_rep_3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n61831), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54054_3_lut (.I0(n26_adj_5283), .I1(baudrate[6]), .I2(n33_adj_5104), 
            .I3(GND_net), .O(n71144));   // verilog/uart_rx.v(119[33:55])
    defparam i54054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54055_3_lut (.I0(n71144), .I1(baudrate[7]), .I2(n35_adj_5096), 
            .I3(GND_net), .O(n71145));   // verilog/uart_rx.v(119[33:55])
    defparam i54055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51485_4_lut (.I0(n39_adj_5099), .I1(n37_adj_5092), .I2(n35_adj_5096), 
            .I3(n68587), .O(n68575));
    defparam i51485_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54317_4_lut (.I0(n38_adj_5282), .I1(n28_adj_5285), .I2(n41_adj_5098), 
            .I3(n68573), .O(n71407));   // verilog/uart_rx.v(119[33:55])
    defparam i54317_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i53767_3_lut (.I0(n71145), .I1(baudrate[8]), .I2(n37_adj_5092), 
            .I3(GND_net), .O(n70857));   // verilog/uart_rx.v(119[33:55])
    defparam i53767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54454_4_lut (.I0(n70857), .I1(n71407), .I2(n41_adj_5098), 
            .I3(n68575), .O(n71544));   // verilog/uart_rx.v(119[33:55])
    defparam i54454_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54455_3_lut (.I0(n71544), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n71545));   // verilog/uart_rx.v(119[33:55])
    defparam i54455_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54411_3_lut (.I0(n71545), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n71501));   // verilog/uart_rx.v(119[33:55])
    defparam i54411_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48106_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n65187));
    defparam i48106_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i54536_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n65231), .I3(n48_adj_5226), .O(n294[14]));
    defparam i54536_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48177_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n65231), .I3(baudrate[9]), .O(n61846));
    defparam i48177_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54349_3_lut (.I0(n71501), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i54349_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8053[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54547_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n65022), .I3(n48_adj_5277), .O(n294[11]));
    defparam i54547_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48182_4_lut (.I0(n65187), .I1(n64529), .I2(n65185), .I3(n64483), 
            .O(n65263));
    defparam i48182_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52103_4_lut (.I0(n33_adj_5055), .I1(n21_adj_5284), .I2(n19_adj_5279), 
            .I3(n17_adj_5278), .O(n69193));
    defparam i52103_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53085_4_lut (.I0(n15_adj_5054), .I1(n13_adj_5053), .I2(n2956), 
            .I3(baudrate[2]), .O(n70175));
    defparam i53085_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i48150_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n65022), .I3(baudrate[12]), .O(n65231));
    defparam i48150_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8079[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8105[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53545_4_lut (.I0(n21_adj_5284), .I1(n19_adj_5279), .I2(n17_adj_5278), 
            .I3(n70175), .O(n70635));
    defparam i53545_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i53539_4_lut (.I0(n27_adj_5051), .I1(n25_adj_5050), .I2(n23_adj_5049), 
            .I3(n70635), .O(n70629));
    defparam i53539_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52107_4_lut (.I0(n33_adj_5055), .I1(n31_adj_5048), .I2(n29_adj_5047), 
            .I3(n70629), .O(n69197));
    defparam i52107_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5286));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53728_3_lut (.I0(n10_adj_5286), .I1(baudrate[13]), .I2(n33_adj_5055), 
            .I3(GND_net), .O(n70818));   // verilog/uart_rx.v(119[33:55])
    defparam i53728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53729_3_lut (.I0(n70818), .I1(baudrate[14]), .I2(n35_adj_5027), 
            .I3(GND_net), .O(n70819));   // verilog/uart_rx.v(119[33:55])
    defparam i53729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5287), .I1(baudrate[17]), 
            .I2(n41), .I3(GND_net), .O(n36_adj_5288));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52096_4_lut (.I0(n39_adj_5052), .I1(n37_adj_5026), .I2(n35_adj_5027), 
            .I3(n69193), .O(n69186));
    defparam i52096_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54209_4_lut (.I0(n36_adj_5288), .I1(n16_adj_5289), .I2(n41), 
            .I3(n69182), .O(n71299));   // verilog/uart_rx.v(119[33:55])
    defparam i54209_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52720_3_lut (.I0(n70819), .I1(baudrate[15]), .I2(n37_adj_5026), 
            .I3(GND_net), .O(n69810));   // verilog/uart_rx.v(119[33:55])
    defparam i52720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i44760_1_lut (.I0(n25376), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61800));
    defparam i44760_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5290), .I1(baudrate[9]), 
            .I2(n25_adj_5050), .I3(GND_net), .O(n22_adj_5291));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54207_4_lut (.I0(n22_adj_5291), .I1(n12_adj_5292), .I2(n25_adj_5050), 
            .I3(n69207), .O(n71297));   // verilog/uart_rx.v(119[33:55])
    defparam i54207_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54208_3_lut (.I0(n71297), .I1(baudrate[10]), .I2(n27_adj_5051), 
            .I3(GND_net), .O(n71298));   // verilog/uart_rx.v(119[33:55])
    defparam i54208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54043_3_lut (.I0(n71298), .I1(baudrate[11]), .I2(n29_adj_5047), 
            .I3(GND_net), .O(n71133));   // verilog/uart_rx.v(119[33:55])
    defparam i54043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53906_4_lut (.I0(n39_adj_5052), .I1(n37_adj_5026), .I2(n35_adj_5027), 
            .I3(n69197), .O(n70996));
    defparam i53906_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54414_4_lut (.I0(n69810), .I1(n71299), .I2(n41), .I3(n69186), 
            .O(n71504));   // verilog/uart_rx.v(119[33:55])
    defparam i54414_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52718_3_lut (.I0(n71133), .I1(baudrate[12]), .I2(n31_adj_5048), 
            .I3(GND_net), .O(n69808));   // verilog/uart_rx.v(119[33:55])
    defparam i52718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48151_1_lut (.I0(n65231), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61837));
    defparam i48151_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54468_4_lut (.I0(n69808), .I1(n71504), .I2(n41), .I3(n70996), 
            .O(n71558));   // verilog/uart_rx.v(119[33:55])
    defparam i54468_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54469_3_lut (.I0(n71558), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n71559));   // verilog/uart_rx.v(119[33:55])
    defparam i54469_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54465_3_lut (.I0(n71559), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n71555));   // verilog/uart_rx.v(119[33:55])
    defparam i54465_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8235[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8261[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8287[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1058 (.I0(n64627), .I1(n64629), .I2(n64485), 
            .I3(n64625), .O(n25379));
    defparam i1_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8287[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8287[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8287[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8287[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8287[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8287[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8287[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8287[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8287[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8287[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8287[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8287[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8287[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8287[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8287[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8287[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8287[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8287[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8287[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8287[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8261[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8261[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8261[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8261[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8261[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8261[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n64629));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5292));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52117_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n69207));
    defparam i52117_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5290));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5289));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52092_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n69182));
    defparam i52092_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5287));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54645_2_lut_4_lut (.I0(n71501), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25411), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i54645_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51483_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n68573));
    defparam i51483_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_adj_1059 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64131), .I3(GND_net), .O(n64079));
    defparam i1_2_lut_3_lut_adj_1059.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1060 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64167), .I3(GND_net), .O(n64205));
    defparam i1_2_lut_3_lut_adj_1060.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1061 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64167), .I3(GND_net), .O(n64169));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1061.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1062 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64131), .I3(GND_net), .O(n64151));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1062.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_4_lut_adj_1063 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n64543));
    defparam i1_2_lut_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1064 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n64545));
    defparam i1_2_lut_4_lut_adj_1064.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5293));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5224), 
            .O(n15_adj_5294));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5294), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5293), 
            .I3(n60695), .O(n72443));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51529_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n68619));
    defparam i51529_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54661_2_lut_4_lut (.I0(n71342), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25379), .O(n294[1]));
    defparam i54661_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_3_lut_adj_1065 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64131), .I3(GND_net), .O(n64133));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1065.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1066 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n64167), .I3(GND_net), .O(n64097));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1066.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54639_2_lut_4_lut (.I0(n71101), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25437), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i54639_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51966_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n69056));
    defparam i51966_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51996_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n69086));
    defparam i51996_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1067 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n64505));
    defparam i1_2_lut_4_lut_adj_1067.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52356_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n69446));
    defparam i52356_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63701), .I3(n48_adj_5152), .O(n32_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54633_2_lut_4_lut (.I0(n71115), .I1(baudrate[5]), .I2(n61512), 
            .I3(n25353), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i54633_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i52363_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n69453));
    defparam i52363_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut (.I0(n25388), .I1(n48_adj_5175), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5198));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i54498_2_lut_4_lut (.I0(n71117), .I1(baudrate[4]), .I2(n61510), 
            .I3(n65267), .O(n294[19]));
    defparam i54498_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i47945_1_lut_2_lut (.I0(baudrate[17]), .I1(n25423), .I2(GND_net), 
            .I3(GND_net), .O(n61820));
    defparam i47945_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i4031_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam i4031_2_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i5971_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21488));   // verilog/uart_rx.v(119[33:55])
    defparam i5971_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52283_2_lut_3_lut (.I0(n25388), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n68374));   // verilog/uart_rx.v(119[33:55])
    defparam i52283_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i51418_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n68508));
    defparam i51418_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54729_2_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n27511));
    defparam i54729_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63707), .I3(n48_adj_5134), .O(n18_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i51424_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n68514));
    defparam i51424_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 equal_349_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(98[17:39])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51628_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5175), .I2(n25388), 
            .I3(GND_net), .O(n68718));   // verilog/uart_rx.v(119[33:55])
    defparam i51628_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i51448_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n68538));
    defparam i51448_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51452_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n68542));
    defparam i51452_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1068 (.I0(n71555), .I1(baudrate[20]), .I2(n2938), 
            .I3(n63717), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1068.LUT_INIT = 16'h7100;
    SB_LUT4 i54636_2_lut_4_lut (.I0(n71555), .I1(baudrate[20]), .I2(n2938), 
            .I3(n65263), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i54636_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1069 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n63625));
    defparam i1_3_lut_4_lut_adj_1069.LUT_INIT = 16'hfffe;
    SB_LUT4 i48037_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n65116));
    defparam i48037_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48041_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n65120));
    defparam i48041_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1070 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n64409));
    defparam i1_2_lut_4_lut_adj_1070.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_4_lut_adj_1071 (.I0(n64267), .I1(n65022), .I2(n8053[11]), 
            .I3(n48_adj_5277), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1071.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_4_lut_adj_1072 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n64475));
    defparam i1_2_lut_4_lut_adj_1072.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1073 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n64473));
    defparam i1_2_lut_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i54630_2_lut_4_lut (.I0(n46_adj_5193), .I1(baudrate[3]), .I2(n61508), 
            .I3(n25391), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i54630_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i1_2_lut_4_lut_adj_1074 (.I0(n71441), .I1(baudrate[17]), .I2(n2596), 
            .I3(n63711), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1074.LUT_INIT = 16'h7100;
    SB_LUT4 i54568_2_lut_4_lut (.I0(n71441), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25423), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i54568_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i51583_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n68673));   // verilog/uart_rx.v(119[33:55])
    defparam i51583_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_3_lut_4_lut_adj_1075 (.I0(n64463), .I1(n65231), .I2(n7975[14]), 
            .I3(n48_adj_5226), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1075.LUT_INIT = 16'h0010;
    SB_LUT4 i48178_2_lut_3_lut_4_lut (.I0(n64463), .I1(n65231), .I2(baudrate[8]), 
            .I3(baudrate[9]), .O(n65259));
    defparam i48178_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54525_2_lut_3_lut_4_lut (.I0(n64463), .I1(n65231), .I2(n48_adj_5152), 
            .I3(baudrate[9]), .O(n294[15]));
    defparam i54525_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i51606_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n68696));   // verilog/uart_rx.v(119[33:55])
    defparam i51606_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i4202_2_lut_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam i4202_2_lut_4_lut.LUT_INIT = 16'hb2bb;
    SB_LUT4 i51619_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n68709));   // verilog/uart_rx.v(119[33:55])
    defparam i51619_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51651_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n68741));   // verilog/uart_rx.v(119[33:55])
    defparam i51651_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i4200_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9783));   // verilog/uart_rx.v(119[33:55])
    defparam i4200_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i1_2_lut_4_lut_adj_1076 (.I0(n71351), .I1(baudrate[16]), .I2(n2476), 
            .I3(n63709), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1076.LUT_INIT = 16'h7100;
    SB_LUT4 i54564_2_lut_4_lut (.I0(n71351), .I1(baudrate[16]), .I2(n2476), 
            .I3(n65018), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i54564_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_3_lut_4_lut_adj_1077 (.I0(baudrate[2]), .I1(n42_adj_5172), 
            .I2(baudrate[3]), .I3(n21490), .O(n62307));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1077.LUT_INIT = 16'hff4f;
    SB_LUT4 i4038_2_lut_3_lut (.I0(baudrate[2]), .I1(n42_adj_5172), .I2(n21490), 
            .I3(GND_net), .O(n44_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam i4038_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 i1_2_lut_4_lut_adj_1078 (.I0(n71063), .I1(baudrate[21]), .I2(n3046), 
            .I3(n63719), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1078.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_866_i36_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n63697), .I3(n48_adj_5206), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i54658_2_lut_4_lut (.I0(n71063), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25376), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i54658_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51547_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n68637));
    defparam i51547_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_adj_1079 (.I0(baudrate[30]), .I1(baudrate[31]), 
            .I2(baudrate[27]), .I3(baudrate[24]), .O(n63623));
    defparam i1_3_lut_4_lut_adj_1079.LUT_INIT = 16'hfffe;
    SB_LUT4 i48138_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n65219));
    defparam i48138_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48181_1_lut_2_lut (.I0(baudrate[7]), .I1(n65259), .I2(GND_net), 
            .I3(GND_net), .O(n61854));
    defparam i48181_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i54501_2_lut_3_lut (.I0(baudrate[7]), .I1(n65259), .I2(n48_adj_5206), 
            .I3(GND_net), .O(n294[17]));
    defparam i54501_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_4_lut_adj_1080 (.I0(n60415), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n63821));
    defparam i1_3_lut_4_lut_adj_1080.LUT_INIT = 16'hfdfc;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51466_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n68556));
    defparam i51466_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51472_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n68562));
    defparam i51472_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47949_1_lut (.I0(n65022), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n61828));
    defparam i47949_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52305_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n69395));
    defparam i52305_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52273_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n69363));
    defparam i52273_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1081 (.I0(baudrate[3]), .I1(n42_adj_5167), 
            .I2(baudrate[4]), .I3(n21504), .O(n62259));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1081.LUT_INIT = 16'hff4f;
    SB_LUT4 i4209_2_lut_3_lut (.I0(baudrate[3]), .I1(n42_adj_5167), .I2(n21504), 
            .I3(GND_net), .O(n44_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam i4209_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54515_2_lut_4_lut (.I0(n71294), .I1(baudrate[7]), .I2(n1261), 
            .I3(n65259), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i54515_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1082 (.I0(n71294), .I1(baudrate[7]), .I2(n1261), 
            .I3(n63699), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1082.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51639_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n68729));   // verilog/uart_rx.v(119[33:55])
    defparam i51639_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1083 (.I0(n71395), .I1(baudrate[11]), .I2(n1831), 
            .I3(n63703), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1083.LUT_INIT = 16'h7100;
    SB_LUT4 i54539_2_lut_4_lut (.I0(n71395), .I1(baudrate[11]), .I2(n1831), 
            .I3(n65231), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i54539_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52239_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n69329));
    defparam i52239_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1084 (.I0(n71340), .I1(baudrate[14]), .I2(n2227), 
            .I3(n63705), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1084.LUT_INIT = 16'h7100;
    SB_LUT4 i54555_2_lut_4_lut (.I0(n71340), .I1(baudrate[14]), .I2(n2227), 
            .I3(n65022), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i54555_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52181_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n69271));
    defparam i52181_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1085 (.I0(n71355), .I1(baudrate[18]), .I2(n2713), 
            .I3(n63713), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1085.LUT_INIT = 16'h7100;
    SB_LUT4 i54572_2_lut_4_lut (.I0(n71355), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25426), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i54572_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52019_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n69109));
    defparam i52019_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52051_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n69141));
    defparam i52051_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1792, ENCODER1_A_N_keep, 
            \encoder1_position[31] , GND_net, \encoder1_position[30] , 
            \encoder1_position[29] , \encoder1_position[28] , \encoder1_position[27] , 
            \encoder1_position[26] , \encoder1_position[25] , \encoder1_position[24] , 
            \encoder1_position[23] , \encoder1_position[22] , \encoder1_position[21] , 
            \encoder1_position[20] , \encoder1_position[19] , \encoder1_position[18] , 
            \encoder1_position[17] , \encoder1_position[16] , \encoder1_position[15] , 
            \encoder1_position[14] , \encoder1_position[13] , \encoder1_position[12] , 
            \encoder1_position[11] , \encoder1_position[10] , \encoder1_position[9] , 
            \encoder1_position[8] , \encoder1_position[7] , \encoder1_position[6] , 
            \encoder1_position[5] , \encoder1_position[4] , \encoder1_position[3] , 
            \encoder1_position[2] , n1829, n1831, VCC_net, b_prev, 
            \a_new[1] , \b_new[1] , n29239, a_prev, position_31__N_3836, 
            n29125, n29124, n1797, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1792;
    input ENCODER1_A_N_keep;
    output \encoder1_position[31] ;
    input GND_net;
    output \encoder1_position[30] ;
    output \encoder1_position[29] ;
    output \encoder1_position[28] ;
    output \encoder1_position[27] ;
    output \encoder1_position[26] ;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output n1829;
    output n1831;
    input VCC_net;
    output b_prev;
    output \a_new[1] ;
    output \b_new[1] ;
    input n29239;
    output a_prev;
    output position_31__N_3836;
    input n29125;
    input n29124;
    output n1797;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n54514, n54513, n54512, n54511, n54510, 
        n54509, n54508, n54507, n54506, n54505, n54504, n54503, 
        n54502, n54501, n54500, n54499, n54498, n54497, n54496, 
        n54495, n54494, n54493, n54492, n54491, n54490, n54489, 
        n54488, n54487, n54486, n54485, n54484;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1792), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1792), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2041_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[31] ), .I3(n54514), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2041_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[30] ), .I3(n54513), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_32 (.CI(n54513), .I0(direction_N_3840), 
            .I1(\encoder1_position[30] ), .CO(n54514));
    SB_LUT4 position_2041_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[29] ), .I3(n54512), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_31 (.CI(n54512), .I0(direction_N_3840), 
            .I1(\encoder1_position[29] ), .CO(n54513));
    SB_LUT4 position_2041_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[28] ), .I3(n54511), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_30 (.CI(n54511), .I0(direction_N_3840), 
            .I1(\encoder1_position[28] ), .CO(n54512));
    SB_LUT4 position_2041_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[27] ), .I3(n54510), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_29 (.CI(n54510), .I0(direction_N_3840), 
            .I1(\encoder1_position[27] ), .CO(n54511));
    SB_LUT4 position_2041_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[26] ), .I3(n54509), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_28 (.CI(n54509), .I0(direction_N_3840), 
            .I1(\encoder1_position[26] ), .CO(n54510));
    SB_LUT4 position_2041_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[25] ), .I3(n54508), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_27 (.CI(n54508), .I0(direction_N_3840), 
            .I1(\encoder1_position[25] ), .CO(n54509));
    SB_LUT4 position_2041_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[24] ), .I3(n54507), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_26 (.CI(n54507), .I0(direction_N_3840), 
            .I1(\encoder1_position[24] ), .CO(n54508));
    SB_LUT4 position_2041_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[23] ), .I3(n54506), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_25 (.CI(n54506), .I0(direction_N_3840), 
            .I1(\encoder1_position[23] ), .CO(n54507));
    SB_LUT4 position_2041_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[22] ), .I3(n54505), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_24 (.CI(n54505), .I0(direction_N_3840), 
            .I1(\encoder1_position[22] ), .CO(n54506));
    SB_LUT4 position_2041_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[21] ), .I3(n54504), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_23 (.CI(n54504), .I0(direction_N_3840), 
            .I1(\encoder1_position[21] ), .CO(n54505));
    SB_LUT4 position_2041_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[20] ), .I3(n54503), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_22 (.CI(n54503), .I0(direction_N_3840), 
            .I1(\encoder1_position[20] ), .CO(n54504));
    SB_LUT4 position_2041_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[19] ), .I3(n54502), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_21 (.CI(n54502), .I0(direction_N_3840), 
            .I1(\encoder1_position[19] ), .CO(n54503));
    SB_LUT4 position_2041_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[18] ), .I3(n54501), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_20 (.CI(n54501), .I0(direction_N_3840), 
            .I1(\encoder1_position[18] ), .CO(n54502));
    SB_LUT4 position_2041_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[17] ), .I3(n54500), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_19 (.CI(n54500), .I0(direction_N_3840), 
            .I1(\encoder1_position[17] ), .CO(n54501));
    SB_LUT4 position_2041_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[16] ), .I3(n54499), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_18 (.CI(n54499), .I0(direction_N_3840), 
            .I1(\encoder1_position[16] ), .CO(n54500));
    SB_LUT4 position_2041_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[15] ), .I3(n54498), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_17 (.CI(n54498), .I0(direction_N_3840), 
            .I1(\encoder1_position[15] ), .CO(n54499));
    SB_LUT4 position_2041_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[14] ), .I3(n54497), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_16 (.CI(n54497), .I0(direction_N_3840), 
            .I1(\encoder1_position[14] ), .CO(n54498));
    SB_LUT4 position_2041_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[13] ), .I3(n54496), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_15 (.CI(n54496), .I0(direction_N_3840), 
            .I1(\encoder1_position[13] ), .CO(n54497));
    SB_LUT4 position_2041_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[12] ), .I3(n54495), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_14 (.CI(n54495), .I0(direction_N_3840), 
            .I1(\encoder1_position[12] ), .CO(n54496));
    SB_LUT4 position_2041_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[11] ), .I3(n54494), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_13 (.CI(n54494), .I0(direction_N_3840), 
            .I1(\encoder1_position[11] ), .CO(n54495));
    SB_LUT4 position_2041_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[10] ), .I3(n54493), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_12 (.CI(n54493), .I0(direction_N_3840), 
            .I1(\encoder1_position[10] ), .CO(n54494));
    SB_LUT4 position_2041_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[9] ), .I3(n54492), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_11 (.CI(n54492), .I0(direction_N_3840), 
            .I1(\encoder1_position[9] ), .CO(n54493));
    SB_LUT4 position_2041_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[8] ), .I3(n54491), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_10 (.CI(n54491), .I0(direction_N_3840), 
            .I1(\encoder1_position[8] ), .CO(n54492));
    SB_LUT4 position_2041_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[7] ), .I3(n54490), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_9 (.CI(n54490), .I0(direction_N_3840), 
            .I1(\encoder1_position[7] ), .CO(n54491));
    SB_LUT4 position_2041_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[6] ), .I3(n54489), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_8 (.CI(n54489), .I0(direction_N_3840), 
            .I1(\encoder1_position[6] ), .CO(n54490));
    SB_LUT4 position_2041_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[5] ), .I3(n54488), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_7 (.CI(n54488), .I0(direction_N_3840), 
            .I1(\encoder1_position[5] ), .CO(n54489));
    SB_LUT4 position_2041_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[4] ), .I3(n54487), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_6 (.CI(n54487), .I0(direction_N_3840), 
            .I1(\encoder1_position[4] ), .CO(n54488));
    SB_LUT4 position_2041_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[3] ), .I3(n54486), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_5 (.CI(n54486), .I0(direction_N_3840), 
            .I1(\encoder1_position[3] ), .CO(n54487));
    SB_LUT4 position_2041_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder1_position[2] ), .I3(n54485), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_4 (.CI(n54485), .I0(direction_N_3840), 
            .I1(\encoder1_position[2] ), .CO(n54486));
    SB_LUT4 position_2041_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1829), .I3(n54484), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_3 (.CI(n54484), .I0(direction_N_3840), 
            .I1(n1829), .CO(n54485));
    SB_LUT4 position_2041_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1831), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1831), 
            .CO(n54484));
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1792), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1792), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1792), .D(n29239));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i0 (.Q(n1831), .C(n1792), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1792), .D(n29125));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1797), .C(n1792), .D(n29124));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i1 (.Q(n1829), .C(n1792), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i2 (.Q(\encoder1_position[2] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i3 (.Q(\encoder1_position[3] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i4 (.Q(\encoder1_position[4] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i5 (.Q(\encoder1_position[5] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i6 (.Q(\encoder1_position[6] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i7 (.Q(\encoder1_position[7] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i8 (.Q(\encoder1_position[8] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i9 (.Q(\encoder1_position[9] ), .C(n1792), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i10 (.Q(\encoder1_position[10] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i11 (.Q(\encoder1_position[11] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i12 (.Q(\encoder1_position[12] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i13 (.Q(\encoder1_position[13] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i14 (.Q(\encoder1_position[14] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i15 (.Q(\encoder1_position[15] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i16 (.Q(\encoder1_position[16] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i17 (.Q(\encoder1_position[17] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i18 (.Q(\encoder1_position[18] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i19 (.Q(\encoder1_position[19] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i20 (.Q(\encoder1_position[20] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i21 (.Q(\encoder1_position[21] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i22 (.Q(\encoder1_position[22] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i23 (.Q(\encoder1_position[23] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i24 (.Q(\encoder1_position[24] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i25 (.Q(\encoder1_position[25] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i26 (.Q(\encoder1_position[26] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i27 (.Q(\encoder1_position[27] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i28 (.Q(\encoder1_position[28] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i29 (.Q(\encoder1_position[29] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i30 (.Q(\encoder1_position[30] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i31 (.Q(\encoder1_position[31] ), .C(n1792), 
            .E(position_31__N_3836), .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\data[15] , \state[1] , \state[0] , n27489, GND_net, 
            \data[12] , clk16MHz, n6, n5, n5_adj_8, n6_adj_9, n39133, 
            n39146, \current[15] , n29320, \current[1] , n29319, \current[2] , 
            n29318, \current[3] , n29317, \current[4] , n29316, \current[5] , 
            n29315, \current[6] , n29314, \current[7] , n29313, \current[8] , 
            n29312, \current[9] , n29311, \current[10] , n29310, \current[11] , 
            n15, n11, n29880, n29879, n29878, \data[11] , n29877, 
            \data[10] , n29875, \data[9] , n29874, \data[8] , n29872, 
            \data[7] , n29871, \data[6] , n29869, \data[5] , n29868, 
            \data[4] , n29866, \data[3] , n29865, \data[2] , n29840, 
            \data[1] , n9, clk_out, n29119, CS_c, n29114, \current[0] , 
            n29683, \data[0] , VCC_net, n25298, n25289, state_7__N_4319, 
            CS_CLK_c, n25328, n25345, n25316) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \data[15] ;
    output \state[1] ;
    output \state[0] ;
    output n27489;
    input GND_net;
    output \data[12] ;
    input clk16MHz;
    output n6;
    output n5;
    output n5_adj_8;
    output n6_adj_9;
    output n39133;
    output n39146;
    output \current[15] ;
    input n29320;
    output \current[1] ;
    input n29319;
    output \current[2] ;
    input n29318;
    output \current[3] ;
    input n29317;
    output \current[4] ;
    input n29316;
    output \current[5] ;
    input n29315;
    output \current[6] ;
    input n29314;
    output \current[7] ;
    input n29313;
    output \current[8] ;
    input n29312;
    output \current[9] ;
    input n29311;
    output \current[10] ;
    input n29310;
    output \current[11] ;
    output n15;
    output n11;
    input n29880;
    input n29879;
    input n29878;
    output \data[11] ;
    input n29877;
    output \data[10] ;
    input n29875;
    output \data[9] ;
    input n29874;
    output \data[8] ;
    input n29872;
    output \data[7] ;
    input n29871;
    output \data[6] ;
    input n29869;
    output \data[5] ;
    input n29868;
    output \data[4] ;
    input n29866;
    output \data[3] ;
    input n29865;
    output \data[2] ;
    input n29840;
    output \data[1] ;
    input n9;
    output clk_out;
    input n29119;
    output CS_c;
    input n29114;
    output \current[0] ;
    input n29683;
    output \data[0] ;
    input VCC_net;
    output n25298;
    output n25289;
    output state_7__N_4319;
    output CS_CLK_c;
    output n25328;
    output n25345;
    output n25316;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [13:0]n241;
    
    wire clk_slow_N_4232;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire clk_slow_N_4233;
    wire [7:0]n37;
    
    wire n27625, n29075, n22406;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire delay_counter_15__N_4314;
    wire [2:0]n17;
    
    wire n10011, n39469, n27582, n28549, n6_adj_5022, n22410, n22412, 
        n22414, n63269, n10, n12, n68371, n2, n54578, n54577, 
        n54576, n54575, n54574, n54573, n54572, n54571, n54570, 
        n54569, n54568, n54567, n54566, n54552, n54551, n54550, 
        n54549, n68378, n54548, n68379, n54547, n68387, n54546;
    
    SB_LUT4 i54527_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n27489));
    defparam i54527_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2243_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2243_1_lut.LUT_INIT = 16'h5555;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 equal_337_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_8));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_332_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_9));   // verilog/tli4970.v(54[9:26])
    defparam equal_332_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i23370_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n39133));
    defparam i23370_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23382_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n39146));
    defparam i23382_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2179_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2179_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27489), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_2044__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27625), 
            .D(n37[7]), .R(n29075));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27625), 
            .D(n37[6]), .R(n29075));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27625), 
            .D(n37[5]), .R(n29075));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27625), 
            .D(n37[4]), .R(n29075));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29320));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29319));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29318));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29317));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29316));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29315));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29314));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29313));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29312));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29311));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29310));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27625), 
            .D(n22406));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 mux_2153_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n10011));
    defparam mux_2153_i2_3_lut.LUT_INIT = 16'h3535;
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n27582), .D(n39469), 
            .S(n28549));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n27582), .D(n10011), 
            .R(n28549));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5022));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_5022), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54550_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n39469));
    defparam i54550_2_lut.LUT_INIT = 16'h1111;
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29880));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29879));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29878));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29877));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29875));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29874));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29872));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29871));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29869));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29868));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29866));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29865));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29840));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29119));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27625), 
            .D(n22410));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29114));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27625), 
            .D(n22412));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27625), 
            .D(n22414));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29683));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNSR delay_counter_2048_2049__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 i2_3_lut (.I0(delay_counter[1]), .I1(delay_counter[4]), .I2(delay_counter[3]), 
            .I3(GND_net), .O(n63269));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_983 (.I0(delay_counter[11]), .I1(delay_counter[9]), 
            .I2(delay_counter[8]), .I3(delay_counter[7]), .O(n10));
    defparam i4_4_lut_adj_983.LUT_INIT = 16'h8000;
    SB_LUT4 i2180_4_lut (.I0(delay_counter[0]), .I1(delay_counter[5]), .I2(delay_counter[2]), 
            .I3(n63269), .O(n12));
    defparam i2180_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i5_4_lut (.I0(n12), .I1(n10), .I2(delay_counter[10]), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'hc080;
    SB_LUT4 i6801_3_lut (.I0(\state[0] ), .I1(n68371), .I2(\state[1] ), 
            .I3(GND_net), .O(n22406));   // verilog/tli4970.v(55[24:39])
    defparam i6801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2521_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));
    defparam i2521_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 counter_2050_2051_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n54578), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2050_2051_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n54577), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_3 (.CI(n54577), .I0(GND_net), .I1(counter[1]), 
            .CO(n54578));
    SB_LUT4 counter_2050_2051_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n54577));
    SB_LUT4 delay_counter_2048_2049_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n54576), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2048_2049_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n54575), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_12 (.CI(n54575), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n54576));
    SB_LUT4 delay_counter_2048_2049_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n54574), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_11 (.CI(n54574), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n54575));
    SB_LUT4 delay_counter_2048_2049_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n54573), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_10 (.CI(n54573), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n54574));
    SB_LUT4 delay_counter_2048_2049_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n54572), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_9 (.CI(n54572), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n54573));
    SB_LUT4 delay_counter_2048_2049_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n54571), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_8 (.CI(n54571), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n54572));
    SB_LUT4 delay_counter_2048_2049_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n54570), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_7 (.CI(n54570), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n54571));
    SB_LUT4 delay_counter_2048_2049_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n54569), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_6 (.CI(n54569), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n54570));
    SB_LUT4 delay_counter_2048_2049_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n54568), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_5 (.CI(n54568), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n54569));
    SB_LUT4 delay_counter_2048_2049_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n54567), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_4 (.CI(n54567), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n54568));
    SB_LUT4 delay_counter_2048_2049_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n54566), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_3 (.CI(n54566), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n54567));
    SB_LUT4 delay_counter_2048_2049_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n54566));
    SB_LUT4 bit_counter_2044_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n54552), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2044_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n54551), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_8 (.CI(n54551), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n54552));
    SB_LUT4 bit_counter_2044_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n54550), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_7 (.CI(n54550), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n54551));
    SB_LUT4 bit_counter_2044_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n54549), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_6 (.CI(n54549), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n54550));
    SB_LUT4 bit_counter_2044_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n54548), .O(n68378)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_5 (.CI(n54548), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n54549));
    SB_LUT4 bit_counter_2044_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n54547), .O(n68379)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_4 (.CI(n54547), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n54548));
    SB_LUT4 bit_counter_2044_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n54546), .O(n68387)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_3 (.CI(n54546), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n54547));
    SB_LUT4 bit_counter_2044_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n68371)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n54546));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n25298));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_984 (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n25289));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut_adj_984.LUT_INIT = 16'hfeff;
    SB_LUT4 i13214_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29075));   // verilog/tli4970.v(55[24:39])
    defparam i13214_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i11840_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27625));
    defparam i11840_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i6808_3_lut (.I0(\state[0] ), .I1(n68378), .I2(\state[1] ), 
            .I3(GND_net), .O(n22414));   // verilog/tli4970.v(55[24:39])
    defparam i6808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6806_3_lut (.I0(\state[0] ), .I1(n68379), .I2(\state[1] ), 
            .I3(GND_net), .O(n22412));   // verilog/tli4970.v(55[24:39])
    defparam i6806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6804_3_lut (.I0(\state[0] ), .I1(n68387), .I2(\state[1] ), 
            .I3(GND_net), .O(n22410));   // verilog/tli4970.v(55[24:39])
    defparam i6804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n27582));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i12688_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4314), .O(n28549));
    defparam i12688_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_985 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25328));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_985.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_986 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25345));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_986.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_4_lut_adj_987 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25316));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_987.LUT_INIT = 16'hffbf;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, enable_slow_N_4213, clk16MHz, \state_7__N_4110[0] , 
            ID, baudrate, n29328, n29327, n29326, n29325, n29324, 
            n29323, n29322, n29321, data_ready, \state_7__N_3918[0] , 
            n63193, data, \state[0] , \state_7__N_4126[3] , scl_enable, 
            scl, n6714, sda_enable, n29668, n6, VCC_net, n29663, 
            n29661, n29660, n29659, n29658, n29654, n29652, sda_out, 
            n39034, n10, n25302, n25348, n4, n4_adj_6, n39188, 
            n10_adj_7) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output enable_slow_N_4213;
    input clk16MHz;
    output \state_7__N_4110[0] ;
    output [7:0]ID;
    output [31:0]baudrate;
    input n29328;
    input n29327;
    input n29326;
    input n29325;
    input n29324;
    input n29323;
    input n29322;
    input n29321;
    output data_ready;
    input \state_7__N_3918[0] ;
    output n63193;
    output [7:0]data;
    output \state[0] ;
    input \state_7__N_4126[3] ;
    output scl_enable;
    output scl;
    output n6714;
    output sda_enable;
    input n29668;
    input n6;
    input VCC_net;
    input n29663;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29654;
    input n29652;
    output sda_out;
    output n39034;
    output n10;
    output n25302;
    output n25348;
    output n4;
    output n4_adj_6;
    output n39188;
    output n10_adj_7;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n60736, n25161;
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire n68479, n4_c, n47932, n63215, n39479;
    wire [7:0]state_7__N_3885;
    
    wire n53830;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    wire [15:0]n5400;
    
    wire n53831;
    wire [15:0]delay_counter_15__N_3956;
    
    wire n53829, n28, n26, n27, n25, ready_prev;
    wire [0:0]n5934;
    
    wire enable, n71574, n47917;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n47909, n68478, n27480, enable_slow_N_4212, n6939, n28842, 
        n6941, n6942, n6943, n6944, n6945, n55114, n55756, n27671, 
        n29079, n29369, n29368, n29367, n29366, n29365, n29364, 
        n29363, n29362, n29361, n29360, n29359, n29358, n29357, 
        n29356, n29355, n29354, n29353, n29352, n29351, n29350, 
        n29349, n29348;
    wire [2:0]n17;
    
    wire n29337, n29336, n29335, n29334, n29333, n29332, n29331, 
        n29330, n29329, n60014, rw, n29693, n60106, n29112, n60050, 
        n39283, n53843, n53842, n53841, n53840, n53839, n53838, 
        n53837, n53836, n53835, n53834, n53833, n53832, n65154, 
        n68472, n21372, n4_adj_5013, n60756, n60733, n4_adj_5014, 
        n6_c, n12;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n60304;
    
    SB_LUT4 i51869_3_lut (.I0(n60736), .I1(n25161), .I2(state[1]), .I3(GND_net), 
            .O(n68479));
    defparam i51869_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_4_lut (.I0(n68479), .I1(n4_c), .I2(n47932), .I3(state[0]), 
            .O(n63215));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i6838_4_lut (.I0(state[1]), .I1(n39479), .I2(state[2]), .I3(state[0]), 
            .O(state_7__N_3885[1]));   // verilog/eeprom.v(38[3] 80[10])
    defparam i6838_4_lut.LUT_INIT = 16'ha5ba;
    SB_CARRY add_1198_4 (.CI(n53830), .I0(delay_counter[2]), .I1(n5400[9]), 
            .CO(n53831));
    SB_LUT4 add_1198_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5400[9]), 
            .I3(n53829), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_3 (.CI(n53829), .I0(delay_counter[1]), .I1(n5400[9]), 
            .CO(n53830));
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n25161));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i54565_2_lut (.I0(n25161), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5400[9]));
    defparam i54565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_1198_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5400[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5400[9]), 
            .CO(n53829));
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5934[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i54484_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n71574));   // verilog/eeprom.v(27[11:16])
    defparam i54484_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n47917));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23711_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n39479));
    defparam i23711_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut (.I0(n47909), .I1(n71574), .I2(n68478), .I3(state[2]), 
            .O(n27480));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut.LUT_INIT = 16'hafee;
    SB_LUT4 i54512_2_lut (.I0(\state_7__N_4110[0] ), .I1(enable_slow_N_4213), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));
    defparam i54512_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27480), 
            .D(delay_counter_15__N_3956[1]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27480), 
            .D(delay_counter_15__N_3956[2]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27480), 
            .D(delay_counter_15__N_3956[3]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27480), 
            .D(n6939), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27480), 
            .D(delay_counter_15__N_3956[5]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27480), 
            .D(n6941), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27480), 
            .D(n6942), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27480), 
            .D(n6943), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27480), 
            .D(n6944), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27480), .D(n6945), .S(n28842));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27480), .D(delay_counter_15__N_3956[11]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27480), .D(delay_counter_15__N_3956[12]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27480), .D(delay_counter_15__N_3956[13]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27480), .D(delay_counter_15__N_3956[14]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27480), .D(delay_counter_15__N_3956[15]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i2_3_lut (.I0(state[0]), .I1(n25161), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n55114));
    defparam i2_3_lut.LUT_INIT = 16'hefef;
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n63215), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27671), .D(n55756), .R(n29079));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n29369));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n29368));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n29367));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n29366));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n29365));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n29364));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n29363));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n29362));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n29361));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n29360));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n29359));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n29358));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n29357));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n29356));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n29355));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n29354));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n29353));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n29352));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n29351));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n29350));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n29349));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n29348));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27671), .D(n17[2]), .R(n29079));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27671), .D(n17[1]), .R(n29079));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n29337));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n29336));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n29335));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n29334));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n29333));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n29332));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n29331));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n29330));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n29329));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n29328));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n29327));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n29326));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n29325));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n29324));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n29323));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n29322));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n29321));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27480), 
            .D(delay_counter_15__N_3956[0]), .R(n47909));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_4_lut_4_lut (.I0(state[0]), .I1(n39479), .I2(state[2]), 
            .I3(state[1]), .O(n47909));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i12985_2_lut_4_lut (.I0(state[0]), .I1(n39479), .I2(state[2]), 
            .I3(n27480), .O(n28842));
    defparam i12985_2_lut_4_lut.LUT_INIT = 16'h3a00;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n60014));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n29693));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n60106));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29112));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n60050));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i23519_2_lut (.I0(state[2]), .I1(n39479), .I2(GND_net), .I3(GND_net), 
            .O(n39283));
    defparam i23519_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 add_1198_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5400[9]), 
            .I3(n53843), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1198_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5400[9]), 
            .I3(n53842), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_16 (.CI(n53842), .I0(delay_counter[14]), .I1(n5400[9]), 
            .CO(n53843));
    SB_LUT4 add_1198_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5400[9]), 
            .I3(n53841), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_15 (.CI(n53841), .I0(delay_counter[13]), .I1(n5400[9]), 
            .CO(n53842));
    SB_LUT4 add_1198_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5400[9]), 
            .I3(n53840), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_14 (.CI(n53840), .I0(delay_counter[12]), .I1(n5400[9]), 
            .CO(n53841));
    SB_LUT4 add_1198_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5400[9]), 
            .I3(n53839), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_13 (.CI(n53839), .I0(delay_counter[11]), .I1(n5400[9]), 
            .CO(n53840));
    SB_LUT4 add_1198_12_lut (.I0(n39283), .I1(delay_counter[10]), .I2(n5400[9]), 
            .I3(n53838), .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_12 (.CI(n53838), .I0(delay_counter[10]), .I1(n5400[9]), 
            .CO(n53839));
    SB_LUT4 add_1198_11_lut (.I0(n39283), .I1(delay_counter[9]), .I2(n5400[9]), 
            .I3(n53837), .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_11 (.CI(n53837), .I0(delay_counter[9]), .I1(n5400[9]), 
            .CO(n53838));
    SB_LUT4 add_1198_10_lut (.I0(n39283), .I1(delay_counter[8]), .I2(n5400[9]), 
            .I3(n53836), .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_10 (.CI(n53836), .I0(delay_counter[8]), .I1(n5400[9]), 
            .CO(n53837));
    SB_LUT4 add_1198_9_lut (.I0(n39283), .I1(delay_counter[7]), .I2(n5400[9]), 
            .I3(n53835), .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_9 (.CI(n53835), .I0(delay_counter[7]), .I1(n5400[9]), 
            .CO(n53836));
    SB_LUT4 add_1198_8_lut (.I0(n39283), .I1(delay_counter[6]), .I2(n5400[9]), 
            .I3(n53834), .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_8 (.CI(n53834), .I0(delay_counter[6]), .I1(n5400[9]), 
            .CO(n53835));
    SB_LUT4 add_1198_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5400[9]), 
            .I3(n53833), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_7 (.CI(n53833), .I0(delay_counter[5]), .I1(n5400[9]), 
            .CO(n53834));
    SB_LUT4 add_1198_6_lut (.I0(n39283), .I1(delay_counter[4]), .I2(n5400[9]), 
            .I3(n53832), .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_6 (.CI(n53832), .I0(delay_counter[4]), .I1(n5400[9]), 
            .CO(n53833));
    SB_LUT4 i1_2_lut_3_lut (.I0(ready_prev), .I1(enable_slow_N_4213), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n55756));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hb4b4;
    SB_LUT4 i1_4_lut_4_lut_adj_975 (.I0(state[2]), .I1(state[1]), .I2(state[0]), 
            .I3(\state_7__N_3918[0] ), .O(n27671));
    defparam i1_4_lut_4_lut_adj_975.LUT_INIT = 16'h4140;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state_7__N_3918[0] ), .I1(state[0]), .I2(state[1]), 
            .I3(state[2]), .O(n29079));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i11_4_lut_4_lut (.I0(rw), .I1(state[1]), .I2(state[0]), .I3(n65154), 
            .O(n60014));   // verilog/eeprom.v(27[11:16])
    defparam i11_4_lut_4_lut.LUT_INIT = 16'haace;
    SB_LUT4 i1_4_lut_adj_976 (.I0(state[2]), .I1(state[1]), .I2(\state_7__N_3918[0] ), 
            .I3(state[0]), .O(n4_c));
    defparam i1_4_lut_adj_976.LUT_INIT = 16'hbbba;
    SB_LUT4 i52329_2_lut_3_lut (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(state[1]), .I3(GND_net), .O(n68472));
    defparam i52329_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 add_1198_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5400[9]), 
            .I3(n53831), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_5 (.CI(n53831), .I0(delay_counter[3]), .I1(n5400[9]), 
            .CO(n53832));
    SB_LUT4 i37661_2_lut_3_lut_4_lut (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i37661_2_lut_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 add_1198_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5400[9]), 
            .I3(n53830), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_977 (.I0(byte_counter[1]), .I1(byte_counter[0]), 
            .I2(n21372), .I3(byte_counter[2]), .O(n63193));   // verilog/eeprom.v(35[8] 81[4])
    defparam i2_3_lut_4_lut_adj_977.LUT_INIT = 16'hfeff;
    SB_LUT4 i13251_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[0]), 
            .I3(ID[0]), .O(n29112));
    defparam i13251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13502_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[7]), 
            .I3(ID[7]), .O(n29363));
    defparam i13502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13503_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[6]), 
            .I3(ID[6]), .O(n29364));
    defparam i13503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13504_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[5]), 
            .I3(ID[5]), .O(n29365));
    defparam i13504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13505_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[4]), 
            .I3(ID[4]), .O(n29366));
    defparam i13505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13506_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[3]), 
            .I3(ID[3]), .O(n29367));
    defparam i13506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13507_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[2]), 
            .I3(ID[2]), .O(n29368));
    defparam i13507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13508_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60756), .I2(data[1]), 
            .I3(ID[1]), .O(n29369));
    defparam i13508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13494_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[7]), 
            .I3(baudrate[7]), .O(n29355));
    defparam i13494_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13495_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[6]), 
            .I3(baudrate[6]), .O(n29356));
    defparam i13495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13496_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[5]), 
            .I3(baudrate[5]), .O(n29357));
    defparam i13496_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13497_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[4]), 
            .I3(baudrate[4]), .O(n29358));
    defparam i13497_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13498_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[3]), 
            .I3(baudrate[3]), .O(n29359));
    defparam i13498_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13499_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[2]), 
            .I3(baudrate[2]), .O(n29360));
    defparam i13499_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13500_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[1]), 
            .I3(baudrate[1]), .O(n29361));
    defparam i13500_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13501_3_lut_4_lut (.I0(n4_adj_5013), .I1(n60733), .I2(data[0]), 
            .I3(baudrate[0]), .O(n29362));
    defparam i13501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13476_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[7]), 
            .I3(baudrate[15]), .O(n29337));
    defparam i13476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13487_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[6]), 
            .I3(baudrate[14]), .O(n29348));
    defparam i13487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13488_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[5]), 
            .I3(baudrate[13]), .O(n29349));
    defparam i13488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13489_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[4]), 
            .I3(baudrate[12]), .O(n29350));
    defparam i13489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13490_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[3]), 
            .I3(baudrate[11]), .O(n29351));
    defparam i13490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13491_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[2]), 
            .I3(baudrate[10]), .O(n29352));
    defparam i13491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13492_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[1]), 
            .I3(baudrate[9]), .O(n29353));
    defparam i13492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13493_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60756), .I2(data[0]), 
            .I3(baudrate[8]), .O(n29354));
    defparam i13493_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_323_i4_2_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5014));   // verilog/eeprom.v(66[9:28])
    defparam equal_323_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_978 (.I0(n21372), .I1(byte_counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n60733));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_979 (.I0(state[2]), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n6_c));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(state[0]), .I1(n60736), .I2(state[1]), .I3(n6_c), 
            .O(n21372));
    defparam i4_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_adj_980 (.I0(byte_counter[0]), .I1(n21372), .I2(GND_net), 
            .I3(GND_net), .O(n60756));
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_LUT4 equal_325_i4_2_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5013));   // verilog/eeprom.v(66[9:28])
    defparam equal_325_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i37668_3_lut_4_lut (.I0(n47932), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i37668_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i13468_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[7]), 
            .I3(baudrate[23]), .O(n29329));
    defparam i13468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13469_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[6]), 
            .I3(baudrate[22]), .O(n29330));
    defparam i13469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13470_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[5]), 
            .I3(baudrate[21]), .O(n29331));
    defparam i13470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13471_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[4]), 
            .I3(baudrate[20]), .O(n29332));
    defparam i13471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13472_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[3]), 
            .I3(baudrate[19]), .O(n29333));
    defparam i13472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13473_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[2]), 
            .I3(baudrate[18]), .O(n29334));
    defparam i13473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13474_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[1]), 
            .I3(baudrate[17]), .O(n29335));
    defparam i13474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13475_3_lut_4_lut (.I0(n4_adj_5014), .I1(n60733), .I2(data[0]), 
            .I3(baudrate[16]), .O(n29336));
    defparam i13475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30_4_lut (.I0(\state_7__N_3918[0] ), .I1(n25161), .I2(state[1]), 
            .I3(n60736), .O(n12));
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12), .I1(n68472), .I2(state[0]), .I3(state[2]), 
            .O(n60050));
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i13_4_lut (.I0(data_ready), .I1(state[2]), .I2(n47917), .I3(n39479), 
            .O(n60106));   // verilog/eeprom.v(27[11:16])
    defparam i13_4_lut.LUT_INIT = 16'haca8;
    SB_LUT4 i1_4_lut_adj_981 (.I0(state[1]), .I1(state[0]), .I2(n47932), 
            .I3(state[2]), .O(n29693));
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hee08;
    SB_LUT4 i48075_3_lut (.I0(state[2]), .I1(n55114), .I2(state[1]), .I3(GND_net), 
            .O(n65154));
    defparam i48075_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i20224_3_lut_4_lut (.I0(state[0]), .I1(n25161), .I2(enable_slow_N_4213), 
            .I3(state[1]), .O(n5934[0]));   // verilog/eeprom.v(27[11:16])
    defparam i20224_3_lut_4_lut.LUT_INIT = 16'h10aa;
    SB_LUT4 i52349_2_lut_3_lut (.I0(n39479), .I1(state[0]), .I2(state[1]), 
            .I3(GND_net), .O(n68478));   // verilog/eeprom.v(27[11:16])
    defparam i52349_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_982 (.I0(rw), .I1(saved_addr[0]), .I2(n60736), 
            .I3(\state_7__N_4110[0] ), .O(n60304));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_982.LUT_INIT = 16'hcacc;
    i2c_controller i2c (.\state[0] (\state[0] ), .\state_7__N_4126[3] (\state_7__N_4126[3] ), 
            .clk16MHz(clk16MHz), .scl_enable(scl_enable), .enable_slow_N_4212(enable_slow_N_4212), 
            .\state_7__N_4110[0] (\state_7__N_4110[0] ), .GND_net(GND_net), 
            .scl(scl), .n6714(n6714), .ready_prev(ready_prev), .enable_slow_N_4213(enable_slow_N_4213), 
            .n47932(n47932), .sda_enable(sda_enable), .\saved_addr[0] (saved_addr[0]), 
            .n60304(n60304), .n29668(n29668), .data({data}), .n6(n6), 
            .VCC_net(VCC_net), .n29663(n29663), .n29661(n29661), .n29660(n29660), 
            .n29659(n29659), .n29658(n29658), .n29654(n29654), .n29652(n29652), 
            .sda_out(sda_out), .n39034(n39034), .n10(n10), .n25302(n25302), 
            .n25348(n25348), .n4(n4), .n4_adj_4(n4_adj_6), .n39188(n39188), 
            .n60736(n60736), .enable(enable), .n10_adj_5(n10_adj_7)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state[0] , \state_7__N_4126[3] , clk16MHz, scl_enable, 
            enable_slow_N_4212, \state_7__N_4110[0] , GND_net, scl, 
            n6714, ready_prev, enable_slow_N_4213, n47932, sda_enable, 
            \saved_addr[0] , n60304, n29668, data, n6, VCC_net, 
            n29663, n29661, n29660, n29659, n29658, n29654, n29652, 
            sda_out, n39034, n10, n25302, n25348, n4, n4_adj_4, 
            n39188, n60736, enable, n10_adj_5) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[0] ;
    input \state_7__N_4126[3] ;
    input clk16MHz;
    output scl_enable;
    input enable_slow_N_4212;
    output \state_7__N_4110[0] ;
    input GND_net;
    output scl;
    output n6714;
    input ready_prev;
    output enable_slow_N_4213;
    output n47932;
    output sda_enable;
    output \saved_addr[0] ;
    input n60304;
    input n29668;
    output [7:0]data;
    input n6;
    input VCC_net;
    input n29663;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29654;
    input n29652;
    output sda_out;
    output n39034;
    output n10;
    output n25302;
    output n25348;
    output n4;
    output n4_adj_4;
    output n39188;
    output n60736;
    input enable;
    output n10_adj_5;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n61685, n15, i2c_clk_N_4199, scl_enable_N_4200, n27553;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n10_c, n28834;
    wire [5:0]n29;
    
    wire n5, n39496, n39323, n39494, n63485, n62660;
    wire [7:0]n119;
    
    wire n27612;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n28819, n62901, n27533, n60064, n62540, n27531, sda_out_adj_5004, 
        n28, n71578, n11, n61579;
    wire [1:0]n6783;
    
    wire n53850, n53849, n53848, n53847, n53846, n53845, n53844, 
        n54629, n54628, n54627, n54626, n54625, n11_adj_5005, n39032, 
        n11_adj_5006, state_7__N_4109, n11_adj_5007, n4_c, n9, n68477, 
        n6707, n63401, n11_adj_5012;
    
    SB_LUT4 i44646_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state_7__N_4126[3] ), 
            .I3(state[2]), .O(n61685));   // verilog/i2c_controller.v(77[27:43])
    defparam i44646_3_lut_4_lut.LUT_INIT = 16'hffd0;
    SB_LUT4 equal_276_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[3]), .I3(state[2]), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_276_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n27553), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n28834));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n28834), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4199));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23333_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i23333_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFSR counter2_2057_2058__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n6714), .D(n5), 
            .S(n39496));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(state[2]), .C(i2c_clk), .E(n6714), .D(n39323), 
            .S(n39494));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(state[3]), .C(i2c_clk), .E(n6714), .D(n63485), 
            .S(n62660));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27612), .D(n119[1]), 
            .S(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27612), .D(n119[2]), 
            .S(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27612), .D(n119[3]), 
            .R(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27612), .D(n119[4]), 
            .R(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27612), .D(n119[5]), 
            .R(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27612), .D(n119[6]), 
            .R(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_961 (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(GND_net), .I3(GND_net), .O(n47932));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i1_2_lut_adj_961.LUT_INIT = 16'hbbbb;
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27612), .D(n119[7]), 
            .R(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27533), 
            .D(n62901), .S(n60064));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_5004), .C(i2c_clk), .E(n27531), 
            .D(n62540), .S(n60064));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27612), .D(n119[0]), 
            .S(n28819));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_4_lut (.I0(state[3]), .I1(state[1]), .I2(\state[0] ), .I3(state[2]), 
            .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i54488_2_lut (.I0(state[3]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n71578));
    defparam i54488_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_962 (.I0(n11), .I1(n71578), .I2(n28), .I3(n61579), 
            .O(n27531));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1830_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6783[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1830_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i44541_2_lut (.I0(state[2]), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n61579));
    defparam i44541_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n11), .I1(n61579), .I2(state[3]), .I3(state[1]), 
            .O(n60064));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_963 (.I0(n11), .I1(state[1]), .I2(state[3]), 
            .I3(n61579), .O(n27533));
    defparam i1_4_lut_adj_963.LUT_INIT = 16'h0a22;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n60304));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29668));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n6));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29663));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29661));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29660));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29659));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29658));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29654));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29652));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n28834));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i2555_2_lut (.I0(sda_out_adj_5004), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n53850), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n53849), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n53849), .I0(counter[6]), .I1(VCC_net), 
            .CO(n53850));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n53848), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n53848), .I0(counter[5]), .I1(VCC_net), 
            .CO(n53849));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n53847), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n53847), .I0(counter[4]), .I1(VCC_net), 
            .CO(n53848));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n53846), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n53846), .I0(counter[3]), .I1(VCC_net), 
            .CO(n53847));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n53845), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n53845), .I0(counter[2]), .I1(VCC_net), 
            .CO(n53846));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n53844), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n53844), .I0(counter[1]), .I1(VCC_net), 
            .CO(n53845));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n53844));
    SB_LUT4 counter2_2057_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n54629), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2057_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n54628), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_6 (.CI(n54628), .I0(GND_net), .I1(counter2[4]), 
            .CO(n54629));
    SB_LUT4 counter2_2057_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n54627), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_5 (.CI(n54627), .I0(GND_net), .I1(counter2[3]), 
            .CO(n54628));
    SB_LUT4 counter2_2057_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n54626), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_4 (.CI(n54626), .I0(GND_net), .I1(counter2[2]), 
            .CO(n54627));
    SB_LUT4 counter2_2057_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n54625), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_3 (.CI(n54625), .I0(GND_net), .I1(counter2[1]), 
            .CO(n54626));
    SB_LUT4 counter2_2057_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n54625));
    SB_LUT4 i23271_2_lut_4_lut (.I0(state[2]), .I1(state[3]), .I2(\state[0] ), 
            .I3(state[1]), .O(n39034));
    defparam i23271_2_lut_4_lut.LUT_INIT = 16'hfebf;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[3]), 
            .I2(\state[0] ), .I3(state[1]), .O(n11_adj_5005));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i23675_2_lut_3_lut (.I0(state[3]), .I1(state[2]), .I2(\state[0] ), 
            .I3(GND_net), .O(n39032));
    defparam i23675_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i23692_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(state[2]), 
            .I3(state[3]), .O(scl_enable_N_4200));   // verilog/i2c_controller.v(44[32:47])
    defparam i23692_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i54651_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(state[1]), 
            .I3(n6714), .O(n62660));
    defparam i54651_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(state[3]), .I3(state[2]), .O(n11_adj_5006));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i23671_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), .I2(state[2]), 
            .I3(state[3]), .O(state_7__N_4109));
    defparam i23671_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(state[3]), .I1(state[2]), 
            .I2(state[1]), .I3(\state[0] ), .O(n11_adj_5007));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(n4_c), .I3(n9), 
            .O(n63485));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hf0f2;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n25302));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_964 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n25348));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_964.LUT_INIT = 16'hfefe;
    SB_LUT4 i54653_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_5007), 
            .I3(n6714), .O(n39494));   // verilog/i2c_controller.v(151[5:14])
    defparam i54653_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 equal_1562_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(state[3]), .I3(state[2]), .O(n11));
    defparam equal_1562_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hf7ff;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i23424_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39188));
    defparam i23424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_965 (.I0(state[3]), .I1(state[1]), .I2(state[2]), 
            .I3(\state[0] ), .O(n62901));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_965.LUT_INIT = 16'h1110;
    SB_LUT4 i3_4_lut_adj_966 (.I0(n27612), .I1(\state[0] ), .I2(state[2]), 
            .I3(state[3]), .O(n28819));
    defparam i3_4_lut_adj_966.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut_adj_967 (.I0(state[3]), .I1(n68477), .I2(n61685), 
            .I3(\state[0] ), .O(n27612));
    defparam i1_4_lut_adj_967.LUT_INIT = 16'h0544;
    SB_LUT4 i44533_3_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[3]), .O(n60736));
    defparam i44533_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52340_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(n6707), 
            .I3(GND_net), .O(n68477));
    defparam i52340_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_4_lut_adj_968 (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5006), 
            .I2(n11), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'h2a2f;
    SB_LUT4 i54509_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(state[3]), 
            .I3(state[2]), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(44[32:47])
    defparam i54509_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i54664_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5006), 
            .I2(GND_net), .I3(GND_net), .O(n39323));
    defparam i54664_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2_3_lut_4_lut_adj_969 (.I0(state[2]), .I1(state[3]), .I2(n6783[1]), 
            .I3(state[1]), .O(n62540));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_969.LUT_INIT = 16'h1000;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_970 (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_971 (.I0(n10_adj_5), .I1(counter[4]), .I2(counter[3]), 
            .I3(counter[5]), .O(n63401));   // verilog/i2c_controller.v(110[10:22])
    defparam i3_4_lut_adj_971.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_972 (.I0(counter[7]), .I1(counter[0]), .I2(n63401), 
            .I3(counter[6]), .O(n6707));   // verilog/i2c_controller.v(110[10:22])
    defparam i3_4_lut_adj_972.LUT_INIT = 16'hfffe;
    SB_LUT4 i54655_3_lut (.I0(n6714), .I1(n15), .I2(n39034), .I3(GND_net), 
            .O(n39496));
    defparam i54655_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i54522_4_lut (.I0(state_7__N_4109), .I1(n6707), .I2(n11_adj_5005), 
            .I3(n39032), .O(n6714));
    defparam i54522_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_973 (.I0(n11_adj_5012), .I1(n11_adj_5006), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4126[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_973.LUT_INIT = 16'h5575;
    SB_LUT4 i1_2_lut_3_lut_adj_974 (.I0(enable), .I1(\state_7__N_4110[0] ), 
            .I2(enable_slow_N_4213), .I3(GND_net), .O(n27553));
    defparam i1_2_lut_3_lut_adj_974.LUT_INIT = 16'haeae;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[3]), .I3(state[2]), .O(n11_adj_5012));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (setpoint, GND_net, \Kp[1] , \Kp[0] , \Kp[2] , 
            \Ki[4] , n358, PWMLimit, \motor_state[9] , \Kp[3] , \Kp[4] , 
            \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , duty, n39420, 
            \Kp[10] , \Kp[11] , \Kp[12] , n284, IntegralLimit, n258, 
            n359, \Ki[0] , control_update, n22, \Ki[3] , n348, n337, 
            n338, n339, n341, n342, n343, n344, n345, clk16MHz, 
            reset, n349, n350, n351, n352, n353, n354, n355, 
            n356, n357, \control_mode[7] , n17, n48532, \control_mode[1] , 
            \control_mode[0] , \motor_state[8] , n238, \PID_CONTROLLER.integral , 
            \motor_state[7] , n336, \motor_state[6] , \motor_state[5] , 
            \Ki[5] , \motor_state[4] , \Ki[6] , n290, n39, \Ki[7] , 
            \Ki[8] , \Ki[9] , \Ki[10] , deadband, \Ki[11] , \Ki[12] , 
            n29864, n29863, n29862, n29861, n29860, n29859, n29858, 
            n29857, n29856, n29855, n29854, n29853, n29852, n29851, 
            n29850, n29849, n29848, n29847, n29846, n29845, n29844, 
            n29843, n29839, n29097, \Ki[13] , \Ki[14] , \Ki[15] , 
            \Ki[1] , \Ki[2] , n346, n347, n34584, n34686, VCC_net, 
            \motor_state[3] , \motor_state[2] , \motor_state[1] , \Kp[13] , 
            n17_adj_1, \motor_state[22] , \motor_state[21] , \motor_state[20] , 
            \motor_state[19] , \motor_state[18] , \motor_state[17] , \motor_state[16] , 
            \motor_state[15] , \motor_state[14] , \motor_state[13] , \motor_state[12] , 
            n3, \motor_state[10] , \Kp[14] , n20628, n20682, n20719, 
            n34395, n6, \Kp[15] , \encoder1_position_scaled[0] , n15, 
            n68243, n15_adj_2, n53436, n131, n204, n4, n4_adj_3, 
            n8, n12, n20, n31, n37, n34791) /* synthesis syn_module_defined=1 */ ;
    input [23:0]setpoint;
    input GND_net;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Ki[4] ;
    output n358;
    input [23:0]PWMLimit;
    input \motor_state[9] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    output [23:0]duty;
    output n39420;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    output n284;
    input [23:0]IntegralLimit;
    output n258;
    output n359;
    input \Ki[0] ;
    output control_update;
    input n22;
    input \Ki[3] ;
    output n348;
    output n337;
    output n338;
    output n339;
    output n341;
    output n342;
    output n343;
    output n344;
    output n345;
    input clk16MHz;
    input reset;
    output n349;
    output n350;
    output n351;
    output n352;
    output n353;
    output n354;
    output n355;
    output n356;
    output n357;
    input \control_mode[7] ;
    input n17;
    input n48532;
    input \control_mode[1] ;
    input \control_mode[0] ;
    input \motor_state[8] ;
    output n238;
    output [23:0]\PID_CONTROLLER.integral ;
    input \motor_state[7] ;
    output n336;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \Ki[5] ;
    input \motor_state[4] ;
    input \Ki[6] ;
    output n290;
    input n39;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input [23:0]deadband;
    input \Ki[11] ;
    input \Ki[12] ;
    input n29864;
    input n29863;
    input n29862;
    input n29861;
    input n29860;
    input n29859;
    input n29858;
    input n29857;
    input n29856;
    input n29855;
    input n29854;
    input n29853;
    input n29852;
    input n29851;
    input n29850;
    input n29849;
    input n29848;
    input n29847;
    input n29846;
    input n29845;
    input n29844;
    input n29843;
    input n29839;
    input n29097;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Ki[1] ;
    input \Ki[2] ;
    output n346;
    output n347;
    input n34584;
    input n34686;
    input VCC_net;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \Kp[13] ;
    input n17_adj_1;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input n3;
    input \motor_state[10] ;
    input \Kp[14] ;
    input n20628;
    input n20682;
    output n20719;
    input n34395;
    input n6;
    input \Kp[15] ;
    input \encoder1_position_scaled[0] ;
    input n15;
    input n68243;
    input n15_adj_2;
    input n53436;
    input n131;
    input n204;
    output n4;
    input n4_adj_3;
    output n8;
    input n12;
    output n20;
    input n31;
    input n37;
    input n34791;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n9971, n68485, n4743, n72353, n71310, n43, n42;
    wire [23:0]n207;
    
    wire n107;
    wire [23:0]n535;
    wire [23:0]n455;
    
    wire n72356;
    wire [11:0]n19328;
    wire [10:0]n19637;
    
    wire n326, n54069, n38, n180, n70808, n70741, n71124, n296, 
        n54070;
    wire [43:0]n360;
    wire [47:0]n1;
    
    wire n53655, n71125, n53609;
    wire [23:0]n1_adj_5001;
    
    wire n253, n54068, n68484, n72347, n253_adj_4434, n326_adj_4435, 
        n53656, n72350, n399, n105, n472, n545, n618, n691, 
        n68483, n72341, n72344, n68482, n72335, n72338, n764, 
        n122, n53, n837, n195, n910, n53654, n268, n341_c, n414, 
        n487, n560;
    wire [23:0]n233;
    wire [23:0]n285;
    wire [23:0]n310;
    
    wire n5083, n68427, n7063, n180_adj_4436, n54067, n68428, n38_adj_4438, 
        n107_adj_4439, counter_31__N_3714, n53653, n45, n39_c, n41, 
        n43_adj_4443, n37_c, n53652, n35, n29, n31_c, n33, n12_c, 
        n25205, n53610, n21, n19, n17_adj_4445, n9, n69480, n27, 
        n15_c, n13, n11, n69464, n12_adj_4446, n53651, n10, n30, 
        n53608, n68506, n69502, n70349, n25, n23, n71263, n70727, 
        n71388, n16, n6_c, n70950, n70951, n8_c, n24, n69428, 
        n69392, n70774, n69644, n53650, n72035, n4_adj_4448, n72038, 
        n70948, n70949, n53649, n53648, n69459, n69455, n71265, 
        n69646, n71488, n71489, n71460, n53647, n69437, n71315, 
        n69652, n71317, n131_c, n72029, n41_adj_4449, n39_adj_4450, 
        n37_adj_4451, n35_adj_4452, n31_adj_4453, n33_adj_4454, n29_adj_4455, 
        n27_adj_4456, n45_adj_4457, n23_adj_4458, n25_adj_4459, n72032, 
        n43_adj_4460, n5_adj_4461, n54838, n39142, n21_adj_4462, n19_adj_4463, 
        n17_adj_4464, n9_adj_4465, n68843, n15_adj_4466, n13_adj_4467, 
        n11_adj_4468, n68837, n12_adj_4469;
    wire [6:0]n20478;
    wire [5:0]n20574;
    
    wire n54051, n54050, n54049, n10_adj_4470, n39_adj_4471, n41_adj_4472, 
        n54048, n30_adj_4473, n54047, n45_adj_4474, n53646;
    wire [11:0]n19468;
    wire [10:0]n19754;
    
    wire n54450, n54046, n54449, n33_adj_4475, n37_adj_4476, n54448, 
        n15_adj_4477, n17_adj_4478, n19_adj_4479, n53607, n53645, 
        n54447, n53644, n43_adj_4480, n54446, n53815, n54445, n68857, 
        n69865, n54444, n53814, n53813, n54443, n54442, n27_adj_4481, 
        n54441, n53812, n54440, n53643, n29_adj_4482, n53811, n53810, 
        n69861, n71160, n70459, n31_adj_4484, n71347;
    wire [9:0]n19898;
    
    wire n840, n54031, n767, n54030, n53809, n53642, n53641, n21_adj_4486;
    wire [0:0]n10332;
    wire [21:0]n10937;
    
    wire n54432, n54431, n694, n54029, n16_adj_4487, n53606, n54430, 
        n23_adj_4488, n54429, n25_adj_4489, n54428, n9_adj_4490, n54427, 
        n6_adj_4491, n70479, n54426, n621, n54028, n53808, n70480, 
        n11_adj_4493, n8_adj_4494, n54425, n13_adj_4495, n35_adj_4496, 
        n69358, n1096, n54424, n68426, n72011, n548_adj_4497, n54027, 
        n72014, n69343, n12_adj_4498, n68389, n71999, n72002, n1023, 
        n54423, n475_adj_4499, n54026, n10_adj_4500, n30_adj_4501, 
        n53807, n24_adj_4503, n69380, n70274, n70266, n68798, n71249, 
        n68796, n70786, n950, n54422, n68388, n71993, n70679, 
        n71384, n877, n54421, n804, n54420, n16_adj_4504, n402_adj_4505, 
        n54025, n71996, n69704, n731, n54419, n658, n54418, n6_adj_4506, 
        n70944, n70945, n585, n54417, n512, n54416, n439_adj_4507, 
        n54415, n329_adj_4508, n54024, n53806, n53640, n366, n54414, 
        n293_adj_4510, n54413, n256, n54023, n8_adj_4511, n24_adj_4512, 
        n53605, n69287, n220, n54412, n369, n68486, n68489, n53805, 
        n4_adj_4514, n53639, n147, n54411, n70477, n68490, n68491, 
        n5_adj_4515, n74, n183, n54022, n70478;
    wire [20:0]n12545;
    
    wire n54410, n41_adj_4516, n110, n54409, n69277, n70776, n68827, 
        n54408, n68390, n71981, n54407, n68824, n71164, n69706, 
        n69654;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n4_adj_4518, n54406, n72176, n70942, n68455, n68492, n54405, 
        n54404, n1099, n54403, n70943, n69333, n69326, n71267, 
        n69656, n1026, n54402, n71490, n953, n54401, n71491, n53638, 
        n880, n54400, n53804, n71447, n71448, n71458, n71361, 
        n14, n807, n54399, n68680, n71984, n68802, n71074, n69295, 
        n734, n54398, n661, n54397, n588, n54396, n71319, n515, 
        n54395, n53803, n69712, n69662, n71321, n442_adj_4521, n54394, 
        n71337, n41_adj_4522, n508, n4_adj_4523, n45_adj_4524, n54848, 
        n5190, n43_adj_4525, n27_adj_4527, n29_adj_4528, n31_adj_4529, 
        n21_adj_4530, n23_adj_4531, n25_adj_4532, n33_adj_4533, n37_adj_4534, 
        n15_adj_4535, n17_adj_4536, n19_adj_4537, n35_adj_4538, n53604, 
        n9_adj_4539, n11_adj_4540, n13_adj_4541, n69249, n69228, n12_adj_4542, 
        n10_adj_4543, n30_adj_4544, n69269, n70197, n70187, n71966, 
        n71894, n71882, n71864, n71858, n71231, n70639, n71380, 
        n71972, n71888, n71846, n72386, n72380, n72374, n72368, 
        n72362, n16_adj_4545, n6_adj_4546, n70938, n70939, n8_adj_4547, 
        n24_adj_4548, n69184, n69163, n70778, n69664, n4_adj_4549, 
        n70936, n70937, n69213, n72383, n69211, n71269, n69666, 
        n71492, n71493, n72173, n72377, n72371, n72365, n71456, 
        n69190, n71323, n72359, n9_adj_4551, n11_adj_4552, n13_adj_4553, 
        n15_adj_4554, n21_adj_4555, n19_adj_4556, n17_adj_4557, n11_adj_4558, 
        n13_adj_4559, n15_adj_4560, n54393, n9_adj_4561, n17_adj_4562, 
        n19_adj_4563, n21_adj_4564, n23_adj_4565, n25_adj_4566, n27_adj_4567, 
        n29_adj_4568, n33_adj_4569, n54392, n69672, n71325;
    wire [8:0]n20115;
    
    wire n770, n54009, n68266, n68252, n68368, n71969, n223_adj_4571, 
        n54391, n697, n54008, n68271, n68284, n68343, n68296, 
        n150, n54390, n8_adj_4572, n77;
    wire [0:0]n10961;
    wire [21:0]n11420;
    
    wire n54827, n54826, n53802, n53637, n54825;
    wire [19:0]n13820;
    
    wire n54389, n624, n54007, n53636, n54824, n68372, n54823, 
        n399_adj_4574, n54822, n54821, n472_adj_4575, n545_adj_4576, 
        n618_adj_4577, n54820, n691_adj_4578, n764_adj_4579, n1096_adj_4580, 
        n54819, n1023_adj_4581, n54818, n837_adj_4582, n54388, n950_adj_4583, 
        n54817, n910_adj_4584, n877_adj_4585, n54816, n54387, n551_adj_4586, 
        n54006, n804_adj_4587, n54815, n104, n35_adj_4588, n54386, 
        n478_adj_4589, n54005, n177, n731_adj_4590, n54814, n250_adj_4591, 
        n658_adj_4592, n54813, n323_adj_4593, n396_adj_4594, n585_adj_4595, 
        n54812, n512_adj_4596, n54811, n439_adj_4597, n54810, n469_adj_4598, 
        n542_adj_4599, n366_adj_4600, n54809, n615, n293_adj_4601, 
        n54808, n688, n220_adj_4602, n54807, n761, n147_adj_4603, 
        n54806, n834, n54385, n5_adj_4604, n74_adj_4605;
    wire [20:0]n12982;
    
    wire n54805, n54804, n54384, n54803, n907, n54802, n1102, 
        n54383, n54801, n54800, n1029, n54382, n980, n54799, n1099_adj_4606, 
        n54798, n956, n54381, n119, n883, n54380, n50, n1026_adj_4607, 
        n54797, n810, n54379, n953_adj_4608, n54796, n737, n54378, 
        n880_adj_4609, n54795, n664, n54377, n807_adj_4610, n54794, 
        n734_adj_4611, n54793, n192, n265, n661_adj_4612, n54792, 
        n591, n54376, n588_adj_4613, n54791, n515_adj_4614, n54790, 
        n518, n54375, n442_adj_4615, n54789, n445_adj_4616, n54374, 
        n338_adj_4617, n369_adj_4618, n54788, n372, n54373, n411, 
        n296_adj_4619, n54787, n299_adj_4620, n54372, n223_adj_4621, 
        n54786, n53801, n226_adj_4623, n54371, n150_adj_4624, n54785, 
        n153, n54370, n484, n557_adj_4625, n8_adj_4626, n77_adj_4627;
    wire [19:0]n14216;
    
    wire n54784, n54783, n11_adj_4628, n80;
    wire [18:0]n14929;
    
    wire n54369, n54782, n54368, n54781, n54367, n54366, n54780, 
        n54365, n630, n1105, n54364, n54779, n1102_adj_4629, n54778, 
        n1032, n54363, n1029_adj_4630, n54777, n959, n54362, n886, 
        n54361, n956_adj_4631, n54776, n813, n54360, n883_adj_4632, 
        n54775, n740, n54359, n810_adj_4633, n54774, n667, n54358, 
        n737_adj_4634, n54773, n594, n54357, n664_adj_4635, n54772, 
        n521, n54356, n591_adj_4636, n54771, n448_adj_4637, n54355, 
        n375, n54354, n518_adj_4638, n54770, n302_adj_4639, n54353, 
        n445_adj_4640, n54769, n372_adj_4641, n54768, n229, n54352, 
        n299_adj_4642, n54767, n156, n54351, n101, n32, n226_adj_4643, 
        n54766, n14_adj_4644, n83;
    wire [9:0]n19994;
    
    wire n840_adj_4645, n54350, n174, n153_adj_4646, n54765, n767_adj_4647, 
        n54349, n694_adj_4648, n54348, n11_adj_4649, n80_adj_4650, 
        n621_adj_4651, n54347;
    wire [6:0]n20433;
    wire [5:0]n20542;
    
    wire n560_adj_4652, n54764, n487_adj_4653, n54763, n548_adj_4654, 
        n54346, n414_adj_4655, n54762, n475_adj_4656, n54345, n402_adj_4657, 
        n54344, n53800, n53635, n329_adj_4659, n54343, n341_adj_4660, 
        n54761, n256_adj_4661, n54342, n247_adj_4662, n183_adj_4663, 
        n54341, n268_adj_4664, n54760, n41_adj_4665, n110_adj_4666, 
        n320_adj_4667, n393_adj_4668, n195_adj_4669, n54759, n466_adj_4670, 
        n53_adj_4671, n122_adj_4672, n405, n54004, n53634, n332_adj_4673, 
        n54003;
    wire [18:0]n15286;
    
    wire n54758, n54757, n54756, n53799, n539_adj_4674, n612, n685, 
        n54755, n259, n54002, n186, n54001, n54754, n44, n113, 
        n1105_adj_4675, n54753, n1032_adj_4676, n54752, n758, n831, 
        n959_adj_4677, n54751, n904, n977, n886_adj_4678, n54750, 
        n813_adj_4679, n54749, n740_adj_4680, n54748, n1050, n53798, 
        n667_adj_4682, n54747;
    wire [17:0]n15902;
    
    wire n54317, n54316, n98, n29_adj_4683, n171, n244_adj_4684, 
        n317_adj_4685, n390_adj_4686, n594_adj_4687, n54746, n463_adj_4688, 
        n536_adj_4689, n54315, n609, n521_adj_4690, n54745, n54314, 
        n53797, n682, n1108, n54313, n1035, n54312, n448_adj_4691, 
        n54744, n962, n54311, n755, n828, n901, n974, n375_adj_4692, 
        n54743, n1047, n889, n54310, n302_adj_4693, n54742, n816, 
        n54309, n229_adj_4694, n54741, n743, n54308, n53633, n53796, 
        n156_adj_4695, n54740, n670, n54307, n597, n54306, n53795, 
        n14_adj_4697, n83_adj_4698, n524, n54305, n451_adj_4699, n54304, 
        n1120, n116, n47, n53794, n189, n262;
    wire [17:0]n16222;
    
    wire n54739, n378, n54303, n54738, n305_adj_4701, n54302, n335, 
        n408, n232, n54301, n53793, n481, n54737, n159, n54300, 
        n17_adj_4703, n86, n54736, n554_adj_4704, n1108_adj_4705, 
        n54735, n627, n1035_adj_4706, n54734, n700, n962_adj_4707, 
        n54733, n95, n889_adj_4708, n54732, n26, n816_adj_4709, 
        n54731, n62402, n490, n53977, n743_adj_4710, n54730;
    wire [4:0]n20644;
    
    wire n417, n53976, n168, n241_adj_4711, n314_adj_4712, n387_adj_4713, 
        n670_adj_4714, n54729, n344_adj_4715, n53975, n460_adj_4716, 
        n271, n53974, n597_adj_4717, n54728, n53632, n198, n53973, 
        n533, n56, n125, n606, n524_adj_4718, n54727;
    wire [7:0]n20292;
    
    wire n700_adj_4719, n53972, n627_adj_4720, n53971, n451_adj_4721, 
        n54726, n554_adj_4722, n53970, n47_adj_4723;
    wire [23:0]n1_adj_5002;
    
    wire n53792, n679, n378_adj_4725, n54725;
    wire [23:0]n36;
    
    wire n53791, n53631, n752, n481_adj_4727, n53969, n53603, n408_adj_4728, 
        n53968;
    wire [16:0]n16743;
    
    wire n54278, n53602, n53601, n335_adj_4729, n53967, n53790, 
        n305_adj_4732, n54724, n54277, n262_adj_4733, n53966, n825, 
        n53789, n898, n232_adj_4735, n54723, n54276, n189_adj_4736, 
        n53965, n53788, n53630, n971, n1044, n159_adj_4739, n54722, 
        n1111, n54275, n47_adj_4740, n116_adj_4741, n1038, n54274, 
        n1117, n965, n54273, n53787, n17_adj_4744, n86_adj_4745, 
        n92, n892, n54272, n819, n54271, n53786;
    wire [16:0]n17028;
    
    wire n54721, n746, n54270, n53785, n54720, n673, n54269, n23_adj_4748, 
        n165, n238_adj_4749, n311, n384_adj_4750, n457_adj_4751, n530, 
        n603, n676, n600, n54268, n53784, n54719, n527, n54267, 
        n749, n822, n895, n1111_adj_4754, n54718, n454, n54266, 
        n968, n381, n54265, n1038_adj_4755, n54717, n53783, n308_adj_4757, 
        n54264, n53782, n1041, n965_adj_4759, n54716, n235_adj_4760, 
        n54263, n53629, n53781, n1114, n162, n54262, n892_adj_4762, 
        n54715, n20_adj_4763, n89, n53780, n113_adj_4765, n44_adj_4766, 
        n186_adj_4767, n259_adj_4768, n332_adj_4769, n405_adj_4770, 
        n478_adj_4771, n551_adj_4772, n624_adj_4773, n819_adj_4774, 
        n54714, n697_adj_4775, n770_adj_4776, n104_adj_4777, n35_adj_4778, 
        n177_adj_4779, n250_adj_4780, n323_adj_4781, n746_adj_4782, 
        n54713, n53779, n53778, n53628, n53777, n396_adj_4786, n469_adj_4787, 
        n542_adj_4788, n615_adj_4789, n688_adj_4790, n761_adj_4791, 
        n834_adj_4792, n41_adj_4793, n907_adj_4794, n980_adj_4795, n101_adj_4796, 
        n32_adj_4797, n39_adj_4798, n53627, n673_adj_4799, n54712, 
        n174_adj_4800;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire n53776, n600_adj_4802, n54711, n53775, n53626, n527_adj_4804, 
        n54710, n53774, n53625, n53773, n454_adj_4807, n54709, n53772, 
        n381_adj_4809, n54708, n308_adj_4810, n54707, n53771, n235_adj_4812, 
        n54706, n53624, n247_adj_4813, n53770, n162_adj_4815, n54705, 
        n20_adj_4816, n89_adj_4817;
    wire [15:0]n17714;
    
    wire n54704, n54703, n68301, n39485, n320_adj_4819;
    wire [23:0]n1_adj_5003;
    
    wire n53769, n53768, n53767, n1114_adj_4823, n54702, n53766, 
        n53765, n1041_adj_4826, n54701, n53623, n53622, n53764, 
        n53763, n53762, n968_adj_4831, n54700, n53761, n895_adj_4833, 
        n54699, n53621, n53760, n53620, n53759, n822_adj_4836, n54698, 
        n53758, n53757, n749_adj_4839, n54697, n53756, n676_adj_4841, 
        n54696, n393_adj_4842, n53755, n603_adj_4844, n54695, n466_adj_4845, 
        n37_adj_4846, n53619, n53754, n53618, n53753, n530_adj_4849, 
        n54694, n53752, n53751, n457_adj_4852, n54693, n384_adj_4853, 
        n54692, n311_adj_4854, n54691, n539_adj_4855, n53750, n53617, 
        n53749, n53616, n53748, n53747, n238_adj_4860, n54690, n35_adj_4861, 
        n612_adj_4862, n165_adj_4863, n54689, n53615, n23_adj_4865, 
        n92_adj_4866;
    wire [14:0]n18276;
    
    wire n54688, n685_adj_4867, n758_adj_4868, n53614, n1117_adj_4869, 
        n54687, n53613, n630_adj_4870, n53915, n557_adj_4871, n53914, 
        n1044_adj_4872, n54686, n484_adj_4873, n53913, n971_adj_4874, 
        n54685, n411_adj_4875, n53912, n898_adj_4876, n54684, n831_adj_4877, 
        n53612, n338_adj_4878, n53911, n825_adj_4879, n54683, n53611, 
        n904_adj_4881, n265_adj_4882, n53910, n752_adj_4883, n54682, 
        n192_adj_4884, n53909, n679_adj_4885, n54681, n50_adj_4886, 
        n119_adj_4887, n606_adj_4888, n54680, n533_adj_4889, n54679, 
        n977_adj_4890, n1050_adj_4891, n125_adj_4892, n460_adj_4893, 
        n54678, n56_adj_4894, n387_adj_4895, n54677, n314_adj_4896, 
        n54676, n241_adj_4897, n54675, n168_adj_4898, n54674, n26_adj_4899, 
        n95_adj_4900;
    wire [13:0]n18728;
    
    wire n1120_adj_4901, n54673, n1047_adj_4902, n54672, n974_adj_4903, 
        n54671, n901_adj_4904, n54670, n828_adj_4905, n54669, n755_adj_4906, 
        n54668, n682_adj_4907, n54667, n609_adj_4908, n54666, n536_adj_4909, 
        n54665, n463_adj_4910, n54664, n390_adj_4911, n54663, n317_adj_4912, 
        n54662, n244_adj_4913, n54661, n171_adj_4914, n54660, n29_adj_4915, 
        n98_adj_4916, n62699, n490_adj_4917, n54659;
    wire [4:0]n20623;
    
    wire n417_adj_4918, n54658, n344_adj_4919, n54657, n31_adj_4920, 
        n271_adj_4921, n54656, n198_adj_4922, n54655;
    wire [12:0]n19132;
    
    wire n54654, n54653, n54652, n54651, n54650, n54649, n54648, 
        n54647, n54646, n54645, n33_adj_4923, n54644, n54643, n54642, 
        n54641, n54640, n54639, n27_adj_4924, n54638, n54637, n54636, 
        n54635, n54634, n54633, n54632, n53669, n53668, n54631, 
        n53667, n53666, n24_adj_4925, n54630, n53665, n53664, n53663, 
        n53662, n53661, n53660, n53659, n53658, n53657, n68640, 
        n26_adj_4926, n29_adj_4927;
    wire [8:0]n20192;
    
    wire n54241, n54240, n54239, n54238, n54237, n54236, n54235, 
        n54234, n68652, n54233, n23_adj_4928, n43_adj_4929, n28;
    wire [15:0]n17462;
    
    wire n54213, n54212, n54211, n45_adj_4930, n54210, n54209, n54208, 
        n54207, n54206, n54205, n54204, n54203, n54202, n54201, 
        n54200, n54199, n54198, n25_adj_4931;
    wire [14:0]n18055;
    
    wire n54179, n54178, n54177, n54176, n54175, n54174, n54173, 
        n54172, n54171, n54170, n54169, n54168, n54167, n54166, 
        n54165;
    wire [7:0]n20352;
    
    wire n54164, n54163, n68957, n54162, n54161, n54160, n54159, 
        n54158, n54157, n54565, n54564;
    wire [13:0]n18536;
    
    wire n54139, n54138, n54137, n54563, n54136, n54135, n54562, 
        n54134, n6_adj_4932, n54133, n54561, n68939, n54132, n54131, 
        n54560, n54130, n54129, n54559, n54128, n54127, n54558, 
        n12_adj_4933, n54126, n54557;
    wire [12:0]n18967;
    
    wire n54125, n54124, n54556, n54123, n54122, n54555, n54121, 
        n54120, n54554, n54119, n54118, n54553, n54117, n54116, 
        n54115;
    wire [1:0]n20738;
    
    wire n53302, n54114, n54113, n62_adj_4934, n54096, n54095, n54094, 
        n54093, n10_adj_4935, n54092, n54091, n54090, n54089, n54088, 
        n64571, n54087, n54086, n54085, n54084, n54083, n54082, 
        n54081, n54080, n54079, n54078, n64575, n54077, n54076, 
        n54075, n54074, n54073, n64573, n53272, n64581, n4_adj_4936, 
        n8_adj_4937, n30_adj_4938, n68983, n69937, n69931, n71176, 
        n70491, n71364, n16_adj_4940, n6_adj_4941, n70916, n70917, 
        n8_adj_4942, n24_adj_4943, n65002, n23_adj_4944, n22_adj_4945, 
        n26_adj_4946, n68863, n69068, n68861, n70784, n69694, n4_adj_4949, 
        n4_adj_4950, n64619;
    wire [2:0]n20722;
    
    wire n4_adj_4951, n347_adj_4952, n6_adj_4953, n61219, n70914, 
        n64615, n68_adj_4954, n53327, n54844, n64605, n73003, n64609, 
        n8_adj_4955, n6_adj_4956, n69105, n70915, n54072, n68912, 
        n68903, n71060, n54071, n69696, n71445, n71446, n71363, 
        n68870, n71072, n69702, n71335, n45_adj_4957, n41_adj_4958, 
        n43_adj_4959, n39_adj_4960, n31_adj_4961, n37_adj_4962, n35_adj_4963, 
        n69062, n70015, n72524, n69987, n72519, n69054, n70007, 
        n72539, n70001, n72534, n16_adj_4964, n71963, n68985, n8_adj_4965, 
        n24_adj_4966, n69066, n72532, n69064, n72560, n70559;
    wire [3:0]n20680;
    
    wire n72557, n70009, n70970, n69036, n72522, n70549, n72551, 
        n71192, n72513, n71463, n72510, n69124, n12_adj_4967, n10_adj_4968, 
        n30_adj_4969, n69161, n70099, n70091, n71214, n70593, n71372, 
        n16_adj_4970, n8_adj_4971, n24_adj_4972, n6_adj_4973, n70930, 
        n70931, n69136, n69072, n70780, n69674, n4_adj_4974, n70920, 
        n70921, n12_adj_4975, n69017;
    wire [2:0]n20717;
    
    wire n72545, n10_adj_4976, n30_adj_4977, n4_adj_4978, n69026, 
        n71273, n69686, n71496, n71497, n71452, n6_adj_4979, n70922, 
        n70923, n68987, n72507, n70782, n69684, n68991, n71331, 
        n69692, n71333, n4_adj_4982, n70928, n70929, n69114, n71271, 
        n69676, n71891, n71494, n71495, n71885, n71454, n71879, 
        n69076, n71861, n71327, n69682, n71334, n71329, n39_adj_4984, 
        n71855, n41_adj_4985, n17_adj_4986, n70407, n16_adj_4989, 
        n70409, n71843, n33_adj_4992, n35_adj_4993, n25_adj_4994, 
        n27_adj_4995, n29_adj_4996, n23_adj_4997, n68656, n68644, 
        n30_adj_4999, n34, n71399, n71400;
    
    SB_LUT4 n9971_bdd_4_lut_55175 (.I0(n9971), .I1(n68485), .I2(setpoint[3]), 
            .I3(n4743), .O(n72353));
    defparam n9971_bdd_4_lut_55175.LUT_INIT = 16'he4aa;
    SB_LUT4 i53981_3_lut (.I0(n71310), .I1(setpoint[21]), .I2(n43), .I3(GND_net), 
            .O(n42));   // verilog/motorControl.v(45[16:33])
    defparam i53981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n72353_bdd_4_lut (.I0(n72353), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4743), .O(n72356));
    defparam n72353_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5095_5_lut (.I0(GND_net), .I1(n19637[2]), .I2(n326), .I3(n54069), 
            .O(n19328[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54034_4_lut (.I0(n42), .I1(n70808), .I2(n43), .I3(n70741), 
            .O(n71124));   // verilog/motorControl.v(45[16:33])
    defparam i54034_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5095_5 (.CI(n54069), .I0(n19637[2]), .I1(n326), .CO(n54070));
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n1[9]), .I3(n53655), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54035_3_lut (.I0(n71124), .I1(setpoint[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n71125));   // verilog/motorControl.v(45[16:33])
    defparam i54035_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n53609), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5095_4_lut (.I0(GND_net), .I1(n19637[1]), .I2(n253), .I3(n54068), 
            .O(n19328[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9971_bdd_4_lut_55170 (.I0(n9971), .I1(n68484), .I2(setpoint[2]), 
            .I3(n4743), .O(n72347));
    defparam n9971_bdd_4_lut_55170.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4434));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4435));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_25_11 (.CI(n53655), .I0(n360[9]), .I1(n1[9]), .CO(n53656));
    SB_LUT4 n72347_bdd_4_lut (.I0(n72347), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4743), .O(n72350));
    defparam n72347_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53683_3_lut (.I0(n71125), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i53683_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23654_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n39420));   // verilog/motorControl.v(42[14] 73[8])
    defparam i23654_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n9971_bdd_4_lut_55165 (.I0(n9971), .I1(n68483), .I2(setpoint[1]), 
            .I3(n4743), .O(n72341));
    defparam n9971_bdd_4_lut_55165.LUT_INIT = 16'he4aa;
    SB_LUT4 n72341_bdd_4_lut (.I0(n72341), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4743), .O(n72344));
    defparam n72341_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9971_bdd_4_lut_55160 (.I0(n9971), .I1(n68482), .I2(setpoint[0]), 
            .I3(n4743), .O(n72335));
    defparam n9971_bdd_4_lut_55160.LUT_INIT = 16'he4aa;
    SB_LUT4 n72335_bdd_4_lut (.I0(n72335), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4743), .O(n72338));
    defparam n72335_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n1[8]), .I3(n53654), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_c));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n359));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n359), .I2(GND_net), .I3(GND_net), 
            .O(n1[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51672_2_lut (.I0(PWMLimit[21]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68427));
    defparam i51672_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(control_update), .I1(n22), .I2(n105), .I3(GND_net), 
            .O(n7063));
    defparam i2_3_lut.LUT_INIT = 16'h2020;
    SB_CARRY add_25_10 (.CI(n53654), .I0(n360[8]), .I1(n1[8]), .CO(n53655));
    SB_CARRY add_5095_4 (.CI(n54068), .I0(n19637[1]), .I1(n253), .CO(n54069));
    SB_LUT4 i51815_2_lut (.I0(PWMLimit[2]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68484));
    defparam i51815_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5095_3_lut (.I0(GND_net), .I1(n19637[0]), .I2(n180_adj_4436), 
            .I3(n54067), .O(n19328[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n310[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i22_3_lut (.I0(n310[21]), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n339));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i19_3_lut (.I0(n233[18]), .I1(n285[18]), .I2(n284), 
            .I3(GND_net), .O(n310[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51671_2_lut (.I0(PWMLimit[22]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68428));
    defparam i51671_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i19_3_lut (.I0(n310[18]), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n342));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n343));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5095_3 (.CI(n54067), .I0(n19637[0]), .I1(n180_adj_4436), 
            .CO(n54068));
    SB_LUT4 add_5095_2_lut (.I0(GND_net), .I1(n38_adj_4438), .I2(n107_adj_4439), 
            .I3(GND_net), .O(n19328[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n344));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n345));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5095_2 (.CI(GND_net), .I0(n38_adj_4438), .I1(n107_adj_4439), 
            .CO(n54067));
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n72338), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_LUT4 mux_21_i11_3_lut (.I0(n233[10]), .I1(n285[10]), .I2(n284), 
            .I3(GND_net), .O(n310[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i11_3_lut (.I0(n310[10]), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n349));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n1[7]), .I3(n53653), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n350));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n351));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n353));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n354));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n356));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n357));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_25_9 (.CI(n53653), .I0(n360[7]), .I1(n1[7]), .CO(n53654));
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4443));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n1[6]), .I3(n53652), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(\control_mode[7] ), .I1(n105), .I2(control_update), 
            .I3(n17), .O(n12_c));
    defparam i5_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i6_4_lut (.I0(n48532), .I1(n12_c), .I2(\control_mode[1] ), 
            .I3(\control_mode[0] ), .O(n25205));
    defparam i6_4_lut.LUT_INIT = 16'h4000;
    SB_CARRY add_25_8 (.CI(n53652), .I0(n360[6]), .I1(n1[6]), .CO(n53653));
    SB_CARRY sub_15_add_2_11 (.CI(n53609), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n53610));
    SB_LUT4 i52390_4_lut (.I0(n21), .I1(n19), .I2(n17_adj_4445), .I3(n9), 
            .O(n69480));
    defparam i52390_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52374_4_lut (.I0(n27), .I1(n15_c), .I2(n13), .I3(n11), 
            .O(n69464));
    defparam i52374_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4446));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n1[5]), .I3(n53651), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4446), .I1(n535[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_25_7 (.CI(n53651), .I0(n360[5]), .I1(n1[5]), .CO(n53652));
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n53608), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52412_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n68506), 
            .O(n69502));
    defparam i52412_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53259_4_lut (.I0(n19), .I1(n17_adj_4445), .I2(n15_c), .I3(n69502), 
            .O(n70349));
    defparam i53259_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i54173_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n70349), 
            .O(n71263));
    defparam i54173_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53637_4_lut (.I0(n31_c), .I1(n29), .I2(n27), .I3(n71263), 
            .O(n70727));
    defparam i53637_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54298_4_lut (.I0(n37_c), .I1(n35), .I2(n33), .I3(n70727), 
            .O(n71388));
    defparam i54298_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4443), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53860_3_lut (.I0(n6_c), .I1(n535[10]), .I2(n21), .I3(GND_net), 
            .O(n70950));   // verilog/motorControl.v(47[25:43])
    defparam i53860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53861_3_lut (.I0(n70950), .I1(n535[11]), .I2(n23), .I3(GND_net), 
            .O(n70951));   // verilog/motorControl.v(47[25:43])
    defparam i53861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4445), 
            .I3(GND_net), .O(n8_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16), .I1(n535[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52338_4_lut (.I0(n43_adj_4443), .I1(n25), .I2(n23), .I3(n69480), 
            .O(n69428));
    defparam i52338_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53684_4_lut (.I0(n24), .I1(n8_c), .I2(n45), .I3(n69392), 
            .O(n70774));   // verilog/motorControl.v(47[25:43])
    defparam i53684_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52554_3_lut (.I0(n70951), .I1(n535[12]), .I2(n25), .I3(GND_net), 
            .O(n69644));   // verilog/motorControl.v(47[25:43])
    defparam i52554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n1[4]), .I3(n53650), 
            .O(n455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n53650), .I0(n360[4]), .I1(n1[4]), .CO(n53651));
    SB_LUT4 n9971_bdd_4_lut_55021 (.I0(n9971), .I1(n68428), .I2(setpoint[22]), 
            .I3(n4743), .O(n72035));
    defparam n9971_bdd_4_lut_55021.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4448));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 n72035_bdd_4_lut (.I0(n72035), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4743), .O(n72038));
    defparam n72035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i53858_3_lut (.I0(n4_adj_4448), .I1(n535[13]), .I2(n27), .I3(GND_net), 
            .O(n70948));   // verilog/motorControl.v(47[25:43])
    defparam i53858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53859_3_lut (.I0(n70948), .I1(n535[14]), .I2(n29), .I3(GND_net), 
            .O(n70949));   // verilog/motorControl.v(47[25:43])
    defparam i53859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n1[3]), .I3(n53649), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_5 (.CI(n53649), .I0(n360[3]), .I1(n1[3]), .CO(n53650));
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n1[2]), .I3(n53648), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52369_4_lut (.I0(n33), .I1(n31_c), .I2(n29), .I3(n69464), 
            .O(n69459));
    defparam i52369_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54175_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n69455), 
            .O(n71265));   // verilog/motorControl.v(47[25:43])
    defparam i54175_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52556_3_lut (.I0(n70949), .I1(n535[15]), .I2(n31_c), .I3(GND_net), 
            .O(n69646));   // verilog/motorControl.v(47[25:43])
    defparam i52556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54398_4_lut (.I0(n69646), .I1(n71265), .I2(n35), .I3(n69459), 
            .O(n71488));   // verilog/motorControl.v(47[25:43])
    defparam i54398_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_25_4 (.CI(n53648), .I0(n360[2]), .I1(n1[2]), .CO(n53649));
    SB_LUT4 i54399_3_lut (.I0(n71488), .I1(n535[18]), .I2(n37_c), .I3(GND_net), 
            .O(n71489));   // verilog/motorControl.v(47[25:43])
    defparam i54399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54370_3_lut (.I0(n71489), .I1(n535[19]), .I2(n39_c), .I3(GND_net), 
            .O(n71460));   // verilog/motorControl.v(47[25:43])
    defparam i54370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n1[1]), .I3(n53647), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52347_4_lut (.I0(n43_adj_4443), .I1(n41), .I2(n39_c), .I3(n71388), 
            .O(n69437));
    defparam i52347_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54225_4_lut (.I0(n69644), .I1(n70774), .I2(n45), .I3(n69428), 
            .O(n71315));   // verilog/motorControl.v(47[25:43])
    defparam i54225_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52562_3_lut (.I0(n71460), .I1(n535[20]), .I2(n41), .I3(GND_net), 
            .O(n69652));   // verilog/motorControl.v(47[25:43])
    defparam i52562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54227_4_lut (.I0(n69652), .I1(n71315), .I2(n45), .I3(n69437), 
            .O(n71317));   // verilog/motorControl.v(47[25:43])
    defparam i54227_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54228_3_lut (.I0(n71317), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(GND_net), .O(n131_c));   // verilog/motorControl.v(47[25:43])
    defparam i54228_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n9971_bdd_4_lut_54907 (.I0(n9971), .I1(n68427), .I2(setpoint[21]), 
            .I3(n4743), .O(n72029));
    defparam n9971_bdd_4_lut_54907.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4449));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n455[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4450));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4451));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4452));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4453));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4454));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4455));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4456));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4457));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4458));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n455[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4459));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n72029_bdd_4_lut (.I0(n72029), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4743), .O(n72032));
    defparam n72029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4460));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n5_adj_4461), .I1(n54838), .I2(n7063), .I3(n39142), 
            .O(n4743));
    defparam i3_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i51684_2_lut (.I0(PWMLimit[3]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68485));
    defparam i51684_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51753_4_lut (.I0(n21_adj_4462), .I1(n19_adj_4463), .I2(n17_adj_4464), 
            .I3(n9_adj_4465), .O(n68843));
    defparam i51753_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51747_4_lut (.I0(n27_adj_4456), .I1(n15_adj_4466), .I2(n13_adj_4467), 
            .I3(n11_adj_4468), .O(n68837));
    defparam i51747_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_25_3 (.CI(n53647), .I0(n360[1]), .I1(n1[1]), .CO(n53648));
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n1[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4454), 
            .I3(GND_net), .O(n12_adj_4469));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_15_add_2_10 (.CI(n53608), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n53609));
    SB_LUT4 add_5195_8_lut (.I0(GND_net), .I1(n20574[5]), .I2(n560), .I3(n54051), 
            .O(n20478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_7_lut (.I0(GND_net), .I1(n20574[4]), .I2(n487), .I3(n54050), 
            .O(n20478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_7 (.CI(n54050), .I0(n20574[4]), .I1(n487), .CO(n54051));
    SB_LUT4 add_5195_6_lut (.I0(GND_net), .I1(n20574[3]), .I2(n414), .I3(n54049), 
            .O(n20478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n1[0]), .CO(n53647));
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4467), 
            .I3(GND_net), .O(n10_adj_4470));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n238), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4471));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4472));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5195_6 (.CI(n54049), .I0(n20574[3]), .I1(n414), .CO(n54050));
    SB_LUT4 add_5195_5_lut (.I0(GND_net), .I1(n20574[2]), .I2(n341_c), 
            .I3(n54048), .O(n20478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_5 (.CI(n54048), .I0(n20574[2]), .I1(n341_c), .CO(n54049));
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_4469), .I1(n535[17]), .I2(n35_adj_4452), 
            .I3(GND_net), .O(n30_adj_4473));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5195_4_lut (.I0(GND_net), .I1(n20574[1]), .I2(n268), .I3(n54047), 
            .O(n20478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4474));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5195_4 (.CI(n54047), .I0(n20574[1]), .I1(n268), .CO(n54048));
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n53646), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5105_13_lut (.I0(GND_net), .I1(n19754[10]), .I2(n910), 
            .I3(n54450), .O(n19468[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_3_lut (.I0(GND_net), .I1(n20574[0]), .I2(n195), .I3(n54046), 
            .O(n20478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_3 (.CI(n54046), .I0(n20574[0]), .I1(n195), .CO(n54047));
    SB_LUT4 add_5105_12_lut (.I0(GND_net), .I1(n19754[9]), .I2(n837), 
            .I3(n54449), .O(n19468[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_12 (.CI(n54449), .I0(n19754[9]), .I1(n837), .CO(n54450));
    SB_LUT4 add_5195_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n54046));
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4475));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n233[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4476));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5105_11_lut (.I0(GND_net), .I1(n19754[8]), .I2(n764), 
            .I3(n54448), .O(n19468[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_11 (.CI(n54448), .I0(n19754[8]), .I1(n764), .CO(n54449));
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4477));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4478));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4479));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n53607), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n53645), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5105_10_lut (.I0(GND_net), .I1(n19754[7]), .I2(n691), 
            .I3(n54447), .O(n19468[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_24 (.CI(n53645), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n53646));
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n53644), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_10 (.CI(n54447), .I0(n19754[7]), .I1(n691), .CO(n54448));
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4480));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5105_9_lut (.I0(GND_net), .I1(n19754[6]), .I2(n618), .I3(n54446), 
            .O(n19468[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_9 (.CI(n54446), .I0(n19754[6]), .I1(n618), .CO(n54447));
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[23]), 
            .I3(n53815), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5105_8_lut (.I0(GND_net), .I1(n19754[5]), .I2(n545), .I3(n54445), 
            .O(n19468[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_8 (.CI(n54445), .I0(n19754[5]), .I1(n545), .CO(n54446));
    SB_LUT4 i52775_4_lut (.I0(n13_adj_4467), .I1(n11_adj_4468), .I2(n9_adj_4465), 
            .I3(n68857), .O(n69865));
    defparam i52775_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_5105_7_lut (.I0(GND_net), .I1(n19754[4]), .I2(n472), .I3(n54444), 
            .O(n19468[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[22]), 
            .I3(n53814), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n53814), .I0(GND_net), .I1(n1_adj_5001[22]), 
            .CO(n53815));
    SB_CARRY add_16_23 (.CI(n53644), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n53645));
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[21]), 
            .I3(n53813), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_7 (.CI(n54444), .I0(n19754[4]), .I1(n472), .CO(n54445));
    SB_LUT4 add_5105_6_lut (.I0(GND_net), .I1(n19754[3]), .I2(n399), .I3(n54443), 
            .O(n19468[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_6 (.CI(n54443), .I0(n19754[3]), .I1(n399), .CO(n54444));
    SB_LUT4 add_5105_5_lut (.I0(GND_net), .I1(n19754[2]), .I2(n326_adj_4435), 
            .I3(n54442), .O(n19468[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4481));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_33_add_3_23 (.CI(n53813), .I0(GND_net), .I1(n1_adj_5001[21]), 
            .CO(n53814));
    SB_CARRY add_5105_5 (.CI(n54442), .I0(n19754[2]), .I1(n326_adj_4435), 
            .CO(n54443));
    SB_LUT4 add_5105_4_lut (.I0(GND_net), .I1(n19754[1]), .I2(n253_adj_4434), 
            .I3(n54441), .O(n19468[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_4 (.CI(n54441), .I0(n19754[1]), .I1(n253_adj_4434), 
            .CO(n54442));
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[20]), 
            .I3(n53812), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n53812), .I0(GND_net), .I1(n1_adj_5001[20]), 
            .CO(n53813));
    SB_LUT4 add_5105_3_lut (.I0(GND_net), .I1(n19754[0]), .I2(n180), .I3(n54440), 
            .O(n19468[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n53643), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_3 (.CI(n54440), .I0(n19754[0]), .I1(n180), .CO(n54441));
    SB_LUT4 add_5105_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n19468[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5105_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5105_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n54440));
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4482));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_16_22 (.CI(n53643), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n53644));
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[19]), 
            .I3(n53811), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_21 (.CI(n53811), .I0(GND_net), .I1(n1_adj_5001[19]), 
            .CO(n53812));
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[18]), 
            .I3(n53810), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52771_4_lut (.I0(n19_adj_4463), .I1(n17_adj_4464), .I2(n15_adj_4466), 
            .I3(n69865), .O(n69861));
    defparam i52771_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i54070_4_lut (.I0(n25_adj_4459), .I1(n23_adj_4458), .I2(n21_adj_4462), 
            .I3(n69861), .O(n71160));
    defparam i54070_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53369_4_lut (.I0(n31_adj_4453), .I1(n29_adj_4455), .I2(n27_adj_4456), 
            .I3(n71160), .O(n70459));
    defparam i53369_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4484));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54257_4_lut (.I0(n37_adj_4451), .I1(n35_adj_4452), .I2(n33_adj_4454), 
            .I3(n70459), .O(n71347));
    defparam i54257_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5118_12_lut (.I0(GND_net), .I1(n19898[9]), .I2(n840), 
            .I3(n54031), .O(n19637[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_20 (.CI(n53810), .I0(GND_net), .I1(n1_adj_5001[18]), 
            .CO(n53811));
    SB_LUT4 add_5118_11_lut (.I0(GND_net), .I1(n19898[8]), .I2(n767), 
            .I3(n54030), .O(n19637[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[17]), 
            .I3(n53809), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n53809), .I0(GND_net), .I1(n1_adj_5001[17]), 
            .CO(n53810));
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n53642), .O(n238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_9 (.CI(n53607), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n53608));
    SB_CARRY add_16_21 (.CI(n53642), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n53643));
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n53641), .O(n233[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_11 (.CI(n54030), .I0(n19898[8]), .I1(n767), .CO(n54031));
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n233[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4486));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n336), .I1(n10937[21]), .I2(GND_net), 
            .I3(n54432), .O(n10332[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n10937[20]), .I2(GND_net), 
            .I3(n54431), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_10_lut (.I0(GND_net), .I1(n19898[7]), .I2(n694), 
            .I3(n54029), .O(n19637[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_10 (.CI(n54029), .I0(n19898[7]), .I1(n694), .CO(n54030));
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4460), 
            .I3(GND_net), .O(n16_adj_4487));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n53606), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_23 (.CI(n54431), .I0(n10937[20]), .I1(GND_net), 
            .CO(n54432));
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n10937[19]), .I2(GND_net), 
            .I3(n54430), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4488));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_24_add_1225_22 (.CI(n54430), .I0(n10937[19]), .I1(GND_net), 
            .CO(n54431));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n10937[18]), .I2(GND_net), 
            .I3(n54429), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_21 (.CI(n54429), .I0(n10937[18]), .I1(GND_net), 
            .CO(n54430));
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4489));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n10937[17]), .I2(GND_net), 
            .I3(n54428), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n54428), .I0(n10937[17]), .I1(GND_net), 
            .CO(n54429));
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4490));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n10937[16]), .I2(GND_net), 
            .I3(n54427), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_19 (.CI(n54427), .I0(n10937[16]), .I1(GND_net), 
            .CO(n54428));
    SB_LUT4 i53389_3_lut (.I0(n6_adj_4491), .I1(n535[10]), .I2(n21_adj_4462), 
            .I3(GND_net), .O(n70479));   // verilog/motorControl.v(65[25:41])
    defparam i53389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n10937[15]), .I2(GND_net), 
            .I3(n54426), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_9_lut (.I0(GND_net), .I1(n19898[6]), .I2(n621), .I3(n54028), 
            .O(n19637[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_9 (.CI(n54028), .I0(n19898[6]), .I1(n621), .CO(n54029));
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[16]), 
            .I3(n53808), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53390_3_lut (.I0(n70479), .I1(n535[11]), .I2(n23_adj_4458), 
            .I3(GND_net), .O(n70480));   // verilog/motorControl.v(65[25:41])
    defparam i53390_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_18 (.CI(n54426), .I0(n10937[15]), .I1(GND_net), 
            .CO(n54427));
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4493));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4464), 
            .I3(GND_net), .O(n8_adj_4494));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n10937[14]), .I2(GND_net), 
            .I3(n54425), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_17 (.CI(n54425), .I0(n10937[14]), .I1(GND_net), 
            .CO(n54426));
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4495));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4496));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52268_4_lut (.I0(n21_adj_4486), .I1(n19_adj_4479), .I2(n17_adj_4478), 
            .I3(n9_adj_4490), .O(n69358));
    defparam i52268_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n10937[13]), .I2(n1096), 
            .I3(n54424), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9971_bdd_4_lut_54902 (.I0(n9971), .I1(n68426), .I2(setpoint[20]), 
            .I3(n4743), .O(n72011));
    defparam n9971_bdd_4_lut_54902.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5118_8_lut (.I0(GND_net), .I1(n19898[5]), .I2(n548_adj_4497), 
            .I3(n54027), .O(n19637[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n72011_bdd_4_lut (.I0(n72011), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4743), .O(n72014));
    defparam n72011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i52253_4_lut (.I0(n27_adj_4481), .I1(n15_adj_4477), .I2(n13_adj_4495), 
            .I3(n11_adj_4493), .O(n69343));
    defparam i52253_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33_adj_4475), 
            .I3(GND_net), .O(n12_adj_4498));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5118_8 (.CI(n54027), .I0(n19898[5]), .I1(n548_adj_4497), 
            .CO(n54028));
    SB_CARRY mult_24_add_1225_16 (.CI(n54424), .I0(n10937[13]), .I1(n1096), 
            .CO(n54425));
    SB_LUT4 n9971_bdd_4_lut_54887 (.I0(n9971), .I1(n68389), .I2(setpoint[19]), 
            .I3(n4743), .O(n71999));
    defparam n9971_bdd_4_lut_54887.LUT_INIT = 16'he4aa;
    SB_LUT4 n71999_bdd_4_lut (.I0(n71999), .I1(n535[19]), .I2(n455[19]), 
            .I3(n4743), .O(n72002));
    defparam n71999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n10937[12]), .I2(n1023), 
            .I3(n54423), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_7_lut (.I0(GND_net), .I1(n19898[4]), .I2(n475_adj_4499), 
            .I3(n54026), .O(n19637[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13_adj_4495), 
            .I3(GND_net), .O(n10_adj_4500));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12_adj_4498), .I1(n233[17]), .I2(n35_adj_4496), 
            .I3(GND_net), .O(n30_adj_4501));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n53808), .I0(GND_net), .I1(n1_adj_5001[16]), 
            .CO(n53809));
    SB_CARRY mult_24_add_1225_15 (.CI(n54423), .I0(n10937[12]), .I1(n1023), 
            .CO(n54424));
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[15]), 
            .I3(n53807), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_4487), .I1(n535[22]), .I2(n45_adj_4457), 
            .I3(GND_net), .O(n24_adj_4503));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53184_4_lut (.I0(n13_adj_4495), .I1(n11_adj_4493), .I2(n9_adj_4490), 
            .I3(n69380), .O(n70274));
    defparam i53184_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53176_4_lut (.I0(n19_adj_4479), .I1(n17_adj_4478), .I2(n15_adj_4477), 
            .I3(n70274), .O(n70266));
    defparam i53176_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_16_20 (.CI(n53641), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n53642));
    SB_LUT4 i51708_4_lut (.I0(n43_adj_4460), .I1(n25_adj_4459), .I2(n23_adj_4458), 
            .I3(n68843), .O(n68798));
    defparam i51708_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54159_4_lut (.I0(n25_adj_4489), .I1(n23_adj_4488), .I2(n21_adj_4486), 
            .I3(n70266), .O(n71249));
    defparam i54159_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53696_4_lut (.I0(n24_adj_4503), .I1(n8_adj_4494), .I2(n45_adj_4457), 
            .I3(n68796), .O(n70786));   // verilog/motorControl.v(65[25:41])
    defparam i53696_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n10937[11]), .I2(n950), 
            .I3(n54422), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9971_bdd_4_lut_54877 (.I0(n9971), .I1(n68388), .I2(setpoint[18]), 
            .I3(n4743), .O(n71993));
    defparam n9971_bdd_4_lut_54877.LUT_INIT = 16'he4aa;
    SB_LUT4 i53589_4_lut (.I0(n31_adj_4484), .I1(n29_adj_4482), .I2(n27_adj_4481), 
            .I3(n71249), .O(n70679));
    defparam i53589_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY mult_24_add_1225_14 (.CI(n54422), .I0(n10937[11]), .I1(n950), 
            .CO(n54423));
    SB_CARRY add_5118_7 (.CI(n54026), .I0(n19898[4]), .I1(n475_adj_4499), 
            .CO(n54027));
    SB_LUT4 i54294_4_lut (.I0(n37_adj_4476), .I1(n35_adj_4496), .I2(n33_adj_4475), 
            .I3(n70679), .O(n71384));
    defparam i54294_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n10937[10]), .I2(n877), 
            .I3(n54421), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_13 (.CI(n54421), .I0(n10937[10]), .I1(n877), 
            .CO(n54422));
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n10937[9]), .I2(n804), 
            .I3(n54420), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43_adj_4480), 
            .I3(GND_net), .O(n16_adj_4504));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5118_6_lut (.I0(GND_net), .I1(n19898[3]), .I2(n402_adj_4505), 
            .I3(n54025), .O(n19637[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_6 (.CI(n54025), .I0(n19898[3]), .I1(n402_adj_4505), 
            .CO(n54026));
    SB_LUT4 n71993_bdd_4_lut (.I0(n71993), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4743), .O(n71996));
    defparam n71993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY unary_minus_33_add_3_17 (.CI(n53807), .I0(GND_net), .I1(n1_adj_5001[15]), 
            .CO(n53808));
    SB_LUT4 i52614_3_lut (.I0(n70480), .I1(n535[12]), .I2(n25_adj_4459), 
            .I3(GND_net), .O(n69704));   // verilog/motorControl.v(65[25:41])
    defparam i52614_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_12 (.CI(n54420), .I0(n10937[9]), .I1(n804), 
            .CO(n54421));
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n10937[8]), .I2(n731), 
            .I3(n54419), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_11 (.CI(n54419), .I0(n10937[8]), .I1(n731), 
            .CO(n54420));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n10937[7]), .I2(n658), 
            .I3(n54418), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53854_3_lut (.I0(n6_adj_4506), .I1(n233[10]), .I2(n21_adj_4486), 
            .I3(GND_net), .O(n70944));   // verilog/motorControl.v(56[14:36])
    defparam i53854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53855_3_lut (.I0(n70944), .I1(n233[11]), .I2(n23_adj_4488), 
            .I3(GND_net), .O(n70945));   // verilog/motorControl.v(56[14:36])
    defparam i53855_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_10 (.CI(n54418), .I0(n10937[7]), .I1(n658), 
            .CO(n54419));
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n10937[6]), .I2(n585), 
            .I3(n54417), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_9 (.CI(n54417), .I0(n10937[6]), .I1(n585), 
            .CO(n54418));
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n10937[5]), .I2(n512), 
            .I3(n54416), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_8 (.CI(n54416), .I0(n10937[5]), .I1(n512), 
            .CO(n54417));
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n10937[4]), .I2(n439_adj_4507), 
            .I3(n54415), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_5_lut (.I0(GND_net), .I1(n19898[2]), .I2(n329_adj_4508), 
            .I3(n54024), .O(n19637[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_5 (.CI(n54024), .I0(n19898[2]), .I1(n329_adj_4508), 
            .CO(n54025));
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[14]), 
            .I3(n53806), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_16 (.CI(n53806), .I0(GND_net), .I1(n1_adj_5001[14]), 
            .CO(n53807));
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n53640), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_7 (.CI(n54415), .I0(n10937[4]), .I1(n439_adj_4507), 
            .CO(n54416));
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n10937[3]), .I2(n366), 
            .I3(n54414), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_19 (.CI(n53640), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n53641));
    SB_CARRY mult_24_add_1225_6 (.CI(n54414), .I0(n10937[3]), .I1(n366), 
            .CO(n54415));
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n10937[2]), .I2(n293_adj_4510), 
            .I3(n54413), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_4_lut (.I0(GND_net), .I1(n19898[1]), .I2(n256), .I3(n54023), 
            .O(n19637[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_8 (.CI(n53606), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n53607));
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_4478), 
            .I3(GND_net), .O(n8_adj_4511));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4504), .I1(n233[22]), .I2(n45_adj_4474), 
            .I3(GND_net), .O(n24_adj_4512));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n53605), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52197_4_lut (.I0(n43_adj_4480), .I1(n25_adj_4489), .I2(n23_adj_4488), 
            .I3(n69358), .O(n69287));
    defparam i52197_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_24_add_1225_5 (.CI(n54413), .I0(n10937[2]), .I1(n293_adj_4510), 
            .CO(n54414));
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n10937[1]), .I2(n220), 
            .I3(n54412), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51682_2_lut (.I0(PWMLimit[4]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68486));
    defparam i51682_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52399_2_lut (.I0(PWMLimit[5]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68489));
    defparam i52399_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_4 (.CI(n54412), .I0(n10937[1]), .I1(n220), 
            .CO(n54413));
    SB_CARRY add_5118_4 (.CI(n54023), .I0(n19898[1]), .I1(n256), .CO(n54024));
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[13]), 
            .I3(n53805), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_4514));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n53639), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n10937[0]), .I2(n147), 
            .I3(n54411), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53387_3_lut (.I0(n4_adj_4514), .I1(n535[13]), .I2(n27_adj_4456), 
            .I3(GND_net), .O(n70477));   // verilog/motorControl.v(65[25:41])
    defparam i53387_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51680_2_lut (.I0(PWMLimit[6]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68490));
    defparam i51680_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51569_2_lut (.I0(PWMLimit[7]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68491));
    defparam i51569_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_3 (.CI(n54411), .I0(n10937[0]), .I1(n147), 
            .CO(n54412));
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4515), .I2(n74), 
            .I3(GND_net), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5118_3_lut (.I0(GND_net), .I1(n19898[0]), .I2(n183), .I3(n54022), 
            .O(n19637[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53388_3_lut (.I0(n70477), .I1(n535[14]), .I2(n29_adj_4455), 
            .I3(GND_net), .O(n70478));   // verilog/motorControl.v(65[25:41])
    defparam i53388_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5_adj_4515), .I1(n74), 
            .CO(n54411));
    SB_LUT4 add_4527_23_lut (.I0(GND_net), .I1(n12545[20]), .I2(GND_net), 
            .I3(n54410), .O(n10937[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5118_3 (.CI(n54022), .I0(n19898[0]), .I1(n183), .CO(n54023));
    SB_LUT4 add_5118_2_lut (.I0(GND_net), .I1(n41_adj_4516), .I2(n110), 
            .I3(GND_net), .O(n19637[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5118_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_22_lut (.I0(GND_net), .I1(n12545[19]), .I2(GND_net), 
            .I3(n54409), .O(n10937[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53686_4_lut (.I0(n24_adj_4512), .I1(n8_adj_4511), .I2(n45_adj_4474), 
            .I3(n69277), .O(n70776));   // verilog/motorControl.v(56[14:36])
    defparam i53686_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4527_22 (.CI(n54409), .I0(n12545[19]), .I1(GND_net), 
            .CO(n54410));
    SB_CARRY add_5118_2 (.CI(GND_net), .I0(n41_adj_4516), .I1(n110), .CO(n54022));
    SB_LUT4 i51737_4_lut (.I0(n33_adj_4454), .I1(n31_adj_4453), .I2(n29_adj_4455), 
            .I3(n68837), .O(n68827));
    defparam i51737_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4527_21_lut (.I0(GND_net), .I1(n12545[18]), .I2(GND_net), 
            .I3(n54408), .O(n10937[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_21 (.CI(n54408), .I0(n12545[18]), .I1(GND_net), 
            .CO(n54409));
    SB_LUT4 n9971_bdd_4_lut_54872 (.I0(n9971), .I1(n68390), .I2(setpoint[12]), 
            .I3(n4743), .O(n71981));
    defparam n9971_bdd_4_lut_54872.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4527_20_lut (.I0(GND_net), .I1(n12545[17]), .I2(GND_net), 
            .I3(n54407), .O(n10937[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54074_4_lut (.I0(n30_adj_4473), .I1(n10_adj_4470), .I2(n35_adj_4452), 
            .I3(n68824), .O(n71164));   // verilog/motorControl.v(65[25:41])
    defparam i54074_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4527_20 (.CI(n54407), .I0(n12545[17]), .I1(GND_net), 
            .CO(n54408));
    SB_LUT4 i52616_3_lut (.I0(n70478), .I1(n535[15]), .I2(n31_adj_4453), 
            .I3(GND_net), .O(n69706));   // verilog/motorControl.v(65[25:41])
    defparam i52616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52564_3_lut (.I0(n70945), .I1(n233[12]), .I2(n25_adj_4489), 
            .I3(GND_net), .O(n69654));   // verilog/motorControl.v(56[14:36])
    defparam i52564_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR counter_2045_2046__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4518));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_4527_19_lut (.I0(GND_net), .I1(n12545[16]), .I2(GND_net), 
            .I3(n54406), .O(n10937[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n72176), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4527_19 (.CI(n54406), .I0(n12545[16]), .I1(GND_net), 
            .CO(n54407));
    SB_LUT4 i53852_3_lut (.I0(n4_adj_4518), .I1(n233[13]), .I2(n27_adj_4481), 
            .I3(GND_net), .O(n70942));   // verilog/motorControl.v(56[14:36])
    defparam i53852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52312_2_lut (.I0(PWMLimit[23]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68455));
    defparam i52312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51679_2_lut (.I0(PWMLimit[8]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68492));
    defparam i51679_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4527_18_lut (.I0(GND_net), .I1(n12545[15]), .I2(GND_net), 
            .I3(n54405), .O(n10937[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_18 (.CI(n54405), .I0(n12545[15]), .I1(GND_net), 
            .CO(n54406));
    SB_LUT4 add_4527_17_lut (.I0(GND_net), .I1(n12545[14]), .I2(GND_net), 
            .I3(n54404), .O(n10937[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_15 (.CI(n53805), .I0(GND_net), .I1(n1_adj_5001[13]), 
            .CO(n53806));
    SB_CARRY add_4527_17 (.CI(n54404), .I0(n12545[14]), .I1(GND_net), 
            .CO(n54405));
    SB_LUT4 add_4527_16_lut (.I0(GND_net), .I1(n12545[13]), .I2(n1099), 
            .I3(n54403), .O(n10937[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53853_3_lut (.I0(n70942), .I1(n233[14]), .I2(n29_adj_4482), 
            .I3(GND_net), .O(n70943));   // verilog/motorControl.v(56[14:36])
    defparam i53853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52243_4_lut (.I0(n33_adj_4475), .I1(n31_adj_4484), .I2(n29_adj_4482), 
            .I3(n69343), .O(n69333));
    defparam i52243_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54177_4_lut (.I0(n30_adj_4501), .I1(n10_adj_4500), .I2(n35_adj_4496), 
            .I3(n69326), .O(n71267));   // verilog/motorControl.v(56[14:36])
    defparam i54177_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_16_18 (.CI(n53639), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n53640));
    SB_LUT4 i52566_3_lut (.I0(n70943), .I1(n233[15]), .I2(n31_adj_4484), 
            .I3(GND_net), .O(n69656));   // verilog/motorControl.v(56[14:36])
    defparam i52566_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4527_16 (.CI(n54403), .I0(n12545[13]), .I1(n1099), .CO(n54404));
    SB_LUT4 add_4527_15_lut (.I0(GND_net), .I1(n12545[12]), .I2(n1026), 
            .I3(n54402), .O(n10937[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_7 (.CI(n53605), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n53606));
    SB_CARRY add_4527_15 (.CI(n54402), .I0(n12545[12]), .I1(n1026), .CO(n54403));
    SB_LUT4 i54400_4_lut (.I0(n69656), .I1(n71267), .I2(n35_adj_4496), 
            .I3(n69333), .O(n71490));   // verilog/motorControl.v(56[14:36])
    defparam i54400_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4527_14_lut (.I0(GND_net), .I1(n12545[11]), .I2(n953), 
            .I3(n54401), .O(n10937[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54401_3_lut (.I0(n71490), .I1(n233[18]), .I2(n37_adj_4476), 
            .I3(GND_net), .O(n71491));   // verilog/motorControl.v(56[14:36])
    defparam i54401_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4527_14 (.CI(n54401), .I0(n12545[11]), .I1(n953), .CO(n54402));
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n53638), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_13_lut (.I0(GND_net), .I1(n12545[10]), .I2(n880), 
            .I3(n54400), .O(n10937[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[12]), 
            .I3(n53804), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54357_4_lut (.I0(n69706), .I1(n71164), .I2(n35_adj_4452), 
            .I3(n68827), .O(n71447));   // verilog/motorControl.v(65[25:41])
    defparam i54357_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54358_3_lut (.I0(n71447), .I1(n535[18]), .I2(n37_adj_4451), 
            .I3(GND_net), .O(n71448));   // verilog/motorControl.v(65[25:41])
    defparam i54358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54368_3_lut (.I0(n71491), .I1(n238), .I2(n39_adj_4471), .I3(GND_net), 
            .O(n71458));   // verilog/motorControl.v(56[14:36])
    defparam i54368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54271_3_lut (.I0(n71448), .I1(n535[19]), .I2(n39_adj_4450), 
            .I3(GND_net), .O(n71361));   // verilog/motorControl.v(65[25:41])
    defparam i54271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i14_3_lut_3_lut (.I0(PWMLimit[7]), .I1(setpoint[7]), 
            .I2(setpoint[6]), .I3(GND_net), .O(n14));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i14_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_4527_13 (.CI(n54400), .I0(n12545[10]), .I1(n880), .CO(n54401));
    SB_LUT4 add_4527_12_lut (.I0(GND_net), .I1(n12545[9]), .I2(n807), 
            .I3(n54399), .O(n10937[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_12 (.CI(n54399), .I0(n12545[9]), .I1(n807), .CO(n54400));
    SB_LUT4 i51590_3_lut_4_lut (.I0(PWMLimit[7]), .I1(setpoint[7]), .I2(setpoint[6]), 
            .I3(PWMLimit[6]), .O(n68680));   // verilog/motorControl.v(45[16:33])
    defparam i51590_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n71981_bdd_4_lut (.I0(n71981), .I1(n535[12]), .I2(n455[12]), 
            .I3(n4743), .O(n71984));
    defparam n71981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51712_4_lut (.I0(n43_adj_4460), .I1(n41_adj_4449), .I2(n39_adj_4450), 
            .I3(n71347), .O(n68802));
    defparam i51712_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53984_4_lut (.I0(n69704), .I1(n70786), .I2(n45_adj_4457), 
            .I3(n68798), .O(n71074));   // verilog/motorControl.v(65[25:41])
    defparam i53984_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52205_4_lut (.I0(n43_adj_4480), .I1(n41_adj_4472), .I2(n39_adj_4471), 
            .I3(n71384), .O(n69295));
    defparam i52205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4527_11_lut (.I0(GND_net), .I1(n12545[8]), .I2(n734), 
            .I3(n54398), .O(n10937[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_11 (.CI(n54398), .I0(n12545[8]), .I1(n734), .CO(n54399));
    SB_LUT4 add_4527_10_lut (.I0(GND_net), .I1(n12545[7]), .I2(n661), 
            .I3(n54397), .O(n10937[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_10 (.CI(n54397), .I0(n12545[7]), .I1(n661), .CO(n54398));
    SB_LUT4 add_4527_9_lut (.I0(GND_net), .I1(n12545[6]), .I2(n588), .I3(n54396), 
            .O(n10937[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_9 (.CI(n54396), .I0(n12545[6]), .I1(n588), .CO(n54397));
    SB_LUT4 i54229_4_lut (.I0(n69654), .I1(n70776), .I2(n45_adj_4474), 
            .I3(n69287), .O(n71319));   // verilog/motorControl.v(56[14:36])
    defparam i54229_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4527_8_lut (.I0(GND_net), .I1(n12545[5]), .I2(n515), .I3(n54395), 
            .O(n10937[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_8 (.CI(n54395), .I0(n12545[5]), .I1(n515), .CO(n54396));
    SB_CARRY unary_minus_33_add_3_14 (.CI(n53804), .I0(GND_net), .I1(n1_adj_5001[12]), 
            .CO(n53805));
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[11]), 
            .I3(n53803), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52622_3_lut (.I0(n71361), .I1(n535[20]), .I2(n41_adj_4449), 
            .I3(GND_net), .O(n69712));   // verilog/motorControl.v(65[25:41])
    defparam i52622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52572_3_lut (.I0(n71458), .I1(n233[20]), .I2(n41_adj_4472), 
            .I3(GND_net), .O(n69662));   // verilog/motorControl.v(56[14:36])
    defparam i52572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54231_4_lut (.I0(n69662), .I1(n71319), .I2(n45_adj_4474), 
            .I3(n69295), .O(n71321));   // verilog/motorControl.v(56[14:36])
    defparam i54231_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4527_7_lut (.I0(GND_net), .I1(n12545[4]), .I2(n442_adj_4521), 
            .I3(n54394), .O(n10937[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i54247_4_lut (.I0(n69712), .I1(n71074), .I2(n45_adj_4457), 
            .I3(n68802), .O(n71337));   // verilog/motorControl.v(65[25:41])
    defparam i54247_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54232_3_lut (.I0(n71321), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i54232_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4522));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n508), .I1(n71337), .I2(n455[23]), .I3(n535[23]), 
            .O(n4_adj_4523));
    defparam i1_4_lut.LUT_INIT = 16'hbfab;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4524));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reduce_or_1169_i1_4_lut (.I0(n54848), .I1(n131_c), .I2(n4_adj_4523), 
            .I3(n25205), .O(n5190));
    defparam reduce_or_1169_i1_4_lut.LUT_INIT = 16'hce0a;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4525));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4527));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4528));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4529));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(n233[10]), .I1(n285[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4530));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4531));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4532));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4533));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(n233[18]), .I1(n285[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4534));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4535));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4536));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n72038), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4537));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4538));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n53604), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4539));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4540));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4541));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52159_4_lut (.I0(n21_adj_4530), .I1(n19_adj_4537), .I2(n17_adj_4536), 
            .I3(n9_adj_4539), .O(n69249));
    defparam i52159_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52138_4_lut (.I0(n27_adj_4527), .I1(n15_adj_4535), .I2(n13_adj_4541), 
            .I3(n11_adj_4540), .O(n69228));
    defparam i52138_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_4533), 
            .I3(GND_net), .O(n12_adj_4542));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4541), 
            .I3(GND_net), .O(n10_adj_4543));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4542), .I1(n285[17]), .I2(n35_adj_4538), 
            .I3(GND_net), .O(n30_adj_4544));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53107_4_lut (.I0(n13_adj_4541), .I1(n11_adj_4540), .I2(n9_adj_4539), 
            .I3(n69269), .O(n70197));
    defparam i53107_4_lut.LUT_INIT = 16'heeef;
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n72032), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i53097_4_lut (.I0(n19_adj_4537), .I1(n17_adj_4536), .I2(n15_adj_4535), 
            .I3(n70197), .O(n70187));
    defparam i53097_4_lut.LUT_INIT = 16'heeef;
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n72014), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n72002), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n71996), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n71966), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n71894), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n71882), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n71864), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n71858), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n71984), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 i54141_4_lut (.I0(n25_adj_4532), .I1(n23_adj_4531), .I2(n21_adj_4530), 
            .I3(n70187), .O(n71231));
    defparam i54141_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53549_4_lut (.I0(n31_adj_4529), .I1(n29_adj_4528), .I2(n27_adj_4527), 
            .I3(n71231), .O(n70639));
    defparam i53549_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54290_4_lut (.I0(n37_adj_4534), .I1(n35_adj_4538), .I2(n33_adj_4533), 
            .I3(n70639), .O(n71380));
    defparam i54290_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n71972), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n71888), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n71846), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n72386), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n72380), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n72374), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n72368), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n72362), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n72356), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n72350), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n72344), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_4525), 
            .I3(GND_net), .O(n16_adj_4545));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53848_3_lut (.I0(n6_adj_4546), .I1(n285[10]), .I2(n21_adj_4530), 
            .I3(GND_net), .O(n70938));   // verilog/motorControl.v(58[23:46])
    defparam i53848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53849_3_lut (.I0(n70938), .I1(n285[11]), .I2(n23_adj_4531), 
            .I3(GND_net), .O(n70939));   // verilog/motorControl.v(58[23:46])
    defparam i53849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_4536), 
            .I3(GND_net), .O(n8_adj_4547));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4545), .I1(n285[22]), .I2(n45_adj_4524), 
            .I3(GND_net), .O(n24_adj_4548));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52094_4_lut (.I0(n43_adj_4525), .I1(n25_adj_4532), .I2(n23_adj_4531), 
            .I3(n69249), .O(n69184));
    defparam i52094_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i53688_4_lut (.I0(n24_adj_4548), .I1(n8_adj_4547), .I2(n45_adj_4524), 
            .I3(n69163), .O(n70778));   // verilog/motorControl.v(58[23:46])
    defparam i53688_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52574_3_lut (.I0(n70939), .I1(n285[12]), .I2(n25_adj_4532), 
            .I3(GND_net), .O(n69664));   // verilog/motorControl.v(58[23:46])
    defparam i52574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_4549));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i53846_3_lut (.I0(n4_adj_4549), .I1(n285[13]), .I2(n27_adj_4527), 
            .I3(GND_net), .O(n70936));   // verilog/motorControl.v(58[23:46])
    defparam i53846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53847_3_lut (.I0(n70936), .I1(n285[14]), .I2(n29_adj_4528), 
            .I3(GND_net), .O(n70937));   // verilog/motorControl.v(58[23:46])
    defparam i53847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52123_4_lut (.I0(n33_adj_4533), .I1(n31_adj_4529), .I2(n29_adj_4528), 
            .I3(n69228), .O(n69213));
    defparam i52123_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9971_bdd_4_lut (.I0(n9971), .I1(n68492), .I2(setpoint[8]), 
            .I3(n4743), .O(n72383));
    defparam n9971_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i54179_4_lut (.I0(n30_adj_4544), .I1(n10_adj_4543), .I2(n35_adj_4538), 
            .I3(n69211), .O(n71269));   // verilog/motorControl.v(58[23:46])
    defparam i54179_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52576_3_lut (.I0(n70937), .I1(n285[15]), .I2(n31_adj_4529), 
            .I3(GND_net), .O(n69666));   // verilog/motorControl.v(58[23:46])
    defparam i52576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n72383_bdd_4_lut (.I0(n72383), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4743), .O(n72386));
    defparam n72383_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i54402_4_lut (.I0(n69666), .I1(n71269), .I2(n35_adj_4538), 
            .I3(n69213), .O(n71492));   // verilog/motorControl.v(58[23:46])
    defparam i54402_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54403_3_lut (.I0(n71492), .I1(n285[18]), .I2(n37_adj_4534), 
            .I3(GND_net), .O(n71493));   // verilog/motorControl.v(58[23:46])
    defparam i54403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9971_bdd_4_lut_55155 (.I0(n9971), .I1(n68455), .I2(setpoint[23]), 
            .I3(n4743), .O(n72173));
    defparam n9971_bdd_4_lut_55155.LUT_INIT = 16'he4aa;
    SB_LUT4 n72173_bdd_4_lut (.I0(n72173), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4743), .O(n72176));
    defparam n72173_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9971_bdd_4_lut_55195 (.I0(n9971), .I1(n68491), .I2(setpoint[7]), 
            .I3(n4743), .O(n72377));
    defparam n9971_bdd_4_lut_55195.LUT_INIT = 16'he4aa;
    SB_LUT4 n72377_bdd_4_lut (.I0(n72377), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4743), .O(n72380));
    defparam n72377_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9971_bdd_4_lut_55190 (.I0(n9971), .I1(n68490), .I2(setpoint[6]), 
            .I3(n4743), .O(n72371));
    defparam n9971_bdd_4_lut_55190.LUT_INIT = 16'he4aa;
    SB_CARRY add_4527_7 (.CI(n54394), .I0(n12545[4]), .I1(n442_adj_4521), 
            .CO(n54395));
    SB_LUT4 n72371_bdd_4_lut (.I0(n72371), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4743), .O(n72374));
    defparam n72371_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9971_bdd_4_lut_55185 (.I0(n9971), .I1(n68489), .I2(setpoint[5]), 
            .I3(n4743), .O(n72365));
    defparam n9971_bdd_4_lut_55185.LUT_INIT = 16'he4aa;
    SB_LUT4 n72365_bdd_4_lut (.I0(n72365), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4743), .O(n72368));
    defparam n72365_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54366_3_lut (.I0(n71493), .I1(n290), .I2(n39), .I3(GND_net), 
            .O(n71456));   // verilog/motorControl.v(58[23:46])
    defparam i54366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52100_4_lut (.I0(n43_adj_4525), .I1(n41_adj_4522), .I2(n39), 
            .I3(n71380), .O(n69190));
    defparam i52100_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54233_4_lut (.I0(n69664), .I1(n70778), .I2(n45_adj_4524), 
            .I3(n69184), .O(n71323));   // verilog/motorControl.v(58[23:46])
    defparam i54233_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9971_bdd_4_lut_55180 (.I0(n9971), .I1(n68486), .I2(setpoint[4]), 
            .I3(n4743), .O(n72359));
    defparam n9971_bdd_4_lut_55180.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_30_i9_2_lut (.I0(PWMLimit[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4551));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4552));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4553));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4554));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i21_2_lut (.I0(PWMLimit[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4555));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4556));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4557));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(deadband[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4558));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4559));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4560));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n72359_bdd_4_lut (.I0(n72359), .I1(n535[4]), .I2(n455[4]), 
            .I3(n4743), .O(n72362));
    defparam n72359_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4527_6_lut (.I0(GND_net), .I1(n12545[3]), .I2(n369), .I3(n54393), 
            .O(n10937[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(deadband[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4561));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4562));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4563));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4564));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4565));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(deadband[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4566));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(deadband[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4567));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(deadband[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4568));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i33_2_lut (.I0(deadband[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4569));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4445));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n455[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4465));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4468));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4467));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4466));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4462));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4463));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4464));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n29864), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n29863), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n29862), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n29861), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n29860), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n29859), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n29858), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n29857), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n29856), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n29855), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n29854), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n29853), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n29852), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n29851), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n29850), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n29849), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n29848), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n29847), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n29846), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n29845), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n29844), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n29843), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n29839), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4527_6 (.CI(n54393), .I0(n12545[3]), .I1(n369), .CO(n54394));
    SB_LUT4 add_4527_5_lut (.I0(GND_net), .I1(n12545[2]), .I2(n296), .I3(n54392), 
            .O(n10937[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_5 (.CI(n54392), .I0(n12545[2]), .I1(n296), .CO(n54393));
    SB_DFFSR counter_2045_2046__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 i52582_3_lut (.I0(n71456), .I1(n285[20]), .I2(n41_adj_4522), 
            .I3(GND_net), .O(n69672));   // verilog/motorControl.v(58[23:46])
    defparam i52582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54235_4_lut (.I0(n69672), .I1(n71323), .I2(n45_adj_4524), 
            .I3(n69190), .O(n71325));   // verilog/motorControl.v(58[23:46])
    defparam i54235_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54236_3_lut (.I0(n71325), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i54236_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29097), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_5139_11_lut (.I0(GND_net), .I1(n20115[8]), .I2(n770), 
            .I3(n54009), .O(n19898[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51491_2_lut (.I0(PWMLimit[9]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68266));
    defparam i51491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51516_2_lut (.I0(PWMLimit[13]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68252));
    defparam i51516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9971_bdd_4_lut_54862 (.I0(n9971), .I1(n68368), .I2(setpoint[11]), 
            .I3(n4743), .O(n71969));
    defparam n9971_bdd_4_lut_54862.LUT_INIT = 16'he4aa;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n53803), .I0(GND_net), .I1(n1_adj_5001[11]), 
            .CO(n53804));
    SB_LUT4 add_4527_4_lut (.I0(GND_net), .I1(n12545[1]), .I2(n223_adj_4571), 
            .I3(n54391), .O(n10937[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_10_lut (.I0(GND_net), .I1(n20115[7]), .I2(n697), 
            .I3(n54008), .O(n19898[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51524_2_lut (.I0(PWMLimit[14]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68271));
    defparam i51524_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52102_2_lut (.I0(PWMLimit[15]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68284));
    defparam i52102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n348));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51648_2_lut (.I0(PWMLimit[10]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68343));
    defparam i51648_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4527_4 (.CI(n54391), .I0(n12545[1]), .I1(n223_adj_4571), 
            .CO(n54392));
    SB_LUT4 i51582_2_lut (.I0(PWMLimit[16]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68296));
    defparam i51582_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4527_3_lut (.I0(GND_net), .I1(n12545[0]), .I2(n150), .I3(n54390), 
            .O(n10937[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_3 (.CI(n54390), .I0(n12545[0]), .I1(n150), .CO(n54391));
    SB_LUT4 add_4527_2_lut (.I0(GND_net), .I1(n8_adj_4572), .I2(n77), 
            .I3(GND_net), .O(n10937[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n11420[21]), .I2(GND_net), 
            .I3(n54827), .O(n10961[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n11420[20]), .I2(GND_net), 
            .I3(n54826), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n54826), .I0(n11420[20]), .I1(GND_net), 
            .CO(n54827));
    SB_CARRY add_4527_2 (.CI(GND_net), .I0(n8_adj_4572), .I1(n77), .CO(n54390));
    SB_CARRY add_5139_10 (.CI(n54008), .I0(n20115[7]), .I1(n697), .CO(n54009));
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[10]), 
            .I3(n53802), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_17 (.CI(n53638), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n53639));
    SB_CARRY sub_15_add_2_6 (.CI(n53604), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n53605));
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n53637), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n11420[19]), .I2(GND_net), 
            .I3(n54825), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4744_22_lut (.I0(GND_net), .I1(n13820[19]), .I2(GND_net), 
            .I3(n54389), .O(n12545[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_9_lut (.I0(GND_net), .I1(n20115[6]), .I2(n624), .I3(n54007), 
            .O(n19898[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_12 (.CI(n53802), .I0(GND_net), .I1(n1_adj_5001[10]), 
            .CO(n53803));
    SB_CARRY mult_23_add_1221_22 (.CI(n54825), .I0(n11420[19]), .I1(GND_net), 
            .CO(n54826));
    SB_CARRY add_16_16 (.CI(n53637), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n53638));
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n53636), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n11420[18]), .I2(GND_net), 
            .I3(n54824), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51718_2_lut (.I0(PWMLimit[17]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68372));
    defparam i51718_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_21 (.CI(n54824), .I0(n11420[18]), .I1(GND_net), 
            .CO(n54825));
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n11420[17]), .I2(GND_net), 
            .I3(n54823), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4574));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_20 (.CI(n54823), .I0(n11420[17]), .I1(GND_net), 
            .CO(n54824));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n11420[16]), .I2(GND_net), 
            .I3(n54822), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n54822), .I0(n11420[16]), .I1(GND_net), 
            .CO(n54823));
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n11420[15]), .I2(GND_net), 
            .I3(n54821), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4575));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_18 (.CI(n54821), .I0(n11420[15]), .I1(GND_net), 
            .CO(n54822));
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4576));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4577));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n11420[14]), .I2(GND_net), 
            .I3(n54820), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4578));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_17 (.CI(n54820), .I0(n11420[14]), .I1(GND_net), 
            .CO(n54821));
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4579));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n11420[13]), .I2(n1096_adj_4580), 
            .I3(n54819), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n54819), .I0(n11420[13]), .I1(n1096_adj_4580), 
            .CO(n54820));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n11420[12]), .I2(n1023_adj_4581), 
            .I3(n54818), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4582));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_15 (.CI(n54818), .I0(n11420[12]), .I1(n1023_adj_4581), 
            .CO(n54819));
    SB_LUT4 add_4744_21_lut (.I0(GND_net), .I1(n13820[18]), .I2(GND_net), 
            .I3(n54388), .O(n12545[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n11420[11]), .I2(n950_adj_4583), 
            .I3(n54817), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_21 (.CI(n54388), .I0(n13820[18]), .I1(GND_net), 
            .CO(n54389));
    SB_CARRY add_5139_9 (.CI(n54007), .I0(n20115[6]), .I1(n624), .CO(n54008));
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4584));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_14 (.CI(n54817), .I0(n11420[11]), .I1(n950_adj_4583), 
            .CO(n54818));
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n11420[10]), .I2(n877_adj_4585), 
            .I3(n54816), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_13 (.CI(n54816), .I0(n11420[10]), .I1(n877_adj_4585), 
            .CO(n54817));
    SB_LUT4 add_4744_20_lut (.I0(GND_net), .I1(n13820[17]), .I2(GND_net), 
            .I3(n54387), .O(n12545[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_20 (.CI(n54387), .I0(n13820[17]), .I1(GND_net), 
            .CO(n54388));
    SB_LUT4 add_5139_8_lut (.I0(GND_net), .I1(n20115[5]), .I2(n551_adj_4586), 
            .I3(n54006), .O(n19898[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n11420[9]), .I2(n804_adj_4587), 
            .I3(n54815), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_12 (.CI(n54815), .I0(n11420[9]), .I1(n804_adj_4587), 
            .CO(n54816));
    SB_LUT4 add_4744_19_lut (.I0(GND_net), .I1(n13820[16]), .I2(GND_net), 
            .I3(n54386), .O(n12545[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_8 (.CI(n54006), .I0(n20115[5]), .I1(n551_adj_4586), 
            .CO(n54007));
    SB_LUT4 add_5139_7_lut (.I0(GND_net), .I1(n20115[4]), .I2(n478_adj_4589), 
            .I3(n54005), .O(n19898[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_19 (.CI(n54386), .I0(n13820[16]), .I1(GND_net), 
            .CO(n54387));
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n11420[8]), .I2(n731_adj_4590), 
            .I3(n54814), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_11 (.CI(n54814), .I0(n11420[8]), .I1(n731_adj_4590), 
            .CO(n54815));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n11420[7]), .I2(n658_adj_4592), 
            .I3(n54813), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_10 (.CI(n54813), .I0(n11420[7]), .I1(n658_adj_4592), 
            .CO(n54814));
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n11420[6]), .I2(n585_adj_4595), 
            .I3(n54812), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n54812), .I0(n11420[6]), .I1(n585_adj_4595), 
            .CO(n54813));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n11420[5]), .I2(n512_adj_4596), 
            .I3(n54811), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_8 (.CI(n54811), .I0(n11420[5]), .I1(n512_adj_4596), 
            .CO(n54812));
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n11420[4]), .I2(n439_adj_4597), 
            .I3(n54810), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4598));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4599));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_7 (.CI(n54810), .I0(n11420[4]), .I1(n439_adj_4597), 
            .CO(n54811));
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n11420[3]), .I2(n366_adj_4600), 
            .I3(n54809), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n54809), .I0(n11420[3]), .I1(n366_adj_4600), 
            .CO(n54810));
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n11420[2]), .I2(n293_adj_4601), 
            .I3(n54808), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_5 (.CI(n54808), .I0(n11420[2]), .I1(n293_adj_4601), 
            .CO(n54809));
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n11420[1]), .I2(n220_adj_4602), 
            .I3(n54807), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_4 (.CI(n54807), .I0(n11420[1]), .I1(n220_adj_4602), 
            .CO(n54808));
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n11420[0]), .I2(n147_adj_4603), 
            .I3(n54806), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_3 (.CI(n54806), .I0(n11420[0]), .I1(n147_adj_4603), 
            .CO(n54807));
    SB_LUT4 add_4744_18_lut (.I0(GND_net), .I1(n13820[15]), .I2(GND_net), 
            .I3(n54385), .O(n12545[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_4604), .I2(n74_adj_4605), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_18 (.CI(n54385), .I0(n13820[15]), .I1(GND_net), 
            .CO(n54386));
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5_adj_4604), .I1(n74_adj_4605), 
            .CO(n54806));
    SB_LUT4 add_4548_23_lut (.I0(GND_net), .I1(n12982[20]), .I2(GND_net), 
            .I3(n54805), .O(n11420[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4548_22_lut (.I0(GND_net), .I1(n12982[19]), .I2(GND_net), 
            .I3(n54804), .O(n11420[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_17_lut (.I0(GND_net), .I1(n13820[14]), .I2(GND_net), 
            .I3(n54384), .O(n12545[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_22 (.CI(n54804), .I0(n12982[19]), .I1(GND_net), 
            .CO(n54805));
    SB_LUT4 add_4548_21_lut (.I0(GND_net), .I1(n12982[18]), .I2(GND_net), 
            .I3(n54803), .O(n11420[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_21 (.CI(n54803), .I0(n12982[18]), .I1(GND_net), 
            .CO(n54804));
    SB_CARRY add_4744_17 (.CI(n54384), .I0(n13820[14]), .I1(GND_net), 
            .CO(n54385));
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51673_2_lut (.I0(PWMLimit[12]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68390));
    defparam i51673_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_20_lut (.I0(GND_net), .I1(n12982[17]), .I2(GND_net), 
            .I3(n54802), .O(n11420[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_16_lut (.I0(GND_net), .I1(n13820[13]), .I2(n1102), 
            .I3(n54383), .O(n12545[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_20 (.CI(n54802), .I0(n12982[17]), .I1(GND_net), 
            .CO(n54803));
    SB_CARRY add_4744_16 (.CI(n54383), .I0(n13820[13]), .I1(n1102), .CO(n54384));
    SB_LUT4 add_4548_19_lut (.I0(GND_net), .I1(n12982[16]), .I2(GND_net), 
            .I3(n54801), .O(n11420[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_19 (.CI(n54801), .I0(n12982[16]), .I1(GND_net), 
            .CO(n54802));
    SB_LUT4 add_4548_18_lut (.I0(GND_net), .I1(n12982[15]), .I2(GND_net), 
            .I3(n54800), .O(n11420[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_15_lut (.I0(GND_net), .I1(n13820[12]), .I2(n1029), 
            .I3(n54382), .O(n12545[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4548_18 (.CI(n54800), .I0(n12982[15]), .I1(GND_net), 
            .CO(n54801));
    SB_LUT4 add_4548_17_lut (.I0(GND_net), .I1(n12982[14]), .I2(GND_net), 
            .I3(n54799), .O(n11420[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_17 (.CI(n54799), .I0(n12982[14]), .I1(GND_net), 
            .CO(n54800));
    SB_CARRY add_4744_15 (.CI(n54382), .I0(n13820[12]), .I1(n1029), .CO(n54383));
    SB_LUT4 add_4548_16_lut (.I0(GND_net), .I1(n12982[13]), .I2(n1099_adj_4606), 
            .I3(n54798), .O(n11420[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_14_lut (.I0(GND_net), .I1(n13820[11]), .I2(n956), 
            .I3(n54381), .O(n12545[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_14 (.CI(n54381), .I0(n13820[11]), .I1(n956), .CO(n54382));
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4744_13_lut (.I0(GND_net), .I1(n13820[10]), .I2(n883), 
            .I3(n54380), .O(n12545[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_16 (.CI(n54798), .I0(n12982[13]), .I1(n1099_adj_4606), 
            .CO(n54799));
    SB_CARRY add_4744_13 (.CI(n54380), .I0(n13820[10]), .I1(n883), .CO(n54381));
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_15_lut (.I0(GND_net), .I1(n12982[12]), .I2(n1026_adj_4607), 
            .I3(n54797), .O(n11420[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_12_lut (.I0(GND_net), .I1(n13820[9]), .I2(n810), 
            .I3(n54379), .O(n12545[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_15 (.CI(n54797), .I0(n12982[12]), .I1(n1026_adj_4607), 
            .CO(n54798));
    SB_CARRY add_4744_12 (.CI(n54379), .I0(n13820[9]), .I1(n810), .CO(n54380));
    SB_LUT4 add_4548_14_lut (.I0(GND_net), .I1(n12982[11]), .I2(n953_adj_4608), 
            .I3(n54796), .O(n11420[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_11_lut (.I0(GND_net), .I1(n13820[8]), .I2(n737), 
            .I3(n54378), .O(n12545[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_14 (.CI(n54796), .I0(n12982[11]), .I1(n953_adj_4608), 
            .CO(n54797));
    SB_CARRY add_4744_11 (.CI(n54378), .I0(n13820[8]), .I1(n737), .CO(n54379));
    SB_LUT4 add_4548_13_lut (.I0(GND_net), .I1(n12982[10]), .I2(n880_adj_4609), 
            .I3(n54795), .O(n11420[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_13 (.CI(n54795), .I0(n12982[10]), .I1(n880_adj_4609), 
            .CO(n54796));
    SB_LUT4 add_4744_10_lut (.I0(GND_net), .I1(n13820[7]), .I2(n664), 
            .I3(n54377), .O(n12545[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4548_12_lut (.I0(GND_net), .I1(n12982[9]), .I2(n807_adj_4610), 
            .I3(n54794), .O(n11420[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_12 (.CI(n54794), .I0(n12982[9]), .I1(n807_adj_4610), 
            .CO(n54795));
    SB_LUT4 add_4548_11_lut (.I0(GND_net), .I1(n12982[8]), .I2(n734_adj_4611), 
            .I3(n54793), .O(n11420[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4548_11 (.CI(n54793), .I0(n12982[8]), .I1(n734_adj_4611), 
            .CO(n54794));
    SB_CARRY add_4744_10 (.CI(n54377), .I0(n13820[7]), .I1(n664), .CO(n54378));
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_10_lut (.I0(GND_net), .I1(n12982[7]), .I2(n661_adj_4612), 
            .I3(n54792), .O(n11420[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_9_lut (.I0(GND_net), .I1(n13820[6]), .I2(n591), .I3(n54376), 
            .O(n12545[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_10 (.CI(n54792), .I0(n12982[7]), .I1(n661_adj_4612), 
            .CO(n54793));
    SB_LUT4 add_4548_9_lut (.I0(GND_net), .I1(n12982[6]), .I2(n588_adj_4613), 
            .I3(n54791), .O(n11420[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_9 (.CI(n54791), .I0(n12982[6]), .I1(n588_adj_4613), 
            .CO(n54792));
    SB_LUT4 add_4548_8_lut (.I0(GND_net), .I1(n12982[5]), .I2(n515_adj_4614), 
            .I3(n54790), .O(n11420[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_9 (.CI(n54376), .I0(n13820[6]), .I1(n591), .CO(n54377));
    SB_LUT4 add_4744_8_lut (.I0(GND_net), .I1(n13820[5]), .I2(n518), .I3(n54375), 
            .O(n12545[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_8 (.CI(n54790), .I0(n12982[5]), .I1(n515_adj_4614), 
            .CO(n54791));
    SB_CARRY add_4744_8 (.CI(n54375), .I0(n13820[5]), .I1(n518), .CO(n54376));
    SB_LUT4 add_4548_7_lut (.I0(GND_net), .I1(n12982[4]), .I2(n442_adj_4615), 
            .I3(n54789), .O(n11420[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_7 (.CI(n54789), .I0(n12982[4]), .I1(n442_adj_4615), 
            .CO(n54790));
    SB_LUT4 add_4744_7_lut (.I0(GND_net), .I1(n13820[4]), .I2(n445_adj_4616), 
            .I3(n54374), .O(n12545[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4617));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_6_lut (.I0(GND_net), .I1(n12982[3]), .I2(n369_adj_4618), 
            .I3(n54788), .O(n11420[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_7 (.CI(n54374), .I0(n13820[4]), .I1(n445_adj_4616), 
            .CO(n54375));
    SB_CARRY add_4548_6 (.CI(n54788), .I0(n12982[3]), .I1(n369_adj_4618), 
            .CO(n54789));
    SB_LUT4 add_4744_6_lut (.I0(GND_net), .I1(n13820[3]), .I2(n372), .I3(n54373), 
            .O(n12545[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_6 (.CI(n54373), .I0(n13820[3]), .I1(n372), .CO(n54374));
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_5_lut (.I0(GND_net), .I1(n12982[2]), .I2(n296_adj_4619), 
            .I3(n54787), .O(n11420[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_5_lut (.I0(GND_net), .I1(n13820[2]), .I2(n299_adj_4620), 
            .I3(n54372), .O(n12545[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_5 (.CI(n54787), .I0(n12982[2]), .I1(n296_adj_4619), 
            .CO(n54788));
    SB_LUT4 add_4548_4_lut (.I0(GND_net), .I1(n12982[1]), .I2(n223_adj_4621), 
            .I3(n54786), .O(n11420[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[9]), 
            .I3(n53801), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_5 (.CI(n54372), .I0(n13820[2]), .I1(n299_adj_4620), 
            .CO(n54373));
    SB_CARRY add_4548_4 (.CI(n54786), .I0(n12982[1]), .I1(n223_adj_4621), 
            .CO(n54787));
    SB_LUT4 add_4744_4_lut (.I0(GND_net), .I1(n13820[1]), .I2(n226_adj_4623), 
            .I3(n54371), .O(n12545[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4548_3_lut (.I0(GND_net), .I1(n12982[0]), .I2(n150_adj_4624), 
            .I3(n54785), .O(n11420[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_4 (.CI(n54371), .I0(n13820[1]), .I1(n226_adj_4623), 
            .CO(n54372));
    SB_CARRY add_4548_3 (.CI(n54785), .I0(n12982[0]), .I1(n150_adj_4624), 
            .CO(n54786));
    SB_CARRY add_16_15 (.CI(n53636), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n53637));
    SB_LUT4 add_4744_3_lut (.I0(GND_net), .I1(n13820[0]), .I2(n153), .I3(n54370), 
            .O(n12545[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4625));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4548_2_lut (.I0(GND_net), .I1(n8_adj_4626), .I2(n77_adj_4627), 
            .I3(GND_net), .O(n11420[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4548_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4548_2 (.CI(GND_net), .I0(n8_adj_4626), .I1(n77_adj_4627), 
            .CO(n54785));
    SB_LUT4 add_4763_22_lut (.I0(GND_net), .I1(n14216[19]), .I2(GND_net), 
            .I3(n54784), .O(n12982[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_3 (.CI(n54370), .I0(n13820[0]), .I1(n153), .CO(n54371));
    SB_LUT4 add_4763_21_lut (.I0(GND_net), .I1(n14216[18]), .I2(GND_net), 
            .I3(n54783), .O(n12982[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4744_2_lut (.I0(GND_net), .I1(n11_adj_4628), .I2(n80), 
            .I3(GND_net), .O(n12545[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4744_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4744_2 (.CI(GND_net), .I0(n11_adj_4628), .I1(n80), .CO(n54370));
    SB_CARRY add_4763_21 (.CI(n54783), .I0(n14216[18]), .I1(GND_net), 
            .CO(n54784));
    SB_LUT4 add_4800_21_lut (.I0(GND_net), .I1(n14929[18]), .I2(GND_net), 
            .I3(n54369), .O(n13820[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_20_lut (.I0(GND_net), .I1(n14216[17]), .I2(GND_net), 
            .I3(n54782), .O(n12982[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_20_lut (.I0(GND_net), .I1(n14929[17]), .I2(GND_net), 
            .I3(n54368), .O(n13820[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_20 (.CI(n54368), .I0(n14929[17]), .I1(GND_net), 
            .CO(n54369));
    SB_CARRY add_4763_20 (.CI(n54782), .I0(n14216[17]), .I1(GND_net), 
            .CO(n54783));
    SB_LUT4 add_4763_19_lut (.I0(GND_net), .I1(n14216[16]), .I2(GND_net), 
            .I3(n54781), .O(n12982[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_19_lut (.I0(GND_net), .I1(n14929[16]), .I2(GND_net), 
            .I3(n54367), .O(n13820[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_19 (.CI(n54367), .I0(n14929[16]), .I1(GND_net), 
            .CO(n54368));
    SB_CARRY add_4763_19 (.CI(n54781), .I0(n14216[16]), .I1(GND_net), 
            .CO(n54782));
    SB_LUT4 add_4800_18_lut (.I0(GND_net), .I1(n14929[15]), .I2(GND_net), 
            .I3(n54366), .O(n13820[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_18 (.CI(n54366), .I0(n14929[15]), .I1(GND_net), 
            .CO(n54367));
    SB_CARRY unary_minus_33_add_3_11 (.CI(n53801), .I0(GND_net), .I1(n1_adj_5001[9]), 
            .CO(n53802));
    SB_LUT4 add_4763_18_lut (.I0(GND_net), .I1(n14216[15]), .I2(GND_net), 
            .I3(n54780), .O(n12982[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_17_lut (.I0(GND_net), .I1(n14929[14]), .I2(GND_net), 
            .I3(n54365), .O(n13820[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_17 (.CI(n54365), .I0(n14929[14]), .I1(GND_net), 
            .CO(n54366));
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4763_18 (.CI(n54780), .I0(n14216[15]), .I1(GND_net), 
            .CO(n54781));
    SB_LUT4 add_4800_16_lut (.I0(GND_net), .I1(n14929[13]), .I2(n1105), 
            .I3(n54364), .O(n13820[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_17_lut (.I0(GND_net), .I1(n14216[14]), .I2(GND_net), 
            .I3(n54779), .O(n12982[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_16 (.CI(n54364), .I0(n14929[13]), .I1(n1105), .CO(n54365));
    SB_CARRY add_4763_17 (.CI(n54779), .I0(n14216[14]), .I1(GND_net), 
            .CO(n54780));
    SB_LUT4 add_4763_16_lut (.I0(GND_net), .I1(n14216[13]), .I2(n1102_adj_4629), 
            .I3(n54778), .O(n12982[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_15_lut (.I0(GND_net), .I1(n14929[12]), .I2(n1032), 
            .I3(n54363), .O(n13820[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_16 (.CI(n54778), .I0(n14216[13]), .I1(n1102_adj_4629), 
            .CO(n54779));
    SB_CARRY add_4800_15 (.CI(n54363), .I0(n14929[12]), .I1(n1032), .CO(n54364));
    SB_LUT4 add_4763_15_lut (.I0(GND_net), .I1(n14216[12]), .I2(n1029_adj_4630), 
            .I3(n54777), .O(n12982[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_14_lut (.I0(GND_net), .I1(n14929[11]), .I2(n959), 
            .I3(n54362), .O(n13820[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_15 (.CI(n54777), .I0(n14216[12]), .I1(n1029_adj_4630), 
            .CO(n54778));
    SB_CARRY add_4800_14 (.CI(n54362), .I0(n14929[11]), .I1(n959), .CO(n54363));
    SB_LUT4 add_4800_13_lut (.I0(GND_net), .I1(n14929[10]), .I2(n886), 
            .I3(n54361), .O(n13820[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_14_lut (.I0(GND_net), .I1(n14216[11]), .I2(n956_adj_4631), 
            .I3(n54776), .O(n12982[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_13 (.CI(n54361), .I0(n14929[10]), .I1(n886), .CO(n54362));
    SB_CARRY add_4763_14 (.CI(n54776), .I0(n14216[11]), .I1(n956_adj_4631), 
            .CO(n54777));
    SB_LUT4 add_4800_12_lut (.I0(GND_net), .I1(n14929[9]), .I2(n813), 
            .I3(n54360), .O(n13820[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_13_lut (.I0(GND_net), .I1(n14216[10]), .I2(n883_adj_4632), 
            .I3(n54775), .O(n12982[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_12 (.CI(n54360), .I0(n14929[9]), .I1(n813), .CO(n54361));
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n346));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4763_13 (.CI(n54775), .I0(n14216[10]), .I1(n883_adj_4632), 
            .CO(n54776));
    SB_LUT4 add_4800_11_lut (.I0(GND_net), .I1(n14929[8]), .I2(n740), 
            .I3(n54359), .O(n13820[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_12_lut (.I0(GND_net), .I1(n14216[9]), .I2(n810_adj_4633), 
            .I3(n54774), .O(n12982[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i75_2_lut (.I0(\Ki[1] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i75_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4800_11 (.CI(n54359), .I0(n14929[8]), .I1(n740), .CO(n54360));
    SB_CARRY add_4763_12 (.CI(n54774), .I0(n14216[9]), .I1(n810_adj_4633), 
            .CO(n54775));
    SB_LUT4 add_4800_10_lut (.I0(GND_net), .I1(n14929[7]), .I2(n667), 
            .I3(n54358), .O(n13820[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_11_lut (.I0(GND_net), .I1(n14216[8]), .I2(n737_adj_4634), 
            .I3(n54773), .O(n12982[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_10 (.CI(n54358), .I0(n14929[7]), .I1(n667), .CO(n54359));
    SB_CARRY add_4763_11 (.CI(n54773), .I0(n14216[8]), .I1(n737_adj_4634), 
            .CO(n54774));
    SB_LUT4 add_4800_9_lut (.I0(GND_net), .I1(n14929[6]), .I2(n594), .I3(n54357), 
            .O(n13820[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_9 (.CI(n54357), .I0(n14929[6]), .I1(n594), .CO(n54358));
    SB_LUT4 add_4763_10_lut (.I0(GND_net), .I1(n14216[7]), .I2(n664_adj_4635), 
            .I3(n54772), .O(n12982[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_8_lut (.I0(GND_net), .I1(n14929[5]), .I2(n521), .I3(n54356), 
            .O(n13820[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_10 (.CI(n54772), .I0(n14216[7]), .I1(n664_adj_4635), 
            .CO(n54773));
    SB_LUT4 add_4763_9_lut (.I0(GND_net), .I1(n14216[6]), .I2(n591_adj_4636), 
            .I3(n54771), .O(n12982[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_8 (.CI(n54356), .I0(n14929[5]), .I1(n521), .CO(n54357));
    SB_LUT4 add_4800_7_lut (.I0(GND_net), .I1(n14929[4]), .I2(n448_adj_4637), 
            .I3(n54355), .O(n13820[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4800_7 (.CI(n54355), .I0(n14929[4]), .I1(n448_adj_4637), 
            .CO(n54356));
    SB_LUT4 add_4800_6_lut (.I0(GND_net), .I1(n14929[3]), .I2(n375), .I3(n54354), 
            .O(n13820[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_9 (.CI(n54771), .I0(n14216[6]), .I1(n591_adj_4636), 
            .CO(n54772));
    SB_CARRY add_4800_6 (.CI(n54354), .I0(n14929[3]), .I1(n375), .CO(n54355));
    SB_LUT4 add_4763_8_lut (.I0(GND_net), .I1(n14216[5]), .I2(n518_adj_4638), 
            .I3(n54770), .O(n12982[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_5_lut (.I0(GND_net), .I1(n14929[2]), .I2(n302_adj_4639), 
            .I3(n54353), .O(n13820[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_8 (.CI(n54770), .I0(n14216[5]), .I1(n518_adj_4638), 
            .CO(n54771));
    SB_CARRY add_4800_5 (.CI(n54353), .I0(n14929[2]), .I1(n302_adj_4639), 
            .CO(n54354));
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4516));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4763_7_lut (.I0(GND_net), .I1(n14216[4]), .I2(n445_adj_4640), 
            .I3(n54769), .O(n12982[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4763_7 (.CI(n54769), .I0(n14216[4]), .I1(n445_adj_4640), 
            .CO(n54770));
    SB_LUT4 add_4763_6_lut (.I0(GND_net), .I1(n14216[3]), .I2(n372_adj_4641), 
            .I3(n54768), .O(n12982[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_4_lut (.I0(GND_net), .I1(n14929[1]), .I2(n229), .I3(n54352), 
            .O(n13820[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_6 (.CI(n54768), .I0(n14216[3]), .I1(n372_adj_4641), 
            .CO(n54769));
    SB_CARRY add_4800_4 (.CI(n54352), .I0(n14929[1]), .I1(n229), .CO(n54353));
    SB_LUT4 add_4763_5_lut (.I0(GND_net), .I1(n14216[2]), .I2(n299_adj_4642), 
            .I3(n54767), .O(n12982[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_3_lut (.I0(GND_net), .I1(n14929[0]), .I2(n156), .I3(n54351), 
            .O(n13820[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_5 (.CI(n54767), .I0(n14216[2]), .I1(n299_adj_4642), 
            .CO(n54768));
    SB_CARRY add_4800_3 (.CI(n54351), .I0(n14929[0]), .I1(n156), .CO(n54352));
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n349), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4763_4_lut (.I0(GND_net), .I1(n14216[1]), .I2(n226_adj_4643), 
            .I3(n54766), .O(n12982[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4800_2_lut (.I0(GND_net), .I1(n14_adj_4644), .I2(n83), 
            .I3(GND_net), .O(n13820[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4800_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_4 (.CI(n54766), .I0(n14216[1]), .I1(n226_adj_4643), 
            .CO(n54767));
    SB_CARRY add_4800_2 (.CI(GND_net), .I0(n14_adj_4644), .I1(n83), .CO(n54351));
    SB_LUT4 add_5127_12_lut (.I0(GND_net), .I1(n19994[9]), .I2(n840_adj_4645), 
            .I3(n54350), .O(n19754[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4763_3_lut (.I0(GND_net), .I1(n14216[0]), .I2(n153_adj_4646), 
            .I3(n54765), .O(n12982[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_11_lut (.I0(GND_net), .I1(n19994[8]), .I2(n767_adj_4647), 
            .I3(n54349), .O(n19754[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4763_3 (.CI(n54765), .I0(n14216[0]), .I1(n153_adj_4646), 
            .CO(n54766));
    SB_CARRY add_5127_11 (.CI(n54349), .I0(n19994[8]), .I1(n767_adj_4647), 
            .CO(n54350));
    SB_LUT4 add_5127_10_lut (.I0(GND_net), .I1(n19994[7]), .I2(n694_adj_4648), 
            .I3(n54348), .O(n19754[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4763_2_lut (.I0(GND_net), .I1(n11_adj_4649), .I2(n80_adj_4650), 
            .I3(GND_net), .O(n12982[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4763_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5127_10 (.CI(n54348), .I0(n19994[7]), .I1(n694_adj_4648), 
            .CO(n54349));
    SB_CARRY add_4763_2 (.CI(GND_net), .I0(n11_adj_4649), .I1(n80_adj_4650), 
            .CO(n54765));
    SB_LUT4 add_5127_9_lut (.I0(GND_net), .I1(n19994[6]), .I2(n621_adj_4651), 
            .I3(n54347), .O(n19754[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5190_8_lut (.I0(GND_net), .I1(n20542[5]), .I2(n560_adj_4652), 
            .I3(n54764), .O(n20433[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_9 (.CI(n54347), .I0(n19994[6]), .I1(n621_adj_4651), 
            .CO(n54348));
    SB_LUT4 add_5190_7_lut (.I0(GND_net), .I1(n20542[4]), .I2(n487_adj_4653), 
            .I3(n54763), .O(n20433[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_8_lut (.I0(GND_net), .I1(n19994[5]), .I2(n548_adj_4654), 
            .I3(n54346), .O(n19754[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5190_7 (.CI(n54763), .I0(n20542[4]), .I1(n487_adj_4653), 
            .CO(n54764));
    SB_CARRY add_5127_8 (.CI(n54346), .I0(n19994[5]), .I1(n548_adj_4654), 
            .CO(n54347));
    SB_LUT4 add_5190_6_lut (.I0(GND_net), .I1(n20542[3]), .I2(n414_adj_4655), 
            .I3(n54762), .O(n20433[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_7_lut (.I0(GND_net), .I1(n19994[4]), .I2(n475_adj_4656), 
            .I3(n54345), .O(n19754[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_7 (.CI(n54345), .I0(n19994[4]), .I1(n475_adj_4656), 
            .CO(n54346));
    SB_LUT4 add_5127_6_lut (.I0(GND_net), .I1(n19994[3]), .I2(n402_adj_4657), 
            .I3(n54344), .O(n19754[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[8]), 
            .I3(n53800), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n53635), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_14 (.CI(n53635), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n53636));
    SB_CARRY add_5139_7 (.CI(n54005), .I0(n20115[4]), .I1(n478_adj_4589), 
            .CO(n54006));
    SB_CARRY add_5190_6 (.CI(n54762), .I0(n20542[3]), .I1(n414_adj_4655), 
            .CO(n54763));
    SB_CARRY add_5127_6 (.CI(n54344), .I0(n19994[3]), .I1(n402_adj_4657), 
            .CO(n54345));
    SB_LUT4 add_5127_5_lut (.I0(GND_net), .I1(n19994[2]), .I2(n329_adj_4659), 
            .I3(n54343), .O(n19754[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5190_5_lut (.I0(GND_net), .I1(n20542[2]), .I2(n341_adj_4660), 
            .I3(n54761), .O(n20433[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5190_5 (.CI(n54761), .I0(n20542[2]), .I1(n341_adj_4660), 
            .CO(n54762));
    SB_CARRY add_5127_5 (.CI(n54343), .I0(n19994[2]), .I1(n329_adj_4659), 
            .CO(n54344));
    SB_LUT4 add_5127_4_lut (.I0(GND_net), .I1(n19994[1]), .I2(n256_adj_4661), 
            .I3(n54342), .O(n19754[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_4 (.CI(n54342), .I0(n19994[1]), .I1(n256_adj_4661), 
            .CO(n54343));
    SB_CARRY unary_minus_33_add_3_10 (.CI(n53800), .I0(GND_net), .I1(n1_adj_5001[8]), 
            .CO(n53801));
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4662));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5127_3_lut (.I0(GND_net), .I1(n19994[0]), .I2(n183_adj_4663), 
            .I3(n54341), .O(n19754[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5127_3 (.CI(n54341), .I0(n19994[0]), .I1(n183_adj_4663), 
            .CO(n54342));
    SB_LUT4 add_5190_4_lut (.I0(GND_net), .I1(n20542[1]), .I2(n268_adj_4664), 
            .I3(n54760), .O(n20433[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5127_2_lut (.I0(GND_net), .I1(n41_adj_4665), .I2(n110_adj_4666), 
            .I3(GND_net), .O(n19754[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5127_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5190_4 (.CI(n54760), .I0(n20542[1]), .I1(n268_adj_4664), 
            .CO(n54761));
    SB_CARRY add_5127_2 (.CI(GND_net), .I0(n41_adj_4665), .I1(n110_adj_4666), 
            .CO(n54341));
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4668));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5190_3_lut (.I0(GND_net), .I1(n20542[0]), .I2(n195_adj_4669), 
            .I3(n54759), .O(n20433[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n358));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5190_3 (.CI(n54759), .I0(n20542[0]), .I1(n195_adj_4669), 
            .CO(n54760));
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5190_2_lut (.I0(GND_net), .I1(n53_adj_4671), .I2(n122_adj_4672), 
            .I3(GND_net), .O(n20433[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5190_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_6_lut (.I0(GND_net), .I1(n20115[3]), .I2(n405), .I3(n54004), 
            .O(n19898[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5190_2 (.CI(GND_net), .I0(n53_adj_4671), .I1(n122_adj_4672), 
            .CO(n54759));
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n53634), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_6 (.CI(n54004), .I0(n20115[3]), .I1(n405), .CO(n54005));
    SB_CARRY add_16_13 (.CI(n53634), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n53635));
    SB_LUT4 add_5139_5_lut (.I0(GND_net), .I1(n20115[2]), .I2(n332_adj_4673), 
            .I3(n54003), .O(n19898[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_21_lut (.I0(GND_net), .I1(n15286[18]), .I2(GND_net), 
            .I3(n54758), .O(n14216[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_20_lut (.I0(GND_net), .I1(n15286[17]), .I2(GND_net), 
            .I3(n54757), .O(n14216[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_20 (.CI(n54757), .I0(n15286[17]), .I1(GND_net), 
            .CO(n54758));
    SB_LUT4 add_4818_19_lut (.I0(GND_net), .I1(n15286[16]), .I2(GND_net), 
            .I3(n54756), .O(n14216[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_5 (.CI(n54003), .I0(n20115[2]), .I1(n332_adj_4673), 
            .CO(n54004));
    SB_CARRY add_4818_19 (.CI(n54756), .I0(n15286[16]), .I1(GND_net), 
            .CO(n54757));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[7]), 
            .I3(n53799), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4674));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_18_lut (.I0(GND_net), .I1(n15286[15]), .I2(GND_net), 
            .I3(n54755), .O(n14216[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_4_lut (.I0(GND_net), .I1(n20115[1]), .I2(n259), .I3(n54002), 
            .O(n19898[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_18 (.CI(n54755), .I0(n15286[15]), .I1(GND_net), 
            .CO(n54756));
    SB_CARRY add_5139_4 (.CI(n54002), .I0(n20115[1]), .I1(n259), .CO(n54003));
    SB_LUT4 add_5139_3_lut (.I0(GND_net), .I1(n20115[0]), .I2(n186), .I3(n54001), 
            .O(n19898[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_17_lut (.I0(GND_net), .I1(n15286[14]), .I2(GND_net), 
            .I3(n54754), .O(n14216[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_3 (.CI(n54001), .I0(n20115[0]), .I1(n186), .CO(n54002));
    SB_CARRY add_4818_17 (.CI(n54754), .I0(n15286[14]), .I1(GND_net), 
            .CO(n54755));
    SB_LUT4 add_5139_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19898[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_16_lut (.I0(GND_net), .I1(n15286[13]), .I2(n1105_adj_4675), 
            .I3(n54753), .O(n14216[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n54001));
    SB_CARRY add_4818_16 (.CI(n54753), .I0(n15286[13]), .I1(n1105_adj_4675), 
            .CO(n54754));
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n358), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4515));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_15_lut (.I0(GND_net), .I1(n15286[12]), .I2(n1032_adj_4676), 
            .I3(n54752), .O(n14216[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4818_15 (.CI(n54752), .I0(n15286[12]), .I1(n1032_adj_4676), 
            .CO(n54753));
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_14_lut (.I0(GND_net), .I1(n15286[11]), .I2(n959_adj_4677), 
            .I3(n54751), .O(n14216[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_14 (.CI(n54751), .I0(n15286[11]), .I1(n959_adj_4677), 
            .CO(n54752));
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_13_lut (.I0(GND_net), .I1(n15286[10]), .I2(n886_adj_4678), 
            .I3(n54750), .O(n14216[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_13 (.CI(n54750), .I0(n15286[10]), .I1(n886_adj_4678), 
            .CO(n54751));
    SB_LUT4 add_4818_12_lut (.I0(GND_net), .I1(n15286[9]), .I2(n813_adj_4679), 
            .I3(n54749), .O(n14216[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n53799), .I0(GND_net), .I1(n1_adj_5001[7]), 
            .CO(n53800));
    SB_CARRY add_4818_12 (.CI(n54749), .I0(n15286[9]), .I1(n813_adj_4679), 
            .CO(n54750));
    SB_LUT4 add_4818_11_lut (.I0(GND_net), .I1(n15286[8]), .I2(n740_adj_4680), 
            .I3(n54748), .O(n14216[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_11 (.CI(n54748), .I0(n15286[8]), .I1(n740_adj_4680), 
            .CO(n54749));
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[6]), 
            .I3(n53798), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_10_lut (.I0(GND_net), .I1(n15286[7]), .I2(n667_adj_4682), 
            .I3(n54747), .O(n14216[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_10 (.CI(n54747), .I0(n15286[7]), .I1(n667_adj_4682), 
            .CO(n54748));
    SB_LUT4 add_4850_20_lut (.I0(GND_net), .I1(n15902[17]), .I2(GND_net), 
            .I3(n54317), .O(n14929[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_19_lut (.I0(GND_net), .I1(n15902[16]), .I2(GND_net), 
            .I3(n54316), .O(n14929[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n350), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4683));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4850_19 (.CI(n54316), .I0(n15902[16]), .I1(GND_net), 
            .CO(n54317));
    SB_CARRY unary_minus_33_add_3_8 (.CI(n53798), .I0(GND_net), .I1(n1_adj_5001[6]), 
            .CO(n53799));
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4684));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4685));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4686));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_9_lut (.I0(GND_net), .I1(n15286[6]), .I2(n594_adj_4687), 
            .I3(n54746), .O(n14216[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4688));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4689));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4818_9 (.CI(n54746), .I0(n15286[6]), .I1(n594_adj_4687), 
            .CO(n54747));
    SB_LUT4 add_4850_18_lut (.I0(GND_net), .I1(n15902[15]), .I2(GND_net), 
            .I3(n54315), .O(n14929[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_18 (.CI(n54315), .I0(n15902[15]), .I1(GND_net), 
            .CO(n54316));
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4818_8_lut (.I0(GND_net), .I1(n15286[5]), .I2(n521_adj_4690), 
            .I3(n54745), .O(n14216[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_17_lut (.I0(GND_net), .I1(n15902[14]), .I2(GND_net), 
            .I3(n54314), .O(n14929[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_17 (.CI(n54314), .I0(n15902[14]), .I1(GND_net), 
            .CO(n54315));
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[5]), 
            .I3(n53797), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4850_16_lut (.I0(GND_net), .I1(n15902[13]), .I2(n1108), 
            .I3(n54313), .O(n14929[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_16 (.CI(n54313), .I0(n15902[13]), .I1(n1108), .CO(n54314));
    SB_CARRY add_4818_8 (.CI(n54745), .I0(n15286[5]), .I1(n521_adj_4690), 
            .CO(n54746));
    SB_LUT4 add_4850_15_lut (.I0(GND_net), .I1(n15902[12]), .I2(n1035), 
            .I3(n54312), .O(n14929[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_15 (.CI(n54312), .I0(n15902[12]), .I1(n1035), .CO(n54313));
    SB_LUT4 add_4818_7_lut (.I0(GND_net), .I1(n15286[4]), .I2(n448_adj_4691), 
            .I3(n54744), .O(n14216[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_14_lut (.I0(GND_net), .I1(n15902[11]), .I2(n962), 
            .I3(n54311), .O(n14929[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4818_7 (.CI(n54744), .I0(n15286[4]), .I1(n448_adj_4691), 
            .CO(n54745));
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4850_14 (.CI(n54311), .I0(n15902[11]), .I1(n962), .CO(n54312));
    SB_LUT4 add_4818_6_lut (.I0(GND_net), .I1(n15286[3]), .I2(n375_adj_4692), 
            .I3(n54743), .O(n14216[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4818_6 (.CI(n54743), .I0(n15286[3]), .I1(n375_adj_4692), 
            .CO(n54744));
    SB_LUT4 add_4850_13_lut (.I0(GND_net), .I1(n15902[10]), .I2(n889), 
            .I3(n54310), .O(n14929[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_13 (.CI(n54310), .I0(n15902[10]), .I1(n889), .CO(n54311));
    SB_LUT4 add_4818_5_lut (.I0(GND_net), .I1(n15286[2]), .I2(n302_adj_4693), 
            .I3(n54742), .O(n14216[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4818_5 (.CI(n54742), .I0(n15286[2]), .I1(n302_adj_4693), 
            .CO(n54743));
    SB_LUT4 add_4850_12_lut (.I0(GND_net), .I1(n15902[9]), .I2(n816), 
            .I3(n54309), .O(n14929[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_12 (.CI(n54309), .I0(n15902[9]), .I1(n816), .CO(n54310));
    SB_LUT4 add_4818_4_lut (.I0(GND_net), .I1(n15286[1]), .I2(n229_adj_4694), 
            .I3(n54741), .O(n14216[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_11_lut (.I0(GND_net), .I1(n15902[8]), .I2(n743), 
            .I3(n54308), .O(n14929[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n53797), .I0(GND_net), .I1(n1_adj_5001[5]), 
            .CO(n53798));
    SB_CARRY add_4850_11 (.CI(n54308), .I0(n15902[8]), .I1(n743), .CO(n54309));
    SB_CARRY add_4818_4 (.CI(n54741), .I0(n15286[1]), .I1(n229_adj_4694), 
            .CO(n54742));
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n53633), .O(n233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n34584), 
            .I3(n53796), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_3_lut (.I0(GND_net), .I1(n15286[0]), .I2(n156_adj_4695), 
            .I3(n54740), .O(n14216[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_10_lut (.I0(GND_net), .I1(n15902[7]), .I2(n670), 
            .I3(n54307), .O(n14929[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_10 (.CI(n54307), .I0(n15902[7]), .I1(n670), .CO(n54308));
    SB_CARRY unary_minus_33_add_3_6 (.CI(n53796), .I0(GND_net), .I1(n34584), 
            .CO(n53797));
    SB_CARRY add_4818_3 (.CI(n54740), .I0(n15286[0]), .I1(n156_adj_4695), 
            .CO(n54741));
    SB_LUT4 add_4850_9_lut (.I0(GND_net), .I1(n15902[6]), .I2(n597), .I3(n54306), 
            .O(n14929[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_9 (.CI(n54306), .I0(n15902[6]), .I1(n597), .CO(n54307));
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[3]), 
            .I3(n53795), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4818_2_lut (.I0(GND_net), .I1(n14_adj_4697), .I2(n83_adj_4698), 
            .I3(GND_net), .O(n14216[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4818_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_8_lut (.I0(GND_net), .I1(n15902[5]), .I2(n524), .I3(n54305), 
            .O(n14929[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_8 (.CI(n54305), .I0(n15902[5]), .I1(n524), .CO(n54306));
    SB_CARRY unary_minus_33_add_3_5 (.CI(n53795), .I0(GND_net), .I1(n1_adj_5001[3]), 
            .CO(n53796));
    SB_CARRY add_4818_2 (.CI(GND_net), .I0(n14_adj_4697), .I1(n83_adj_4698), 
            .CO(n54740));
    SB_LUT4 add_4850_7_lut (.I0(GND_net), .I1(n15902[4]), .I2(n451_adj_4699), 
            .I3(n54304), .O(n14929[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_7 (.CI(n54304), .I0(n15902[4]), .I1(n451_adj_4699), 
            .CO(n54305));
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_12 (.CI(n53633), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n53634));
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[2]), 
            .I3(n53794), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_20_lut (.I0(GND_net), .I1(n16222[17]), .I2(GND_net), 
            .I3(n54739), .O(n15286[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4850_6_lut (.I0(GND_net), .I1(n15902[3]), .I2(n378), .I3(n54303), 
            .O(n14929[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_19_lut (.I0(GND_net), .I1(n16222[16]), .I2(GND_net), 
            .I3(n54738), .O(n15286[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_6 (.CI(n54303), .I0(n15902[3]), .I1(n378), .CO(n54304));
    SB_LUT4 add_4850_5_lut (.I0(GND_net), .I1(n15902[2]), .I2(n305_adj_4701), 
            .I3(n54302), .O(n14929[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_4 (.CI(n53794), .I0(GND_net), .I1(n1_adj_5001[2]), 
            .CO(n53795));
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4867_19 (.CI(n54738), .I0(n16222[16]), .I1(GND_net), 
            .CO(n54739));
    SB_CARRY add_4850_5 (.CI(n54302), .I0(n15902[2]), .I1(n305_adj_4701), 
            .CO(n54303));
    SB_LUT4 add_4850_4_lut (.I0(GND_net), .I1(n15902[1]), .I2(n232), .I3(n54301), 
            .O(n14929[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5001[1]), 
            .I3(n53793), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_18_lut (.I0(GND_net), .I1(n16222[15]), .I2(GND_net), 
            .I3(n54737), .O(n15286[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_4 (.CI(n54301), .I0(n15902[1]), .I1(n232), .CO(n54302));
    SB_LUT4 add_4850_3_lut (.I0(GND_net), .I1(n15902[0]), .I2(n159), .I3(n54300), 
            .O(n14929[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_18 (.CI(n54737), .I0(n16222[15]), .I1(GND_net), 
            .CO(n54738));
    SB_CARRY add_4850_3 (.CI(n54300), .I0(n15902[0]), .I1(n159), .CO(n54301));
    SB_LUT4 add_4850_2_lut (.I0(GND_net), .I1(n17_adj_4703), .I2(n86), 
            .I3(GND_net), .O(n14929[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4850_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_17_lut (.I0(GND_net), .I1(n16222[14]), .I2(GND_net), 
            .I3(n54736), .O(n15286[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4850_2 (.CI(GND_net), .I0(n17_adj_4703), .I1(n86), .CO(n54300));
    SB_CARRY add_4867_17 (.CI(n54736), .I0(n16222[14]), .I1(GND_net), 
            .CO(n54737));
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4704));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_16_lut (.I0(GND_net), .I1(n16222[13]), .I2(n1108_adj_4705), 
            .I3(n54735), .O(n15286[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_16 (.CI(n54735), .I0(n16222[13]), .I1(n1108_adj_4705), 
            .CO(n54736));
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_15_lut (.I0(GND_net), .I1(n16222[12]), .I2(n1035_adj_4706), 
            .I3(n54734), .O(n15286[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_15 (.CI(n54734), .I0(n16222[12]), .I1(n1035_adj_4706), 
            .CO(n54735));
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_14_lut (.I0(GND_net), .I1(n16222[11]), .I2(n962_adj_4707), 
            .I3(n54733), .O(n15286[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_14 (.CI(n54733), .I0(n16222[11]), .I1(n962_adj_4707), 
            .CO(n54734));
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_13_lut (.I0(GND_net), .I1(n16222[10]), .I2(n889_adj_4708), 
            .I3(n54732), .O(n15286[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_13 (.CI(n54732), .I0(n16222[10]), .I1(n889_adj_4708), 
            .CO(n54733));
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n351), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_12_lut (.I0(GND_net), .I1(n16222[9]), .I2(n816_adj_4709), 
            .I3(n54731), .O(n15286[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_12 (.CI(n54731), .I0(n16222[9]), .I1(n816_adj_4709), 
            .CO(n54732));
    SB_LUT4 add_5207_7_lut (.I0(GND_net), .I1(n62402), .I2(n490), .I3(n53977), 
            .O(n20574[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_11_lut (.I0(GND_net), .I1(n16222[8]), .I2(n743_adj_4710), 
            .I3(n54730), .O(n15286[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5207_6_lut (.I0(GND_net), .I1(n20644[3]), .I2(n417), .I3(n53976), 
            .O(n20574[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4711));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5207_6 (.CI(n53976), .I0(n20644[3]), .I1(n417), .CO(n53977));
    SB_CARRY add_4867_11 (.CI(n54730), .I0(n16222[8]), .I1(n743_adj_4710), 
            .CO(n54731));
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4712));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4713));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_10_lut (.I0(GND_net), .I1(n16222[7]), .I2(n670_adj_4714), 
            .I3(n54729), .O(n15286[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5207_5_lut (.I0(GND_net), .I1(n20644[2]), .I2(n344_adj_4715), 
            .I3(n53975), .O(n20574[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4716));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4867_10 (.CI(n54729), .I0(n16222[7]), .I1(n670_adj_4714), 
            .CO(n54730));
    SB_CARRY add_5207_5 (.CI(n53975), .I0(n20644[2]), .I1(n344_adj_4715), 
            .CO(n53976));
    SB_LUT4 add_5207_4_lut (.I0(GND_net), .I1(n20644[1]), .I2(n271), .I3(n53974), 
            .O(n20574[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_9_lut (.I0(GND_net), .I1(n16222[6]), .I2(n597_adj_4717), 
            .I3(n54728), .O(n15286[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_4 (.CI(n53974), .I0(n20644[1]), .I1(n271), .CO(n53975));
    SB_CARRY unary_minus_33_add_3_3 (.CI(n53793), .I0(GND_net), .I1(n1_adj_5001[1]), 
            .CO(n53794));
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n53632), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n53632), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n53633));
    SB_LUT4 add_5207_3_lut (.I0(GND_net), .I1(n20644[0]), .I2(n198), .I3(n53973), 
            .O(n20574[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_3 (.CI(n53973), .I0(n20644[0]), .I1(n198), .CO(n53974));
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n34686), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4867_9 (.CI(n54728), .I0(n16222[6]), .I1(n597_adj_4717), 
            .CO(n54729));
    SB_LUT4 add_5207_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20574[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n53973));
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_8_lut (.I0(GND_net), .I1(n16222[5]), .I2(n524_adj_4718), 
            .I3(n54727), .O(n15286[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_10_lut (.I0(GND_net), .I1(n20292[7]), .I2(n700_adj_4719), 
            .I3(n53972), .O(n20115[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_9_lut (.I0(GND_net), .I1(n20292[6]), .I2(n627_adj_4720), 
            .I3(n53971), .O(n20115[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n34686), 
            .CO(n53793));
    SB_CARRY add_4867_8 (.CI(n54727), .I0(n16222[5]), .I1(n524_adj_4718), 
            .CO(n54728));
    SB_LUT4 add_4867_7_lut (.I0(GND_net), .I1(n16222[4]), .I2(n451_adj_4721), 
            .I3(n54726), .O(n15286[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_9 (.CI(n53971), .I0(n20292[6]), .I1(n627_adj_4720), 
            .CO(n53972));
    SB_LUT4 add_5158_8_lut (.I0(GND_net), .I1(n20292[5]), .I2(n554_adj_4722), 
            .I3(n53970), .O(n20115[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_7 (.CI(n54726), .I0(n16222[4]), .I1(n451_adj_4721), 
            .CO(n54727));
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_5002[23]), 
            .I3(n53792), .O(n47_adj_4723)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5158_8 (.CI(n53970), .I0(n20292[5]), .I1(n554_adj_4722), 
            .CO(n53971));
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_6_lut (.I0(GND_net), .I1(n16222[3]), .I2(n378_adj_4725), 
            .I3(n54725), .O(n15286[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[22]), 
            .I3(n53791), .O(n36[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n53631), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5158_7_lut (.I0(GND_net), .I1(n20292[4]), .I2(n481_adj_4727), 
            .I3(n53969), .O(n20115[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_7 (.CI(n53969), .I0(n20292[4]), .I1(n481_adj_4727), 
            .CO(n53970));
    SB_CARRY unary_minus_27_add_3_24 (.CI(n53791), .I0(GND_net), .I1(n1_adj_5002[22]), 
            .CO(n53792));
    SB_CARRY add_4867_6 (.CI(n54725), .I0(n16222[3]), .I1(n378_adj_4725), 
            .CO(n54726));
    SB_CARRY sub_15_add_2_5 (.CI(n53603), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n53604));
    SB_LUT4 add_5158_6_lut (.I0(GND_net), .I1(n20292[3]), .I2(n408_adj_4728), 
            .I3(n53968), .O(n20115[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_19_lut (.I0(GND_net), .I1(n16743[16]), .I2(GND_net), 
            .I3(n54278), .O(n15902[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_4 (.CI(n53602), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n53603));
    SB_CARRY sub_15_add_2_3 (.CI(n53601), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n53602));
    SB_CARRY add_5158_6 (.CI(n53968), .I0(n20292[3]), .I1(n408_adj_4728), 
            .CO(n53969));
    SB_LUT4 add_5158_5_lut (.I0(GND_net), .I1(n20292[2]), .I2(n335_adj_4729), 
            .I3(n53967), .O(n20115[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[21]), 
            .I3(n53790), .O(n36[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_5_lut (.I0(GND_net), .I1(n16222[2]), .I2(n305_adj_4732), 
            .I3(n54724), .O(n15286[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_18_lut (.I0(GND_net), .I1(n16743[15]), .I2(GND_net), 
            .I3(n54277), .O(n15902[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_18 (.CI(n54277), .I0(n16743[15]), .I1(GND_net), 
            .CO(n54278));
    SB_CARRY add_5158_5 (.CI(n53967), .I0(n20292[2]), .I1(n335_adj_4729), 
            .CO(n53968));
    SB_LUT4 add_5158_4_lut (.I0(GND_net), .I1(n20292[1]), .I2(n262_adj_4733), 
            .I3(n53966), .O(n20115[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n53790), .I0(GND_net), .I1(n1_adj_5002[21]), 
            .CO(n53791));
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5158_4 (.CI(n53966), .I0(n20292[1]), .I1(n262_adj_4733), 
            .CO(n53967));
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[20]), 
            .I3(n53789), .O(n36[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_22 (.CI(n53789), .I0(GND_net), .I1(n1_adj_5002[20]), 
            .CO(n53790));
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_10 (.CI(n53631), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n53632));
    SB_CARRY add_4867_5 (.CI(n54724), .I0(n16222[2]), .I1(n305_adj_4732), 
            .CO(n54725));
    SB_LUT4 add_4867_4_lut (.I0(GND_net), .I1(n16222[1]), .I2(n232_adj_4735), 
            .I3(n54723), .O(n15286[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_17_lut (.I0(GND_net), .I1(n16743[14]), .I2(GND_net), 
            .I3(n54276), .O(n15902[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_17 (.CI(n54276), .I0(n16743[14]), .I1(GND_net), 
            .CO(n54277));
    SB_LUT4 add_5158_3_lut (.I0(GND_net), .I1(n20292[0]), .I2(n189_adj_4736), 
            .I3(n53965), .O(n20115[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[19]), 
            .I3(n53788), .O(n36[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n53630), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_4 (.CI(n54723), .I0(n16222[1]), .I1(n232_adj_4735), 
            .CO(n54724));
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4867_3_lut (.I0(GND_net), .I1(n16222[0]), .I2(n159_adj_4739), 
            .I3(n54722), .O(n15286[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_16_lut (.I0(GND_net), .I1(n16743[13]), .I2(n1111), 
            .I3(n54275), .O(n15902[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_16 (.CI(n54275), .I0(n16743[13]), .I1(n1111), .CO(n54276));
    SB_CARRY add_5158_3 (.CI(n53965), .I0(n20292[0]), .I1(n189_adj_4736), 
            .CO(n53966));
    SB_LUT4 add_5158_2_lut (.I0(GND_net), .I1(n47_adj_4740), .I2(n116_adj_4741), 
            .I3(GND_net), .O(n20115[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_15_lut (.I0(GND_net), .I1(n16743[12]), .I2(n1038), 
            .I3(n54274), .O(n15902[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_15 (.CI(n54274), .I0(n16743[12]), .I1(n1038), .CO(n54275));
    SB_CARRY add_5158_2 (.CI(GND_net), .I0(n47_adj_4740), .I1(n116_adj_4741), 
            .CO(n53965));
    SB_CARRY unary_minus_27_add_3_21 (.CI(n53788), .I0(GND_net), .I1(n1_adj_5002[19]), 
            .CO(n53789));
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4867_3 (.CI(n54722), .I0(n16222[0]), .I1(n159_adj_4739), 
            .CO(n54723));
    SB_LUT4 add_4897_14_lut (.I0(GND_net), .I1(n16743[11]), .I2(n965), 
            .I3(n54273), .O(n15902[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[18]), 
            .I3(n53787), .O(n36[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_2_lut (.I0(GND_net), .I1(n17_adj_4744), .I2(n86_adj_4745), 
            .I3(GND_net), .O(n15286[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_14 (.CI(n54273), .I0(n16743[11]), .I1(n965), .CO(n54274));
    SB_CARRY unary_minus_27_add_3_20 (.CI(n53787), .I0(GND_net), .I1(n1_adj_5002[18]), 
            .CO(n53788));
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4897_13_lut (.I0(GND_net), .I1(n16743[10]), .I2(n892), 
            .I3(n54272), .O(n15902[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_13 (.CI(n54272), .I0(n16743[10]), .I1(n892), .CO(n54273));
    SB_CARRY add_4867_2 (.CI(GND_net), .I0(n17_adj_4744), .I1(n86_adj_4745), 
            .CO(n54722));
    SB_LUT4 add_4897_12_lut (.I0(GND_net), .I1(n16743[9]), .I2(n819), 
            .I3(n54271), .O(n15902[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_12 (.CI(n54271), .I0(n16743[9]), .I1(n819), .CO(n54272));
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[17]), 
            .I3(n53786), .O(n36[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_19_lut (.I0(GND_net), .I1(n17028[16]), .I2(GND_net), 
            .I3(n54721), .O(n16222[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_11_lut (.I0(GND_net), .I1(n16743[8]), .I2(n746), 
            .I3(n54270), .O(n15902[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n53786), .I0(GND_net), .I1(n1_adj_5002[17]), 
            .CO(n53787));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[16]), 
            .I3(n53785), .O(n36[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_18_lut (.I0(GND_net), .I1(n17028[15]), .I2(GND_net), 
            .I3(n54720), .O(n16222[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_11 (.CI(n54270), .I0(n16743[8]), .I1(n746), .CO(n54271));
    SB_LUT4 add_4897_10_lut (.I0(GND_net), .I1(n16743[7]), .I2(n673), 
            .I3(n54269), .O(n15902[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_18 (.CI(n53785), .I0(GND_net), .I1(n1_adj_5002[16]), 
            .CO(n53786));
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n352), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4748));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4750));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4751));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_18 (.CI(n54720), .I0(n17028[15]), .I1(GND_net), 
            .CO(n54721));
    SB_CARRY add_4897_10 (.CI(n54269), .I0(n16743[7]), .I1(n673), .CO(n54270));
    SB_LUT4 add_4897_9_lut (.I0(GND_net), .I1(n16743[6]), .I2(n600), .I3(n54268), 
            .O(n15902[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[15]), 
            .I3(n53784), .O(n36[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_17_lut (.I0(GND_net), .I1(n17028[14]), .I2(GND_net), 
            .I3(n54719), .O(n16222[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_9 (.CI(n54268), .I0(n16743[6]), .I1(n600), .CO(n54269));
    SB_LUT4 add_4897_8_lut (.I0(GND_net), .I1(n16743[5]), .I2(n527), .I3(n54267), 
            .O(n15902[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_9 (.CI(n53630), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n53631));
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_17 (.CI(n54719), .I0(n17028[14]), .I1(GND_net), 
            .CO(n54720));
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4897_8 (.CI(n54267), .I0(n16743[5]), .I1(n527), .CO(n54268));
    SB_LUT4 add_4913_16_lut (.I0(GND_net), .I1(n17028[13]), .I2(n1111_adj_4754), 
            .I3(n54718), .O(n16222[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_7_lut (.I0(GND_net), .I1(n16743[4]), .I2(n454), .I3(n54266), 
            .O(n15902[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_7 (.CI(n54266), .I0(n16743[4]), .I1(n454), .CO(n54267));
    SB_CARRY unary_minus_27_add_3_17 (.CI(n53784), .I0(GND_net), .I1(n1_adj_5002[15]), 
            .CO(n53785));
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_16 (.CI(n54718), .I0(n17028[13]), .I1(n1111_adj_4754), 
            .CO(n54719));
    SB_LUT4 add_4897_6_lut (.I0(GND_net), .I1(n16743[3]), .I2(n381), .I3(n54265), 
            .O(n15902[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_15_lut (.I0(GND_net), .I1(n17028[12]), .I2(n1038_adj_4755), 
            .I3(n54717), .O(n16222[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_6 (.CI(n54265), .I0(n16743[3]), .I1(n381), .CO(n54266));
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[14]), 
            .I3(n53783), .O(n36[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n53783), .I0(GND_net), .I1(n1_adj_5002[14]), 
            .CO(n53784));
    SB_CARRY add_4913_15 (.CI(n54717), .I0(n17028[12]), .I1(n1038_adj_4755), 
            .CO(n54718));
    SB_LUT4 add_4897_5_lut (.I0(GND_net), .I1(n16743[2]), .I2(n308_adj_4757), 
            .I3(n54264), .O(n15902[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_5 (.CI(n54264), .I0(n16743[2]), .I1(n308_adj_4757), 
            .CO(n54265));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[13]), 
            .I3(n53782), .O(n36[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4913_14_lut (.I0(GND_net), .I1(n17028[11]), .I2(n965_adj_4759), 
            .I3(n54716), .O(n16222[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_4_lut (.I0(GND_net), .I1(n16743[1]), .I2(n235_adj_4760), 
            .I3(n54263), .O(n15902[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_4 (.CI(n54263), .I0(n16743[1]), .I1(n235_adj_4760), 
            .CO(n54264));
    SB_CARRY unary_minus_27_add_3_15 (.CI(n53782), .I0(GND_net), .I1(n1_adj_5002[13]), 
            .CO(n53783));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n53629), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_8 (.CI(n53629), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n53630));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[12]), 
            .I3(n53781), .O(n36[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_14 (.CI(n54716), .I0(n17028[11]), .I1(n965_adj_4759), 
            .CO(n54717));
    SB_LUT4 add_4897_3_lut (.I0(GND_net), .I1(n16743[0]), .I2(n162), .I3(n54262), 
            .O(n15902[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_3 (.CI(n54262), .I0(n16743[0]), .I1(n162), .CO(n54263));
    SB_LUT4 add_4913_13_lut (.I0(GND_net), .I1(n17028[10]), .I2(n892_adj_4762), 
            .I3(n54715), .O(n16222[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4897_2_lut (.I0(GND_net), .I1(n20_adj_4763), .I2(n89), 
            .I3(GND_net), .O(n15902[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4897_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n53781), .I0(GND_net), .I1(n1_adj_5002[12]), 
            .CO(n53782));
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[11]), 
            .I3(n53780), .O(n36[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4765));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4766));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_13 (.CI(n54715), .I0(n17028[10]), .I1(n892_adj_4762), 
            .CO(n54716));
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4767));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4768));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4769));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4770));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4771));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4772));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4773));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4913_12_lut (.I0(GND_net), .I1(n17028[9]), .I2(n819_adj_4774), 
            .I3(n54714), .O(n16222[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4775));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4776));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4777));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4778));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4779));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4780));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4781));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4913_12 (.CI(n54714), .I0(n17028[9]), .I1(n819_adj_4774), 
            .CO(n54715));
    SB_LUT4 add_4913_11_lut (.I0(GND_net), .I1(n17028[8]), .I2(n746_adj_4782), 
            .I3(n54713), .O(n16222[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_13 (.CI(n53780), .I0(GND_net), .I1(n1_adj_5002[11]), 
            .CO(n53781));
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[10]), 
            .I3(n53779), .O(n36[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n53779), .I0(GND_net), .I1(n1_adj_5002[10]), 
            .CO(n53780));
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[9]), 
            .I3(n53778), .O(n36[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4913_11 (.CI(n54713), .I0(n17028[8]), .I1(n746_adj_4782), 
            .CO(n54714));
    SB_CARRY unary_minus_27_add_3_11 (.CI(n53778), .I0(GND_net), .I1(n1_adj_5002[9]), 
            .CO(n53779));
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n53628), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n71969_bdd_4_lut (.I0(n71969), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4743), .O(n71972));
    defparam n71969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_16_7 (.CI(n53628), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n53629));
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[8]), 
            .I3(n53777), .O(n36[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4897_2 (.CI(GND_net), .I0(n20_adj_4763), .I1(n89), .CO(n54262));
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4786));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4787));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4788));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4789));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4790));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4791));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4792));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4793));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4794));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4795));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4796));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4797));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4798));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n53627), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_10 (.CI(n53777), .I0(GND_net), .I1(n1_adj_5002[8]), 
            .CO(n53778));
    SB_LUT4 add_4913_10_lut (.I0(GND_net), .I1(n17028[7]), .I2(n673_adj_4799), 
            .I3(n54712), .O(n16222[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4800));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n53601));
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[7]), 
            .I3(n53776), .O(n36[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n53776), .I0(GND_net), .I1(n1_adj_5002[7]), 
            .CO(n53777));
    SB_CARRY add_4913_10 (.CI(n54712), .I0(n17028[7]), .I1(n673_adj_4799), 
            .CO(n54713));
    SB_LUT4 add_4913_9_lut (.I0(GND_net), .I1(n17028[6]), .I2(n600_adj_4802), 
            .I3(n54711), .O(n16222[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4913_9 (.CI(n54711), .I0(n17028[6]), .I1(n600_adj_4802), 
            .CO(n54712));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[6]), 
            .I3(n53775), .O(n36[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_6 (.CI(n53627), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n53628));
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n53626), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_8 (.CI(n53775), .I0(GND_net), .I1(n1_adj_5002[6]), 
            .CO(n53776));
    SB_LUT4 add_4913_8_lut (.I0(GND_net), .I1(n17028[5]), .I2(n527_adj_4804), 
            .I3(n54710), .O(n16222[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[5]), 
            .I3(n53774), .O(n36[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_5 (.CI(n53626), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n53627));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n53625), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n53774), .I0(GND_net), .I1(n1_adj_5002[5]), 
            .CO(n53775));
    SB_CARRY add_4913_8 (.CI(n54710), .I0(n17028[5]), .I1(n527_adj_4804), 
            .CO(n54711));
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[4]), 
            .I3(n53773), .O(n36[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_6 (.CI(n53773), .I0(GND_net), .I1(n1_adj_5002[4]), 
            .CO(n53774));
    SB_LUT4 add_4913_7_lut (.I0(GND_net), .I1(n17028[4]), .I2(n454_adj_4807), 
            .I3(n54709), .O(n16222[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[3]), 
            .I3(n53772), .O(n36[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n53772), .I0(GND_net), .I1(n1_adj_5002[3]), 
            .CO(n53773));
    SB_CARRY add_4913_7 (.CI(n54709), .I0(n17028[4]), .I1(n454_adj_4807), 
            .CO(n54710));
    SB_LUT4 add_4913_6_lut (.I0(GND_net), .I1(n17028[3]), .I2(n381_adj_4809), 
            .I3(n54708), .O(n16222[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4913_6 (.CI(n54708), .I0(n17028[3]), .I1(n381_adj_4809), 
            .CO(n54709));
    SB_LUT4 add_4913_5_lut (.I0(GND_net), .I1(n17028[2]), .I2(n308_adj_4810), 
            .I3(n54707), .O(n16222[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4913_5 (.CI(n54707), .I0(n17028[2]), .I1(n308_adj_4810), 
            .CO(n54708));
    SB_CARRY add_16_4 (.CI(n53625), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n53626));
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[2]), 
            .I3(n53771), .O(n36[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_4_lut (.I0(GND_net), .I1(n17028[1]), .I2(n235_adj_4812), 
            .I3(n54706), .O(n16222[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n53624), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_4 (.CI(n53771), .I0(GND_net), .I1(n1_adj_5002[2]), 
            .CO(n53772));
    SB_CARRY add_4913_4 (.CI(n54706), .I0(n17028[1]), .I1(n235_adj_4812), 
            .CO(n54707));
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4813));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5002[1]), 
            .I3(n53770), .O(n36[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4913_3_lut (.I0(GND_net), .I1(n17028[0]), .I2(n162_adj_4815), 
            .I3(n54705), .O(n16222[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n53770), .I0(GND_net), .I1(n1_adj_5002[1]), 
            .CO(n53771));
    SB_CARRY add_4913_3 (.CI(n54705), .I0(n17028[0]), .I1(n162_adj_4815), 
            .CO(n54706));
    SB_LUT4 add_4913_2_lut (.I0(GND_net), .I1(n20_adj_4816), .I2(n89_adj_4817), 
            .I3(GND_net), .O(n16222[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4913_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4913_2 (.CI(GND_net), .I0(n20_adj_4816), .I1(n89_adj_4817), 
            .CO(n54705));
    SB_LUT4 add_4954_18_lut (.I0(GND_net), .I1(n17714[15]), .I2(GND_net), 
            .I3(n54704), .O(n17028[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_17_lut (.I0(GND_net), .I1(n17714[14]), .I2(GND_net), 
            .I3(n54703), .O(n17028[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_3 (.CI(n53624), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n53625));
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n39485), .I1(GND_net), .I2(n1_adj_5002[0]), 
            .I3(VCC_net), .O(n68301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5002[0]), 
            .CO(n53770));
    SB_CARRY add_4954_17 (.CI(n54703), .I0(n17714[14]), .I1(GND_net), 
            .CO(n54704));
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n53624));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[23]), 
            .I3(n53769), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[22]), 
            .I3(n53768), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n53768), .I0(GND_net), .I1(n1_adj_5003[22]), 
            .CO(n53769));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[21]), 
            .I3(n53767), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_16_lut (.I0(GND_net), .I1(n17714[13]), .I2(n1114_adj_4823), 
            .I3(n54702), .O(n17028[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n53767), .I0(GND_net), .I1(n1_adj_5003[21]), 
            .CO(n53768));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[20]), 
            .I3(n53766), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n53766), .I0(GND_net), .I1(n1_adj_5003[20]), 
            .CO(n53767));
    SB_CARRY add_4954_16 (.CI(n54702), .I0(n17714[13]), .I1(n1114_adj_4823), 
            .CO(n54703));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[19]), 
            .I3(n53765), .O(n290)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n53765), .I0(GND_net), .I1(n1_adj_5003[19]), 
            .CO(n53766));
    SB_LUT4 add_4954_15_lut (.I0(GND_net), .I1(n17714[12]), .I2(n1041_adj_4826), 
            .I3(n54701), .O(n17028[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(n17_adj_1), 
            .I3(n53623), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n53622), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[18]), 
            .I3(n53764), .O(n285[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n53764), .I0(GND_net), .I1(n1_adj_5003[18]), 
            .CO(n53765));
    SB_CARRY add_4954_15 (.CI(n54701), .I0(n17714[12]), .I1(n1041_adj_4826), 
            .CO(n54702));
    SB_CARRY sub_15_add_2_24 (.CI(n53622), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n53623));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[17]), 
            .I3(n53763), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n53763), .I0(GND_net), .I1(n1_adj_5003[17]), 
            .CO(n53764));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[16]), 
            .I3(n53762), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n53762), .I0(GND_net), .I1(n1_adj_5003[16]), 
            .CO(n53763));
    SB_LUT4 add_4954_14_lut (.I0(GND_net), .I1(n17714[11]), .I2(n968_adj_4831), 
            .I3(n54700), .O(n17028[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[15]), 
            .I3(n53761), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_14 (.CI(n54700), .I0(n17714[11]), .I1(n968_adj_4831), 
            .CO(n54701));
    SB_LUT4 add_4954_13_lut (.I0(GND_net), .I1(n17714[10]), .I2(n895_adj_4833), 
            .I3(n54699), .O(n17028[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n53621), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_23 (.CI(n53621), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n53622));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n53761), .I0(GND_net), .I1(n1_adj_5003[15]), 
            .CO(n53762));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[14]), 
            .I3(n53760), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_13 (.CI(n54699), .I0(n17714[10]), .I1(n895_adj_4833), 
            .CO(n54700));
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n53620), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_22 (.CI(n53620), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n53621));
    SB_CARRY unary_minus_20_add_3_16 (.CI(n53760), .I0(GND_net), .I1(n1_adj_5003[14]), 
            .CO(n53761));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[13]), 
            .I3(n53759), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_12_lut (.I0(GND_net), .I1(n17714[9]), .I2(n822_adj_4836), 
            .I3(n54698), .O(n17028[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n53759), .I0(GND_net), .I1(n1_adj_5003[13]), 
            .CO(n53760));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[12]), 
            .I3(n53758), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_12 (.CI(n54698), .I0(n17714[9]), .I1(n822_adj_4836), 
            .CO(n54699));
    SB_CARRY unary_minus_20_add_3_14 (.CI(n53758), .I0(GND_net), .I1(n1_adj_5003[12]), 
            .CO(n53759));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[11]), 
            .I3(n53757), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_11_lut (.I0(GND_net), .I1(n17714[8]), .I2(n749_adj_4839), 
            .I3(n54697), .O(n17028[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n53757), .I0(GND_net), .I1(n1_adj_5003[11]), 
            .CO(n53758));
    SB_CARRY add_4954_11 (.CI(n54697), .I0(n17714[8]), .I1(n749_adj_4839), 
            .CO(n54698));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[10]), 
            .I3(n53756), .O(n285[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_10_lut (.I0(GND_net), .I1(n17714[7]), .I2(n676_adj_4841), 
            .I3(n54696), .O(n17028[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4842));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n53756), .I0(GND_net), .I1(n1_adj_5003[10]), 
            .CO(n53757));
    SB_CARRY add_4954_10 (.CI(n54696), .I0(n17714[7]), .I1(n676_adj_4841), 
            .CO(n54697));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[9]), 
            .I3(n53755), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_9_lut (.I0(GND_net), .I1(n17714[6]), .I2(n603_adj_4844), 
            .I3(n54695), .O(n17028[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4845));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4846));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n53619), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_21 (.CI(n53619), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n53620));
    SB_CARRY unary_minus_20_add_3_11 (.CI(n53755), .I0(GND_net), .I1(n1_adj_5003[9]), 
            .CO(n53756));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[8]), 
            .I3(n53754), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_9 (.CI(n54695), .I0(n17714[6]), .I1(n603_adj_4844), 
            .CO(n54696));
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n53618), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n53618), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n53619));
    SB_CARRY unary_minus_20_add_3_10 (.CI(n53754), .I0(GND_net), .I1(n1_adj_5003[8]), 
            .CO(n53755));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[7]), 
            .I3(n53753), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_8_lut (.I0(GND_net), .I1(n17714[5]), .I2(n530_adj_4849), 
            .I3(n54694), .O(n17028[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n53753), .I0(GND_net), .I1(n1_adj_5003[7]), 
            .CO(n53754));
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[6]), 
            .I3(n53752), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_8 (.CI(n54694), .I0(n17714[5]), .I1(n530_adj_4849), 
            .CO(n54695));
    SB_CARRY unary_minus_20_add_3_8 (.CI(n53752), .I0(GND_net), .I1(n1_adj_5003[6]), 
            .CO(n53753));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[5]), 
            .I3(n53751), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_7_lut (.I0(GND_net), .I1(n17714[4]), .I2(n457_adj_4852), 
            .I3(n54693), .O(n17028[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_7 (.CI(n54693), .I0(n17714[4]), .I1(n457_adj_4852), 
            .CO(n54694));
    SB_LUT4 add_4954_6_lut (.I0(GND_net), .I1(n17714[3]), .I2(n384_adj_4853), 
            .I3(n54692), .O(n17028[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_6 (.CI(n54692), .I0(n17714[3]), .I1(n384_adj_4853), 
            .CO(n54693));
    SB_LUT4 add_4954_5_lut (.I0(GND_net), .I1(n17714[2]), .I2(n311_adj_4854), 
            .I3(n54691), .O(n17028[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4855));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n53751), .I0(GND_net), .I1(n1_adj_5003[5]), 
            .CO(n53752));
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[4]), 
            .I3(n53750), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n53750), .I0(GND_net), .I1(n1_adj_5003[4]), 
            .CO(n53751));
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n53617), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_19 (.CI(n53617), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n53618));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[3]), 
            .I3(n53749), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_5 (.CI(n54691), .I0(n17714[2]), .I1(n311_adj_4854), 
            .CO(n54692));
    SB_CARRY unary_minus_20_add_3_5 (.CI(n53749), .I0(GND_net), .I1(n1_adj_5003[3]), 
            .CO(n53750));
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n53616), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[2]), 
            .I3(n53748), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n53748), .I0(GND_net), .I1(n1_adj_5003[2]), 
            .CO(n53749));
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[1]), 
            .I3(n53747), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4954_4_lut (.I0(GND_net), .I1(n17714[1]), .I2(n238_adj_4860), 
            .I3(n54690), .O(n17028[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4861));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_20_add_3_3 (.CI(n53747), .I0(GND_net), .I1(n1_adj_5003[1]), 
            .CO(n53748));
    SB_CARRY add_4954_4 (.CI(n54690), .I0(n17714[1]), .I1(n238_adj_4860), 
            .CO(n54691));
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4862));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4954_3_lut (.I0(GND_net), .I1(n17714[0]), .I2(n165_adj_4863), 
            .I3(n54689), .O(n17028[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5003[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n53616), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n53617));
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n53615), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5003[0]), 
            .CO(n53747));
    SB_CARRY add_4954_3 (.CI(n54689), .I0(n17714[0]), .I1(n165_adj_4863), 
            .CO(n54690));
    SB_CARRY sub_15_add_2_17 (.CI(n53615), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n53616));
    SB_LUT4 add_4954_2_lut (.I0(GND_net), .I1(n23_adj_4865), .I2(n92_adj_4866), 
            .I3(GND_net), .O(n17028[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4954_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4954_2 (.CI(GND_net), .I0(n23_adj_4865), .I1(n92_adj_4866), 
            .CO(n54689));
    SB_LUT4 add_4991_17_lut (.I0(GND_net), .I1(n18276[14]), .I2(GND_net), 
            .I3(n54688), .O(n17714[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4867));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4868));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n53614), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_16 (.CI(n53614), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n53615));
    SB_LUT4 add_4991_16_lut (.I0(GND_net), .I1(n18276[13]), .I2(n1117_adj_4869), 
            .I3(n54687), .O(n17714[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n53613), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n53613), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n53614));
    SB_LUT4 add_5175_9_lut (.I0(GND_net), .I1(n20433[6]), .I2(n630_adj_4870), 
            .I3(n53915), .O(n20292[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_16 (.CI(n54687), .I0(n18276[13]), .I1(n1117_adj_4869), 
            .CO(n54688));
    SB_LUT4 add_5175_8_lut (.I0(GND_net), .I1(n20433[5]), .I2(n557_adj_4871), 
            .I3(n53914), .O(n20292[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_15_lut (.I0(GND_net), .I1(n18276[12]), .I2(n1044_adj_4872), 
            .I3(n54686), .O(n17714[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_8 (.CI(n53914), .I0(n20433[5]), .I1(n557_adj_4871), 
            .CO(n53915));
    SB_CARRY add_4991_15 (.CI(n54686), .I0(n18276[12]), .I1(n1044_adj_4872), 
            .CO(n54687));
    SB_LUT4 add_5175_7_lut (.I0(GND_net), .I1(n20433[4]), .I2(n484_adj_4873), 
            .I3(n53913), .O(n20292[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_14_lut (.I0(GND_net), .I1(n18276[11]), .I2(n971_adj_4874), 
            .I3(n54685), .O(n17714[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_7 (.CI(n53913), .I0(n20433[4]), .I1(n484_adj_4873), 
            .CO(n53914));
    SB_CARRY add_4991_14 (.CI(n54685), .I0(n18276[11]), .I1(n971_adj_4874), 
            .CO(n54686));
    SB_LUT4 add_5175_6_lut (.I0(GND_net), .I1(n20433[3]), .I2(n411_adj_4875), 
            .I3(n53912), .O(n20292[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_13_lut (.I0(GND_net), .I1(n18276[10]), .I2(n898_adj_4876), 
            .I3(n54684), .O(n17714[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_6 (.CI(n53912), .I0(n20433[3]), .I1(n411_adj_4875), 
            .CO(n53913));
    SB_CARRY add_4991_13 (.CI(n54684), .I0(n18276[10]), .I1(n898_adj_4876), 
            .CO(n54685));
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4877));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n53612), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n53612), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n53613));
    SB_LUT4 add_5175_5_lut (.I0(GND_net), .I1(n20433[2]), .I2(n338_adj_4878), 
            .I3(n53911), .O(n20292[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_12_lut (.I0(GND_net), .I1(n18276[9]), .I2(n825_adj_4879), 
            .I3(n54683), .O(n17714[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(n3), 
            .I3(n53611), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n53611), .I0(setpoint[11]), .I1(n3), 
            .CO(n53612));
    SB_CARRY add_5175_5 (.CI(n53911), .I0(n20433[2]), .I1(n338_adj_4878), 
            .CO(n53912));
    SB_CARRY add_4991_12 (.CI(n54683), .I0(n18276[9]), .I1(n825_adj_4879), 
            .CO(n54684));
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4881));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5175_4_lut (.I0(GND_net), .I1(n20433[1]), .I2(n265_adj_4882), 
            .I3(n53910), .O(n20292[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_11_lut (.I0(GND_net), .I1(n18276[8]), .I2(n752_adj_4883), 
            .I3(n54682), .O(n17714[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_4 (.CI(n53910), .I0(n20433[1]), .I1(n265_adj_4882), 
            .CO(n53911));
    SB_CARRY add_4991_11 (.CI(n54682), .I0(n18276[8]), .I1(n752_adj_4883), 
            .CO(n54683));
    SB_LUT4 add_5175_3_lut (.I0(GND_net), .I1(n20433[0]), .I2(n192_adj_4884), 
            .I3(n53909), .O(n20292[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_10_lut (.I0(GND_net), .I1(n18276[7]), .I2(n679_adj_4885), 
            .I3(n54681), .O(n17714[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_3 (.CI(n53909), .I0(n20433[0]), .I1(n192_adj_4884), 
            .CO(n53910));
    SB_CARRY add_4991_10 (.CI(n54681), .I0(n18276[7]), .I1(n679_adj_4885), 
            .CO(n54682));
    SB_LUT4 add_5175_2_lut (.I0(GND_net), .I1(n50_adj_4886), .I2(n119_adj_4887), 
            .I3(GND_net), .O(n20292[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5175_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_9_lut (.I0(GND_net), .I1(n18276[6]), .I2(n606_adj_4888), 
            .I3(n54680), .O(n17714[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5175_2 (.CI(GND_net), .I0(n50_adj_4886), .I1(n119_adj_4887), 
            .CO(n53909));
    SB_CARRY add_4991_9 (.CI(n54680), .I0(n18276[6]), .I1(n606_adj_4888), 
            .CO(n54681));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n53610), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4991_8_lut (.I0(GND_net), .I1(n18276[5]), .I2(n533_adj_4889), 
            .I3(n54679), .O(n17714[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4890));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4891));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4991_8 (.CI(n54679), .I0(n18276[5]), .I1(n533_adj_4889), 
            .CO(n54680));
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4892));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4991_7_lut (.I0(GND_net), .I1(n18276[4]), .I2(n460_adj_4893), 
            .I3(n54678), .O(n17714[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_7 (.CI(n54678), .I0(n18276[4]), .I1(n460_adj_4893), 
            .CO(n54679));
    SB_LUT4 mult_24_i38_2_lut (.I0(\Ki[0] ), .I1(n341), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4894));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4991_6_lut (.I0(GND_net), .I1(n18276[3]), .I2(n387_adj_4895), 
            .I3(n54677), .O(n17714[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_6 (.CI(n54677), .I0(n18276[3]), .I1(n387_adj_4895), 
            .CO(n54678));
    SB_LUT4 add_4991_5_lut (.I0(GND_net), .I1(n18276[2]), .I2(n314_adj_4896), 
            .I3(n54676), .O(n17714[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_5 (.CI(n54676), .I0(n18276[2]), .I1(n314_adj_4896), 
            .CO(n54677));
    SB_LUT4 add_4991_4_lut (.I0(GND_net), .I1(n18276[1]), .I2(n241_adj_4897), 
            .I3(n54675), .O(n17714[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_4 (.CI(n54675), .I0(n18276[1]), .I1(n241_adj_4897), 
            .CO(n54676));
    SB_LUT4 add_4991_3_lut (.I0(GND_net), .I1(n18276[0]), .I2(n168_adj_4898), 
            .I3(n54674), .O(n17714[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_3 (.CI(n54674), .I0(n18276[0]), .I1(n168_adj_4898), 
            .CO(n54675));
    SB_LUT4 add_4991_2_lut (.I0(GND_net), .I1(n26_adj_4899), .I2(n95_adj_4900), 
            .I3(GND_net), .O(n17714[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4991_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4991_2 (.CI(GND_net), .I0(n26_adj_4899), .I1(n95_adj_4900), 
            .CO(n54674));
    SB_LUT4 add_5025_16_lut (.I0(GND_net), .I1(n18728[13]), .I2(n1120_adj_4901), 
            .I3(n54673), .O(n18276[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5025_15_lut (.I0(GND_net), .I1(n18728[12]), .I2(n1047_adj_4902), 
            .I3(n54672), .O(n18276[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_15 (.CI(n54672), .I0(n18728[12]), .I1(n1047_adj_4902), 
            .CO(n54673));
    SB_LUT4 add_5025_14_lut (.I0(GND_net), .I1(n18728[11]), .I2(n974_adj_4903), 
            .I3(n54671), .O(n18276[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_14 (.CI(n54671), .I0(n18728[11]), .I1(n974_adj_4903), 
            .CO(n54672));
    SB_LUT4 add_5025_13_lut (.I0(GND_net), .I1(n18728[10]), .I2(n901_adj_4904), 
            .I3(n54670), .O(n18276[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_13 (.CI(n54670), .I0(n18728[10]), .I1(n901_adj_4904), 
            .CO(n54671));
    SB_LUT4 add_5025_12_lut (.I0(GND_net), .I1(n18728[9]), .I2(n828_adj_4905), 
            .I3(n54669), .O(n18276[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_12 (.CI(n54669), .I0(n18728[9]), .I1(n828_adj_4905), 
            .CO(n54670));
    SB_LUT4 add_5025_11_lut (.I0(GND_net), .I1(n18728[8]), .I2(n755_adj_4906), 
            .I3(n54668), .O(n18276[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_11 (.CI(n54668), .I0(n18728[8]), .I1(n755_adj_4906), 
            .CO(n54669));
    SB_LUT4 add_5025_10_lut (.I0(GND_net), .I1(n18728[7]), .I2(n682_adj_4907), 
            .I3(n54667), .O(n18276[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_10 (.CI(n54667), .I0(n18728[7]), .I1(n682_adj_4907), 
            .CO(n54668));
    SB_LUT4 add_5025_9_lut (.I0(GND_net), .I1(n18728[6]), .I2(n609_adj_4908), 
            .I3(n54666), .O(n18276[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_9 (.CI(n54666), .I0(n18728[6]), .I1(n609_adj_4908), 
            .CO(n54667));
    SB_LUT4 add_5025_8_lut (.I0(GND_net), .I1(n18728[5]), .I2(n536_adj_4909), 
            .I3(n54665), .O(n18276[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_8 (.CI(n54665), .I0(n18728[5]), .I1(n536_adj_4909), 
            .CO(n54666));
    SB_LUT4 add_5025_7_lut (.I0(GND_net), .I1(n18728[4]), .I2(n463_adj_4910), 
            .I3(n54664), .O(n18276[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_7 (.CI(n54664), .I0(n18728[4]), .I1(n463_adj_4910), 
            .CO(n54665));
    SB_LUT4 add_5025_6_lut (.I0(GND_net), .I1(n18728[3]), .I2(n390_adj_4911), 
            .I3(n54663), .O(n18276[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_6 (.CI(n54663), .I0(n18728[3]), .I1(n390_adj_4911), 
            .CO(n54664));
    SB_LUT4 add_5025_5_lut (.I0(GND_net), .I1(n18728[2]), .I2(n317_adj_4912), 
            .I3(n54662), .O(n18276[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_5 (.CI(n54662), .I0(n18728[2]), .I1(n317_adj_4912), 
            .CO(n54663));
    SB_LUT4 add_5025_4_lut (.I0(GND_net), .I1(n18728[1]), .I2(n244_adj_4913), 
            .I3(n54661), .O(n18276[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_4 (.CI(n54661), .I0(n18728[1]), .I1(n244_adj_4913), 
            .CO(n54662));
    SB_LUT4 add_5025_3_lut (.I0(GND_net), .I1(n18728[0]), .I2(n171_adj_4914), 
            .I3(n54660), .O(n18276[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_3 (.CI(n54660), .I0(n18728[0]), .I1(n171_adj_4914), 
            .CO(n54661));
    SB_LUT4 add_5025_2_lut (.I0(GND_net), .I1(n29_adj_4915), .I2(n98_adj_4916), 
            .I3(GND_net), .O(n18276[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5025_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5025_2 (.CI(GND_net), .I0(n29_adj_4915), .I1(n98_adj_4916), 
            .CO(n54660));
    SB_LUT4 add_5203_7_lut (.I0(GND_net), .I1(n62699), .I2(n490_adj_4917), 
            .I3(n54659), .O(n20542[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5203_6_lut (.I0(GND_net), .I1(n20623[3]), .I2(n417_adj_4918), 
            .I3(n54658), .O(n20542[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_6 (.CI(n54658), .I0(n20623[3]), .I1(n417_adj_4918), 
            .CO(n54659));
    SB_LUT4 add_5203_5_lut (.I0(GND_net), .I1(n20623[2]), .I2(n344_adj_4919), 
            .I3(n54657), .O(n20542[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_5 (.CI(n54657), .I0(n20623[2]), .I1(n344_adj_4919), 
            .CO(n54658));
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4920));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_15_add_2_12 (.CI(n53610), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n53611));
    SB_LUT4 add_5203_4_lut (.I0(GND_net), .I1(n20623[1]), .I2(n271_adj_4921), 
            .I3(n54656), .O(n20542[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_4 (.CI(n54656), .I0(n20623[1]), .I1(n271_adj_4921), 
            .CO(n54657));
    SB_LUT4 add_5203_3_lut (.I0(GND_net), .I1(n20628), .I2(n198_adj_4922), 
            .I3(n54655), .O(n20542[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_3 (.CI(n54655), .I0(n20628), .I1(n198_adj_4922), 
            .CO(n54656));
    SB_LUT4 add_5203_2_lut (.I0(GND_net), .I1(n56_adj_4894), .I2(n125_adj_4892), 
            .I3(GND_net), .O(n20542[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_2 (.CI(GND_net), .I0(n56_adj_4894), .I1(n125_adj_4892), 
            .CO(n54655));
    SB_LUT4 add_5055_15_lut (.I0(GND_net), .I1(n19132[12]), .I2(n1050_adj_4891), 
            .I3(n54654), .O(n18728[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5055_14_lut (.I0(GND_net), .I1(n19132[11]), .I2(n977_adj_4890), 
            .I3(n54653), .O(n18728[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_14 (.CI(n54653), .I0(n19132[11]), .I1(n977_adj_4890), 
            .CO(n54654));
    SB_LUT4 add_5055_13_lut (.I0(GND_net), .I1(n19132[10]), .I2(n904_adj_4881), 
            .I3(n54652), .O(n18728[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_13 (.CI(n54652), .I0(n19132[10]), .I1(n904_adj_4881), 
            .CO(n54653));
    SB_LUT4 add_5055_12_lut (.I0(GND_net), .I1(n19132[9]), .I2(n831_adj_4877), 
            .I3(n54651), .O(n18728[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_12 (.CI(n54651), .I0(n19132[9]), .I1(n831_adj_4877), 
            .CO(n54652));
    SB_LUT4 add_5055_11_lut (.I0(GND_net), .I1(n19132[8]), .I2(n758_adj_4868), 
            .I3(n54650), .O(n18728[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_11 (.CI(n54650), .I0(n19132[8]), .I1(n758_adj_4868), 
            .CO(n54651));
    SB_LUT4 add_5055_10_lut (.I0(GND_net), .I1(n19132[7]), .I2(n685_adj_4867), 
            .I3(n54649), .O(n18728[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_10 (.CI(n54649), .I0(n19132[7]), .I1(n685_adj_4867), 
            .CO(n54650));
    SB_LUT4 add_5055_9_lut (.I0(GND_net), .I1(n19132[6]), .I2(n612_adj_4862), 
            .I3(n54648), .O(n18728[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_9 (.CI(n54648), .I0(n19132[6]), .I1(n612_adj_4862), 
            .CO(n54649));
    SB_LUT4 add_5055_8_lut (.I0(GND_net), .I1(n19132[5]), .I2(n539_adj_4855), 
            .I3(n54647), .O(n18728[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_8 (.CI(n54647), .I0(n19132[5]), .I1(n539_adj_4855), 
            .CO(n54648));
    SB_LUT4 add_5055_7_lut (.I0(GND_net), .I1(n19132[4]), .I2(n466_adj_4845), 
            .I3(n54646), .O(n18728[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_7 (.CI(n54646), .I0(n19132[4]), .I1(n466_adj_4845), 
            .CO(n54647));
    SB_LUT4 add_5055_6_lut (.I0(GND_net), .I1(n19132[3]), .I2(n393_adj_4842), 
            .I3(n54645), .O(n18728[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4923));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5055_6 (.CI(n54645), .I0(n19132[3]), .I1(n393_adj_4842), 
            .CO(n54646));
    SB_LUT4 add_5055_5_lut (.I0(GND_net), .I1(n19132[2]), .I2(n320_adj_4819), 
            .I3(n54644), .O(n18728[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_5 (.CI(n54644), .I0(n19132[2]), .I1(n320_adj_4819), 
            .CO(n54645));
    SB_LUT4 add_5055_4_lut (.I0(GND_net), .I1(n19132[1]), .I2(n247_adj_4813), 
            .I3(n54643), .O(n18728[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_4 (.CI(n54643), .I0(n19132[1]), .I1(n247_adj_4813), 
            .CO(n54644));
    SB_LUT4 add_5055_3_lut (.I0(GND_net), .I1(n19132[0]), .I2(n174_adj_4800), 
            .I3(n54642), .O(n18728[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_3 (.CI(n54642), .I0(n19132[0]), .I1(n174_adj_4800), 
            .CO(n54643));
    SB_LUT4 add_5055_2_lut (.I0(GND_net), .I1(n32_adj_4797), .I2(n101_adj_4796), 
            .I3(GND_net), .O(n18728[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5055_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5055_2 (.CI(GND_net), .I0(n32_adj_4797), .I1(n101_adj_4796), 
            .CO(n54642));
    SB_LUT4 add_5081_14_lut (.I0(GND_net), .I1(n19468[11]), .I2(n980_adj_4795), 
            .I3(n54641), .O(n19132[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5081_13_lut (.I0(GND_net), .I1(n19468[10]), .I2(n907_adj_4794), 
            .I3(n54640), .O(n19132[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_13 (.CI(n54640), .I0(n19468[10]), .I1(n907_adj_4794), 
            .CO(n54641));
    SB_LUT4 add_5081_12_lut (.I0(GND_net), .I1(n19468[9]), .I2(n834_adj_4792), 
            .I3(n54639), .O(n19132[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_12 (.CI(n54639), .I0(n19468[9]), .I1(n834_adj_4792), 
            .CO(n54640));
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4924));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5081_11_lut (.I0(GND_net), .I1(n19468[8]), .I2(n761_adj_4791), 
            .I3(n54638), .O(n19132[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_11 (.CI(n54638), .I0(n19468[8]), .I1(n761_adj_4791), 
            .CO(n54639));
    SB_LUT4 add_5081_10_lut (.I0(GND_net), .I1(n19468[7]), .I2(n688_adj_4790), 
            .I3(n54637), .O(n19132[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_10 (.CI(n54637), .I0(n19468[7]), .I1(n688_adj_4790), 
            .CO(n54638));
    SB_LUT4 add_5081_9_lut (.I0(GND_net), .I1(n19468[6]), .I2(n615_adj_4789), 
            .I3(n54636), .O(n19132[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_9 (.CI(n54636), .I0(n19468[6]), .I1(n615_adj_4789), 
            .CO(n54637));
    SB_LUT4 add_5081_8_lut (.I0(GND_net), .I1(n19468[5]), .I2(n542_adj_4788), 
            .I3(n54635), .O(n19132[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_8 (.CI(n54635), .I0(n19468[5]), .I1(n542_adj_4788), 
            .CO(n54636));
    SB_LUT4 add_5081_7_lut (.I0(GND_net), .I1(n19468[4]), .I2(n469_adj_4787), 
            .I3(n54634), .O(n19132[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_7 (.CI(n54634), .I0(n19468[4]), .I1(n469_adj_4787), 
            .CO(n54635));
    SB_LUT4 add_5081_6_lut (.I0(GND_net), .I1(n19468[3]), .I2(n396_adj_4786), 
            .I3(n54633), .O(n19132[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_6 (.CI(n54633), .I0(n19468[3]), .I1(n396_adj_4786), 
            .CO(n54634));
    SB_LUT4 add_5081_5_lut (.I0(GND_net), .I1(n19468[2]), .I2(n323_adj_4781), 
            .I3(n54632), .O(n19132[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_5 (.CI(n54632), .I0(n19468[2]), .I1(n323_adj_4781), 
            .CO(n54633));
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n10961[0]), .I2(n10332[0]), 
            .I3(n53669), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n1[22]), .I3(n53668), 
            .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_24 (.CI(n53668), .I0(n360[22]), .I1(n1[22]), .CO(n53669));
    SB_LUT4 add_5081_4_lut (.I0(GND_net), .I1(n19468[1]), .I2(n250_adj_4780), 
            .I3(n54631), .O(n19132[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n1[21]), .I3(n53667), 
            .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n53667), .I0(n360[21]), .I1(n1[21]), .CO(n53668));
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n1[20]), .I3(n53666), 
            .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n53666), .I0(n360[20]), .I1(n1[20]), .CO(n53667));
    SB_CARRY add_5081_4 (.CI(n54631), .I0(n19468[1]), .I1(n250_adj_4780), 
            .CO(n54632));
    SB_LUT4 LessThan_9_i24_3_lut_3_lut (.I0(setpoint[11]), .I1(setpoint[12]), 
            .I2(PWMLimit[12]), .I3(GND_net), .O(n24_adj_4925));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5081_3_lut (.I0(GND_net), .I1(n19468[0]), .I2(n177_adj_4779), 
            .I3(n54630), .O(n19132[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5081_3 (.CI(n54630), .I0(n19468[0]), .I1(n177_adj_4779), 
            .CO(n54631));
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n1[19]), .I3(n53665), 
            .O(n455[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n53665), .I0(n360[19]), .I1(n1[19]), .CO(n53666));
    SB_LUT4 add_5081_2_lut (.I0(GND_net), .I1(n35_adj_4778), .I2(n104_adj_4777), 
            .I3(GND_net), .O(n19132[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5081_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n1[18]), .I3(n53664), 
            .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n53664), .I0(n360[18]), .I1(n1[18]), .CO(n53665));
    SB_CARRY add_5081_2 (.CI(GND_net), .I0(n35_adj_4778), .I1(n104_adj_4777), 
            .CO(n54630));
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n1[17]), .I3(n53663), 
            .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n53663), .I0(n360[17]), .I1(n1[17]), .CO(n53664));
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n1[16]), .I3(n53662), 
            .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n53662), .I0(n360[16]), .I1(n1[16]), .CO(n53663));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n1[15]), .I3(n53661), 
            .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_17 (.CI(n53661), .I0(n360[15]), .I1(n1[15]), .CO(n53662));
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n1[14]), .I3(n53660), 
            .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_16 (.CI(n53660), .I0(n360[14]), .I1(n1[14]), .CO(n53661));
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n1[13]), .I3(n53659), 
            .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_15 (.CI(n53659), .I0(n360[13]), .I1(n1[13]), .CO(n53660));
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n1[12]), .I3(n53658), 
            .O(n455[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n53658), .I0(n360[12]), .I1(n1[12]), .CO(n53659));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n1[11]), .I3(n53657), 
            .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n53657), .I0(n360[11]), .I1(n1[11]), .CO(n53658));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n1[10]), .I3(n53656), 
            .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_12 (.CI(n53656), .I0(n360[10]), .I1(n1[10]), .CO(n53657));
    SB_LUT4 i51550_2_lut_4_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), .I2(PWMLimit[13]), 
            .I3(setpoint[13]), .O(n68640));
    defparam i51550_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i26_3_lut_3_lut (.I0(setpoint[13]), .I1(setpoint[17]), 
            .I2(PWMLimit[17]), .I3(GND_net), .O(n26_adj_4926));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4927));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5147_11_lut (.I0(GND_net), .I1(n20192[8]), .I2(n770_adj_4776), 
            .I3(n54241), .O(n19994[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5147_10_lut (.I0(GND_net), .I1(n20192[7]), .I2(n697_adj_4775), 
            .I3(n54240), .O(n19994[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_10 (.CI(n54240), .I0(n20192[7]), .I1(n697_adj_4775), 
            .CO(n54241));
    SB_LUT4 add_5147_9_lut (.I0(GND_net), .I1(n20192[6]), .I2(n624_adj_4773), 
            .I3(n54239), .O(n19994[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_9 (.CI(n54239), .I0(n20192[6]), .I1(n624_adj_4773), 
            .CO(n54240));
    SB_LUT4 add_5147_8_lut (.I0(GND_net), .I1(n20192[5]), .I2(n551_adj_4772), 
            .I3(n54238), .O(n19994[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_8 (.CI(n54238), .I0(n20192[5]), .I1(n551_adj_4772), 
            .CO(n54239));
    SB_LUT4 add_5147_7_lut (.I0(GND_net), .I1(n20192[4]), .I2(n478_adj_4771), 
            .I3(n54237), .O(n19994[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_7 (.CI(n54237), .I0(n20192[4]), .I1(n478_adj_4771), 
            .CO(n54238));
    SB_LUT4 add_5147_6_lut (.I0(GND_net), .I1(n20192[3]), .I2(n405_adj_4770), 
            .I3(n54236), .O(n19994[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_6 (.CI(n54236), .I0(n20192[3]), .I1(n405_adj_4770), 
            .CO(n54237));
    SB_LUT4 add_5147_5_lut (.I0(GND_net), .I1(n20192[2]), .I2(n332_adj_4769), 
            .I3(n54235), .O(n19994[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_5 (.CI(n54235), .I0(n20192[2]), .I1(n332_adj_4769), 
            .CO(n54236));
    SB_LUT4 add_5147_4_lut (.I0(GND_net), .I1(n20192[1]), .I2(n259_adj_4768), 
            .I3(n54234), .O(n19994[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_4 (.CI(n54234), .I0(n20192[1]), .I1(n259_adj_4768), 
            .CO(n54235));
    SB_LUT4 i51562_2_lut_4_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), .I2(PWMLimit[14]), 
            .I3(setpoint[14]), .O(n68652));
    defparam i51562_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5147_3_lut (.I0(GND_net), .I1(n20192[0]), .I2(n186_adj_4767), 
            .I3(n54233), .O(n19994[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_3 (.CI(n54233), .I0(n20192[0]), .I1(n186_adj_4767), 
            .CO(n54234));
    SB_LUT4 add_5147_2_lut (.I0(GND_net), .I1(n44_adj_4766), .I2(n113_adj_4765), 
            .I3(GND_net), .O(n19994[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5147_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5147_2 (.CI(GND_net), .I0(n44_adj_4766), .I1(n113_adj_4765), 
            .CO(n54233));
    SB_LUT4 LessThan_30_i23_2_lut (.I0(PWMLimit[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4928));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i43_2_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4929));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i28_3_lut_3_lut (.I0(setpoint[14]), .I1(setpoint[15]), 
            .I2(PWMLimit[15]), .I3(GND_net), .O(n28));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4939_18_lut (.I0(GND_net), .I1(n17462[15]), .I2(GND_net), 
            .I3(n54213), .O(n16743[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4939_17_lut (.I0(GND_net), .I1(n17462[14]), .I2(GND_net), 
            .I3(n54212), .O(n16743[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_17 (.CI(n54212), .I0(n17462[14]), .I1(GND_net), 
            .CO(n54213));
    SB_LUT4 add_4939_16_lut (.I0(GND_net), .I1(n17462[13]), .I2(n1114), 
            .I3(n54211), .O(n16743[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_16 (.CI(n54211), .I0(n17462[13]), .I1(n1114), .CO(n54212));
    SB_LUT4 LessThan_30_i45_2_lut (.I0(PWMLimit[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4930));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4939_15_lut (.I0(GND_net), .I1(n17462[12]), .I2(n1041), 
            .I3(n54210), .O(n16743[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_15 (.CI(n54210), .I0(n17462[12]), .I1(n1041), .CO(n54211));
    SB_LUT4 add_4939_14_lut (.I0(GND_net), .I1(n17462[11]), .I2(n968), 
            .I3(n54209), .O(n16743[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_14 (.CI(n54209), .I0(n17462[11]), .I1(n968), .CO(n54210));
    SB_LUT4 add_4939_13_lut (.I0(GND_net), .I1(n17462[10]), .I2(n895), 
            .I3(n54208), .O(n16743[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_13 (.CI(n54208), .I0(n17462[10]), .I1(n895), .CO(n54209));
    SB_LUT4 add_4939_12_lut (.I0(GND_net), .I1(n17462[9]), .I2(n822), 
            .I3(n54207), .O(n16743[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_12 (.CI(n54207), .I0(n17462[9]), .I1(n822), .CO(n54208));
    SB_LUT4 add_4939_11_lut (.I0(GND_net), .I1(n17462[8]), .I2(n749), 
            .I3(n54206), .O(n16743[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_11 (.CI(n54206), .I0(n17462[8]), .I1(n749), .CO(n54207));
    SB_LUT4 add_4939_10_lut (.I0(GND_net), .I1(n17462[7]), .I2(n676), 
            .I3(n54205), .O(n16743[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_10 (.CI(n54205), .I0(n17462[7]), .I1(n676), .CO(n54206));
    SB_LUT4 add_4939_9_lut (.I0(GND_net), .I1(n17462[6]), .I2(n603), .I3(n54204), 
            .O(n16743[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_9 (.CI(n54204), .I0(n17462[6]), .I1(n603), .CO(n54205));
    SB_LUT4 add_4939_8_lut (.I0(GND_net), .I1(n17462[5]), .I2(n530), .I3(n54203), 
            .O(n16743[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_8 (.CI(n54203), .I0(n17462[5]), .I1(n530), .CO(n54204));
    SB_LUT4 add_4939_7_lut (.I0(GND_net), .I1(n17462[4]), .I2(n457_adj_4751), 
            .I3(n54202), .O(n16743[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_7 (.CI(n54202), .I0(n17462[4]), .I1(n457_adj_4751), 
            .CO(n54203));
    SB_LUT4 add_4939_6_lut (.I0(GND_net), .I1(n17462[3]), .I2(n384_adj_4750), 
            .I3(n54201), .O(n16743[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_6 (.CI(n54201), .I0(n17462[3]), .I1(n384_adj_4750), 
            .CO(n54202));
    SB_LUT4 add_4939_5_lut (.I0(GND_net), .I1(n17462[2]), .I2(n311), .I3(n54200), 
            .O(n16743[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_5 (.CI(n54200), .I0(n17462[2]), .I1(n311), .CO(n54201));
    SB_LUT4 add_4939_4_lut (.I0(GND_net), .I1(n17462[1]), .I2(n238_adj_4749), 
            .I3(n54199), .O(n16743[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_4 (.CI(n54199), .I0(n17462[1]), .I1(n238_adj_4749), 
            .CO(n54200));
    SB_LUT4 add_4939_3_lut (.I0(GND_net), .I1(n17462[0]), .I2(n165), .I3(n54198), 
            .O(n16743[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_3 (.CI(n54198), .I0(n17462[0]), .I1(n165), .CO(n54199));
    SB_LUT4 add_4939_2_lut (.I0(GND_net), .I1(n23_adj_4748), .I2(n92), 
            .I3(GND_net), .O(n16743[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4939_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4939_2 (.CI(GND_net), .I0(n23_adj_4748), .I1(n92), .CO(n54198));
    SB_LUT4 LessThan_30_i25_2_lut (.I0(PWMLimit[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4931));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4977_17_lut (.I0(GND_net), .I1(n18055[14]), .I2(GND_net), 
            .I3(n54179), .O(n17462[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4977_16_lut (.I0(GND_net), .I1(n18055[13]), .I2(n1117), 
            .I3(n54178), .O(n17462[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_16 (.CI(n54178), .I0(n18055[13]), .I1(n1117), .CO(n54179));
    SB_LUT4 add_4977_15_lut (.I0(GND_net), .I1(n18055[12]), .I2(n1044), 
            .I3(n54177), .O(n17462[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_15 (.CI(n54177), .I0(n18055[12]), .I1(n1044), .CO(n54178));
    SB_LUT4 add_4977_14_lut (.I0(GND_net), .I1(n18055[11]), .I2(n971), 
            .I3(n54176), .O(n17462[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_14 (.CI(n54176), .I0(n18055[11]), .I1(n971), .CO(n54177));
    SB_LUT4 add_4977_13_lut (.I0(GND_net), .I1(n18055[10]), .I2(n898), 
            .I3(n54175), .O(n17462[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_13 (.CI(n54175), .I0(n18055[10]), .I1(n898), .CO(n54176));
    SB_LUT4 add_4977_12_lut (.I0(GND_net), .I1(n18055[9]), .I2(n825), 
            .I3(n54174), .O(n17462[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_12 (.CI(n54174), .I0(n18055[9]), .I1(n825), .CO(n54175));
    SB_LUT4 add_4977_11_lut (.I0(GND_net), .I1(n18055[8]), .I2(n752), 
            .I3(n54173), .O(n17462[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_11 (.CI(n54173), .I0(n18055[8]), .I1(n752), .CO(n54174));
    SB_LUT4 add_4977_10_lut (.I0(GND_net), .I1(n18055[7]), .I2(n679), 
            .I3(n54172), .O(n17462[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_10 (.CI(n54172), .I0(n18055[7]), .I1(n679), .CO(n54173));
    SB_LUT4 add_4977_9_lut (.I0(GND_net), .I1(n18055[6]), .I2(n606), .I3(n54171), 
            .O(n17462[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_9 (.CI(n54171), .I0(n18055[6]), .I1(n606), .CO(n54172));
    SB_LUT4 add_4977_8_lut (.I0(GND_net), .I1(n18055[5]), .I2(n533), .I3(n54170), 
            .O(n17462[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_8 (.CI(n54170), .I0(n18055[5]), .I1(n533), .CO(n54171));
    SB_LUT4 add_4977_7_lut (.I0(GND_net), .I1(n18055[4]), .I2(n460_adj_4716), 
            .I3(n54169), .O(n17462[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_7 (.CI(n54169), .I0(n18055[4]), .I1(n460_adj_4716), 
            .CO(n54170));
    SB_LUT4 add_4977_6_lut (.I0(GND_net), .I1(n18055[3]), .I2(n387_adj_4713), 
            .I3(n54168), .O(n17462[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_6 (.CI(n54168), .I0(n18055[3]), .I1(n387_adj_4713), 
            .CO(n54169));
    SB_LUT4 add_4977_5_lut (.I0(GND_net), .I1(n18055[2]), .I2(n314_adj_4712), 
            .I3(n54167), .O(n17462[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_5 (.CI(n54167), .I0(n18055[2]), .I1(n314_adj_4712), 
            .CO(n54168));
    SB_LUT4 add_4977_4_lut (.I0(GND_net), .I1(n18055[1]), .I2(n241_adj_4711), 
            .I3(n54166), .O(n17462[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_4 (.CI(n54166), .I0(n18055[1]), .I1(n241_adj_4711), 
            .CO(n54167));
    SB_LUT4 add_4977_3_lut (.I0(GND_net), .I1(n18055[0]), .I2(n168), .I3(n54165), 
            .O(n17462[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_3 (.CI(n54165), .I0(n18055[0]), .I1(n168), .CO(n54166));
    SB_LUT4 add_4977_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17462[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4977_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4977_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n54165));
    SB_LUT4 add_5165_10_lut (.I0(GND_net), .I1(n20352[7]), .I2(n700), 
            .I3(n54164), .O(n20192[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5165_9_lut (.I0(GND_net), .I1(n20352[6]), .I2(n627), .I3(n54163), 
            .O(n20192[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51867_4_lut (.I0(n21_adj_4555), .I1(n19_adj_4556), .I2(n17_adj_4557), 
            .I3(n9_adj_4551), .O(n68957));
    defparam i51867_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5165_9 (.CI(n54163), .I0(n20352[6]), .I1(n627), .CO(n54164));
    SB_LUT4 add_5165_8_lut (.I0(GND_net), .I1(n20352[5]), .I2(n554_adj_4704), 
            .I3(n54162), .O(n20192[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_8 (.CI(n54162), .I0(n20352[5]), .I1(n554_adj_4704), 
            .CO(n54163));
    SB_LUT4 add_5165_7_lut (.I0(GND_net), .I1(n20352[4]), .I2(n481), .I3(n54161), 
            .O(n20192[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_7 (.CI(n54161), .I0(n20352[4]), .I1(n481), .CO(n54162));
    SB_LUT4 add_5165_6_lut (.I0(GND_net), .I1(n20352[3]), .I2(n408), .I3(n54160), 
            .O(n20192[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_6 (.CI(n54160), .I0(n20352[3]), .I1(n408), .CO(n54161));
    SB_LUT4 add_5165_5_lut (.I0(GND_net), .I1(n20352[2]), .I2(n335), .I3(n54159), 
            .O(n20192[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_5 (.CI(n54159), .I0(n20352[2]), .I1(n335), .CO(n54160));
    SB_LUT4 add_5165_4_lut (.I0(GND_net), .I1(n20352[1]), .I2(n262), .I3(n54158), 
            .O(n20192[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_4 (.CI(n54158), .I0(n20352[1]), .I1(n262), .CO(n54159));
    SB_LUT4 add_5165_3_lut (.I0(GND_net), .I1(n20352[0]), .I2(n189), .I3(n54157), 
            .O(n20192[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_3 (.CI(n54157), .I0(n20352[0]), .I1(n189), .CO(n54158));
    SB_LUT4 add_5165_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n20192[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n54157));
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4922));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n54565), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4921));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n54564), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5012_16_lut (.I0(GND_net), .I1(n18536[13]), .I2(n1120), 
            .I3(n54139), .O(n18055[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5012_15_lut (.I0(GND_net), .I1(n18536[12]), .I2(n1047), 
            .I3(n54138), .O(n18055[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_14 (.CI(n54564), .I0(GND_net), .I1(counter[12]), 
            .CO(n54565));
    SB_CARRY add_5012_15 (.CI(n54138), .I0(n18536[12]), .I1(n1047), .CO(n54139));
    SB_LUT4 add_5012_14_lut (.I0(GND_net), .I1(n18536[11]), .I2(n974), 
            .I3(n54137), .O(n18055[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n54563), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_14 (.CI(n54137), .I0(n18536[11]), .I1(n974), .CO(n54138));
    SB_LUT4 add_5012_13_lut (.I0(GND_net), .I1(n18536[10]), .I2(n901), 
            .I3(n54136), .O(n18055[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_13 (.CI(n54563), .I0(GND_net), .I1(counter[11]), 
            .CO(n54564));
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4919));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5012_13 (.CI(n54136), .I0(n18536[10]), .I1(n901), .CO(n54137));
    SB_LUT4 add_5012_12_lut (.I0(GND_net), .I1(n18536[9]), .I2(n828), 
            .I3(n54135), .O(n18055[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n54562), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_12 (.CI(n54135), .I0(n18536[9]), .I1(n828), .CO(n54136));
    SB_LUT4 add_5012_11_lut (.I0(GND_net), .I1(n18536[8]), .I2(n755), 
            .I3(n54134), .O(n18055[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_12 (.CI(n54562), .I0(GND_net), .I1(counter[10]), 
            .CO(n54563));
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4918));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_944 (.I0(n20682), .I1(n6_adj_4932), .I2(\Ki[4] ), 
            .I3(n341), .O(n20623[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_944.LUT_INIT = 16'h9666;
    SB_CARRY add_5012_11 (.CI(n54134), .I0(n18536[8]), .I1(n755), .CO(n54135));
    SB_LUT4 add_5012_10_lut (.I0(GND_net), .I1(n18536[7]), .I2(n682), 
            .I3(n54133), .O(n18055[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n54561), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51849_4_lut (.I0(n27_adj_4924), .I1(n15_adj_4554), .I2(n13_adj_4553), 
            .I3(n11_adj_4552), .O(n68939));
    defparam i51849_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5012_10 (.CI(n54133), .I0(n18536[7]), .I1(n682), .CO(n54134));
    SB_LUT4 add_5012_9_lut (.I0(GND_net), .I1(n18536[6]), .I2(n609), .I3(n54132), 
            .O(n18055[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_11 (.CI(n54561), .I0(GND_net), .I1(counter[9]), 
            .CO(n54562));
    SB_CARRY add_5012_9 (.CI(n54132), .I0(n18536[6]), .I1(n609), .CO(n54133));
    SB_LUT4 add_5012_8_lut (.I0(GND_net), .I1(n18536[5]), .I2(n536_adj_4689), 
            .I3(n54131), .O(n18055[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n54560), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_8 (.CI(n54131), .I0(n18536[5]), .I1(n536_adj_4689), 
            .CO(n54132));
    SB_LUT4 add_5012_7_lut (.I0(GND_net), .I1(n18536[4]), .I2(n463_adj_4688), 
            .I3(n54130), .O(n18055[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_10 (.CI(n54560), .I0(GND_net), .I1(counter[8]), 
            .CO(n54561));
    SB_CARRY add_5012_7 (.CI(n54130), .I0(n18536[4]), .I1(n463_adj_4688), 
            .CO(n54131));
    SB_LUT4 add_5012_6_lut (.I0(GND_net), .I1(n18536[3]), .I2(n390_adj_4686), 
            .I3(n54129), .O(n18055[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n54559), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_6 (.CI(n54129), .I0(n18536[3]), .I1(n390_adj_4686), 
            .CO(n54130));
    SB_LUT4 add_5012_5_lut (.I0(GND_net), .I1(n18536[2]), .I2(n317_adj_4685), 
            .I3(n54128), .O(n18055[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_9 (.CI(n54559), .I0(GND_net), .I1(counter[7]), 
            .CO(n54560));
    SB_CARRY add_5012_5 (.CI(n54128), .I0(n18536[2]), .I1(n317_adj_4685), 
            .CO(n54129));
    SB_LUT4 add_5012_4_lut (.I0(GND_net), .I1(n18536[1]), .I2(n244_adj_4684), 
            .I3(n54127), .O(n18055[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n54558), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4923), 
            .I3(GND_net), .O(n12_adj_4933));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5012_4 (.CI(n54127), .I0(n18536[1]), .I1(n244_adj_4684), 
            .CO(n54128));
    SB_LUT4 add_5012_3_lut (.I0(GND_net), .I1(n18536[0]), .I2(n171), .I3(n54126), 
            .O(n18055[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_8 (.CI(n54558), .I0(GND_net), .I1(counter[6]), 
            .CO(n54559));
    SB_CARRY add_5012_3 (.CI(n54126), .I0(n18536[0]), .I1(n171), .CO(n54127));
    SB_LUT4 add_5012_2_lut (.I0(GND_net), .I1(n29_adj_4683), .I2(n98), 
            .I3(GND_net), .O(n18055[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5012_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n54557), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5012_2 (.CI(GND_net), .I0(n29_adj_4683), .I1(n98), .CO(n54126));
    SB_LUT4 add_5043_15_lut (.I0(GND_net), .I1(n18967[12]), .I2(n1050), 
            .I3(n54125), .O(n18536[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_7 (.CI(n54557), .I0(GND_net), .I1(counter[5]), 
            .CO(n54558));
    SB_LUT4 add_5043_14_lut (.I0(GND_net), .I1(n18967[11]), .I2(n977), 
            .I3(n54124), .O(n18536[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_14 (.CI(n54124), .I0(n18967[11]), .I1(n977), .CO(n54125));
    SB_LUT4 counter_2045_2046_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n54556), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_13_lut (.I0(GND_net), .I1(n18967[10]), .I2(n904), 
            .I3(n54123), .O(n18536[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_13 (.CI(n54123), .I0(n18967[10]), .I1(n904), .CO(n54124));
    SB_CARRY counter_2045_2046_add_4_6 (.CI(n54556), .I0(GND_net), .I1(counter[4]), 
            .CO(n54557));
    SB_LUT4 add_5043_12_lut (.I0(GND_net), .I1(n18967[9]), .I2(n831), 
            .I3(n54122), .O(n18536[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_12 (.CI(n54122), .I0(n18967[9]), .I1(n831), .CO(n54123));
    SB_LUT4 counter_2045_2046_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n54555), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_11_lut (.I0(GND_net), .I1(n18967[8]), .I2(n758), 
            .I3(n54121), .O(n18536[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_11 (.CI(n54121), .I0(n18967[8]), .I1(n758), .CO(n54122));
    SB_CARRY counter_2045_2046_add_4_5 (.CI(n54555), .I0(GND_net), .I1(counter[3]), 
            .CO(n54556));
    SB_LUT4 add_5043_10_lut (.I0(GND_net), .I1(n18967[7]), .I2(n685), 
            .I3(n54120), .O(n18536[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_10 (.CI(n54120), .I0(n18967[7]), .I1(n685), .CO(n54121));
    SB_LUT4 counter_2045_2046_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n54554), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_9_lut (.I0(GND_net), .I1(n18967[6]), .I2(n612), .I3(n54119), 
            .O(n18536[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_9 (.CI(n54119), .I0(n18967[6]), .I1(n612), .CO(n54120));
    SB_CARRY counter_2045_2046_add_4_4 (.CI(n54554), .I0(GND_net), .I1(counter[2]), 
            .CO(n54555));
    SB_LUT4 add_5043_8_lut (.I0(GND_net), .I1(n18967[5]), .I2(n539_adj_4674), 
            .I3(n54118), .O(n18536[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_8 (.CI(n54118), .I0(n18967[5]), .I1(n539_adj_4674), 
            .CO(n54119));
    SB_LUT4 counter_2045_2046_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n54553), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_7_lut (.I0(GND_net), .I1(n18967[4]), .I2(n466_adj_4670), 
            .I3(n54117), .O(n18536[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_7 (.CI(n54117), .I0(n18967[4]), .I1(n466_adj_4670), 
            .CO(n54118));
    SB_CARRY counter_2045_2046_add_4_3 (.CI(n54553), .I0(GND_net), .I1(counter[1]), 
            .CO(n54554));
    SB_LUT4 add_5043_6_lut (.I0(GND_net), .I1(n18967[3]), .I2(n393_adj_4668), 
            .I3(n54116), .O(n18536[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_6 (.CI(n54116), .I0(n18967[3]), .I1(n393_adj_4668), 
            .CO(n54117));
    SB_LUT4 counter_2045_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5043_5_lut (.I0(GND_net), .I1(n18967[2]), .I2(n320_adj_4667), 
            .I3(n54115), .O(n18536[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_5 (.CI(n54115), .I0(n18967[2]), .I1(n320_adj_4667), 
            .CO(n54116));
    SB_CARRY counter_2045_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n54553));
    SB_LUT4 i1_4_lut_adj_945 (.I0(n20738[0]), .I1(n53302), .I2(\Ki[2] ), 
            .I3(n339), .O(n20719));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h9666;
    SB_LUT4 add_5043_4_lut (.I0(GND_net), .I1(n18967[1]), .I2(n247_adj_4662), 
            .I3(n54114), .O(n18536[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_4 (.CI(n54114), .I0(n18967[1]), .I1(n247_adj_4662), 
            .CO(n54115));
    SB_LUT4 add_5043_3_lut (.I0(GND_net), .I1(n18967[0]), .I2(n174), .I3(n54113), 
            .O(n18536[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_3 (.CI(n54113), .I0(n18967[0]), .I1(n174), .CO(n54114));
    SB_LUT4 add_5043_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18536[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5043_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5043_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n54113));
    SB_LUT4 mult_24_i42_2_lut (.I0(\Ki[0] ), .I1(n339), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4934));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5181_9_lut (.I0(GND_net), .I1(n20478[6]), .I2(n630), .I3(n54096), 
            .O(n20352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5181_8_lut (.I0(GND_net), .I1(n20478[5]), .I2(n557_adj_4625), 
            .I3(n54095), .O(n20352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_8 (.CI(n54095), .I0(n20478[5]), .I1(n557_adj_4625), 
            .CO(n54096));
    SB_LUT4 add_5181_7_lut (.I0(GND_net), .I1(n20478[4]), .I2(n484), .I3(n54094), 
            .O(n20352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_7 (.CI(n54094), .I0(n20478[4]), .I1(n484), .CO(n54095));
    SB_LUT4 add_5181_6_lut (.I0(GND_net), .I1(n20478[3]), .I2(n411), .I3(n54093), 
            .O(n20352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_6 (.CI(n54093), .I0(n20478[3]), .I1(n411), .CO(n54094));
    SB_LUT4 LessThan_30_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4553), 
            .I3(GND_net), .O(n10_adj_4935));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5181_5_lut (.I0(GND_net), .I1(n20478[2]), .I2(n338_adj_4617), 
            .I3(n54092), .O(n20352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_5 (.CI(n54092), .I0(n20478[2]), .I1(n338_adj_4617), 
            .CO(n54093));
    SB_LUT4 add_5181_4_lut (.I0(GND_net), .I1(n20478[1]), .I2(n265), .I3(n54091), 
            .O(n20352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_4 (.CI(n54091), .I0(n20478[1]), .I1(n265), .CO(n54092));
    SB_LUT4 add_5181_3_lut (.I0(GND_net), .I1(n20478[0]), .I2(n192), .I3(n54090), 
            .O(n20352[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_3 (.CI(n54090), .I0(n20478[0]), .I1(n192), .CO(n54091));
    SB_LUT4 add_5181_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20352[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5181_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5181_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n54090));
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4917));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_14_lut (.I0(GND_net), .I1(n19328[11]), .I2(n980), 
            .I3(n54089), .O(n18967[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_13_lut (.I0(GND_net), .I1(n19328[10]), .I2(n907), 
            .I3(n54088), .O(n18967[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_946 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n337), .I3(n336), 
            .O(n64571));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_946.LUT_INIT = 16'h93a0;
    SB_CARRY add_5070_13 (.CI(n54088), .I0(n19328[10]), .I1(n907), .CO(n54089));
    SB_LUT4 add_5070_12_lut (.I0(GND_net), .I1(n19328[9]), .I2(n834), 
            .I3(n54087), .O(n18967[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_12 (.CI(n54087), .I0(n19328[9]), .I1(n834), .CO(n54088));
    SB_LUT4 add_5070_11_lut (.I0(GND_net), .I1(n19328[8]), .I2(n761), 
            .I3(n54086), .O(n18967[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_11 (.CI(n54086), .I0(n19328[8]), .I1(n761), .CO(n54087));
    SB_LUT4 add_5070_10_lut (.I0(GND_net), .I1(n19328[7]), .I2(n688), 
            .I3(n54085), .O(n18967[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_10 (.CI(n54085), .I0(n19328[7]), .I1(n688), .CO(n54086));
    SB_LUT4 add_5070_9_lut (.I0(GND_net), .I1(n19328[6]), .I2(n615), .I3(n54084), 
            .O(n18967[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_9 (.CI(n54084), .I0(n19328[6]), .I1(n615), .CO(n54085));
    SB_LUT4 add_5070_8_lut (.I0(GND_net), .I1(n19328[5]), .I2(n542_adj_4599), 
            .I3(n54083), .O(n18967[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_8 (.CI(n54083), .I0(n19328[5]), .I1(n542_adj_4599), 
            .CO(n54084));
    SB_LUT4 add_5070_7_lut (.I0(GND_net), .I1(n19328[4]), .I2(n469_adj_4598), 
            .I3(n54082), .O(n18967[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_7 (.CI(n54082), .I0(n19328[4]), .I1(n469_adj_4598), 
            .CO(n54083));
    SB_LUT4 add_5070_6_lut (.I0(GND_net), .I1(n19328[3]), .I2(n396_adj_4594), 
            .I3(n54081), .O(n18967[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_6 (.CI(n54081), .I0(n19328[3]), .I1(n396_adj_4594), 
            .CO(n54082));
    SB_LUT4 add_5070_5_lut (.I0(GND_net), .I1(n19328[2]), .I2(n323_adj_4593), 
            .I3(n54080), .O(n18967[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_5 (.CI(n54080), .I0(n19328[2]), .I1(n323_adj_4593), 
            .CO(n54081));
    SB_LUT4 add_5070_4_lut (.I0(GND_net), .I1(n19328[1]), .I2(n250_adj_4591), 
            .I3(n54079), .O(n18967[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_4 (.CI(n54079), .I0(n19328[1]), .I1(n250_adj_4591), 
            .CO(n54080));
    SB_LUT4 add_5070_3_lut (.I0(GND_net), .I1(n19328[0]), .I2(n177), .I3(n54078), 
            .O(n18967[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_947 (.I0(\Ki[5] ), .I1(n34395), .I2(n341), .I3(\Ki[4] ), 
            .O(n64575));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'h6ca0;
    SB_CARRY add_5070_3 (.CI(n54078), .I0(n19328[0]), .I1(n177), .CO(n54079));
    SB_LUT4 add_5070_2_lut (.I0(GND_net), .I1(n35_adj_4588), .I2(n104), 
            .I3(GND_net), .O(n18967[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_2 (.CI(GND_net), .I0(n35_adj_4588), .I1(n104), .CO(n54078));
    SB_LUT4 add_5095_13_lut (.I0(GND_net), .I1(n19637[10]), .I2(n910_adj_4584), 
            .I3(n54077), .O(n19328[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5095_12_lut (.I0(GND_net), .I1(n19637[9]), .I2(n837_adj_4582), 
            .I3(n54076), .O(n19328[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5095_12 (.CI(n54076), .I0(n19637[9]), .I1(n837_adj_4582), 
            .CO(n54077));
    SB_LUT4 add_5095_11_lut (.I0(GND_net), .I1(n19637[8]), .I2(n764_adj_4579), 
            .I3(n54075), .O(n19328[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5095_11 (.CI(n54075), .I0(n19637[8]), .I1(n764_adj_4579), 
            .CO(n54076));
    SB_LUT4 add_5095_10_lut (.I0(GND_net), .I1(n19637[7]), .I2(n691_adj_4578), 
            .I3(n54074), .O(n19328[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5095_10 (.CI(n54074), .I0(n19637[7]), .I1(n691_adj_4578), 
            .CO(n54075));
    SB_LUT4 add_5095_9_lut (.I0(GND_net), .I1(n19637[6]), .I2(n618_adj_4577), 
            .I3(n54073), .O(n19328[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5095_9 (.CI(n54073), .I0(n19637[6]), .I1(n618_adj_4577), 
            .CO(n54074));
    SB_LUT4 i1_4_lut_adj_948 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(n339), .I3(n338), 
            .O(n64573));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n64573), .I1(n53272), .I2(n64575), .I3(n64571), 
            .O(n64581));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i37572_4_lut (.I0(n20738[0]), .I1(\Ki[2] ), .I2(n53302), .I3(n339), 
            .O(n4_adj_4936));   // verilog/motorControl.v(61[29:40])
    defparam i37572_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i37710_4_lut (.I0(n20682), .I1(\Ki[4] ), .I2(n6_adj_4932), 
            .I3(n341), .O(n8_adj_4937));   // verilog/motorControl.v(61[29:40])
    defparam i37710_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n12_adj_4933), .I1(n455[17]), .I2(n35_adj_4861), 
            .I3(GND_net), .O(n30_adj_4938));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 reduce_or_1110_i1_2_lut_3_lut_4_lut (.I0(n39142), .I1(n54838), 
            .I2(n508), .I3(n7063), .O(n5083));
    defparam reduce_or_1110_i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff80;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n6), .I1(n8_adj_4937), .I2(n4_adj_4936), 
            .I3(n64581), .O(n62699));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i52847_4_lut (.I0(n13_adj_4553), .I1(n11_adj_4552), .I2(n9_adj_4551), 
            .I3(n68983), .O(n69937));
    defparam i52847_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52841_4_lut (.I0(n19_adj_4556), .I1(n17_adj_4557), .I2(n15_adj_4554), 
            .I3(n69937), .O(n69931));
    defparam i52841_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4916));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54086_4_lut (.I0(n25_adj_4931), .I1(n23_adj_4928), .I2(n21_adj_4555), 
            .I3(n69931), .O(n71176));
    defparam i54086_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4915));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4914));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4913));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4912));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4911));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4910));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4909));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4908));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4906));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4905));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4903));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4902));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4900));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4899));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4897));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4896));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4895));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4893));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4889));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4888));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4887));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4885));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4884));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4883));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4882));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53401_4_lut (.I0(n31_adj_4920), .I1(n29_adj_4927), .I2(n27_adj_4924), 
            .I3(n71176), .O(n70491));
    defparam i53401_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4879));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4878));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4876));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4875));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4874));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4873));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4872));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4871));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4870));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4869));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54274_4_lut (.I0(n37_adj_4846), .I1(n35_adj_4861), .I2(n33_adj_4923), 
            .I3(n70491), .O(n71364));
    defparam i54274_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4929), 
            .I3(GND_net), .O(n16_adj_4940));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4866));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4865));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53826_3_lut (.I0(n6_adj_4941), .I1(n455[10]), .I2(n21_adj_4555), 
            .I3(GND_net), .O(n70916));   // verilog/motorControl.v(63[16:31])
    defparam i53826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4863));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53827_3_lut (.I0(n70916), .I1(n455[11]), .I2(n23_adj_4928), 
            .I3(GND_net), .O(n70917));   // verilog/motorControl.v(63[16:31])
    defparam i53827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4860));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4854));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4853));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4852));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4849));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4844));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4841));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4839));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4836));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4557), 
            .I3(GND_net), .O(n8_adj_4942));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4833));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_30_i24_3_lut (.I0(n16_adj_4940), .I1(n455[22]), .I2(n45_adj_4930), 
            .I3(GND_net), .O(n24_adj_4943));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4826));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4823));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47928_2_lut (.I0(counter[11]), .I1(counter[13]), .I2(GND_net), 
            .I3(GND_net), .O(n65002));
    defparam i47928_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(counter[8]), .I1(counter[0]), .I2(counter[2]), 
            .I3(counter[3]), .O(n23_adj_4944));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5003[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23717_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n39485));   // verilog/motorControl.v(61[20:40])
    defparam i23717_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4817));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4816));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4815));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4812));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4810));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut (.I0(counter[1]), .I1(counter[6]), .I2(counter[10]), 
            .I3(counter[5]), .O(n22_adj_4945));
    defparam i8_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4809));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut (.I0(n23_adj_4944), .I1(counter[4]), .I2(n65002), 
            .I3(counter[9]), .O(n26_adj_4946));
    defparam i12_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51773_4_lut (.I0(n43_adj_4929), .I1(n25_adj_4931), .I2(n23_adj_4928), 
            .I3(n68957), .O(n68863));
    defparam i51773_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4807));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4804));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54561_4_lut (.I0(counter[7]), .I1(n26_adj_4946), .I2(n22_adj_4945), 
            .I3(counter[12]), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i54561_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4802));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54542_4_lut (.I0(\encoder1_position_scaled[0] ), .I1(n15), 
            .I2(n68243), .I3(n15_adj_2), .O(motor_state[0]));   // verilog/motorControl.v(53[17:33])
    defparam i54542_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4799));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4782));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4774));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n353), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4763));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4762));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4760));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4759));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4757));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4755));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51978_2_lut_4_lut (.I0(deadband[21]), .I1(n455[21]), .I2(deadband[9]), 
            .I3(n455[9]), .O(n69068));
    defparam i51978_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4754));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53694_4_lut (.I0(n24_adj_4943), .I1(n8_adj_4942), .I2(n45_adj_4930), 
            .I3(n68861), .O(n70784));   // verilog/motorControl.v(63[16:31])
    defparam i53694_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4745));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4744));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4741));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n344), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4739));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4736));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4735));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52604_3_lut (.I0(n70917), .I1(n455[12]), .I2(n25_adj_4931), 
            .I3(GND_net), .O(n69694));   // verilog/motorControl.v(63[16:31])
    defparam i52604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4733));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4732));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4729));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4728));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4727));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4725));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5002[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4722));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4721));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4720));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_4949));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4719));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4718));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4717));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n207[23]), .I1(\Kp[2] ), .I2(n4_adj_4950), 
            .I3(n207[22]), .O(n64619));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4715));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_952 (.I0(n207[22]), .I1(n20722[1]), .I2(n4_adj_4951), 
            .I3(\Kp[3] ), .O(n20644[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'hc66c;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4714));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_4952));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_953 (.I0(n20722[1]), .I1(n6_adj_4953), .I2(n347_adj_4952), 
            .I3(n61219), .O(n20644[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i53824_3_lut (.I0(n4_adj_4949), .I1(n455[13]), .I2(n27_adj_4924), 
            .I3(GND_net), .O(n70914));   // verilog/motorControl.v(63[16:31])
    defparam i53824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4710));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(n64615), .I1(n207[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4951));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37782_4_lut (.I0(n20722[1]), .I1(\Kp[3] ), .I2(n4_adj_4951), 
            .I3(n207[22]), .O(n6_adj_4953));   // verilog/motorControl.v(61[20:26])
    defparam i37782_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 mult_23_i46_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_4954));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\Kp[1] ), .I1(\Kp[2] ), .I2(\Kp[0] ), .I3(GND_net), 
            .O(n64615));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i48012_3_lut (.I0(n207[23]), .I1(n64615), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n61219));   // verilog/motorControl.v(61[20:26])
    defparam i48012_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i37591_3_lut (.I0(n207[23]), .I1(n53327), .I2(n54844), .I3(GND_net), 
            .O(n20722[1]));   // verilog/motorControl.v(61[20:26])
    defparam i37591_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\Kp[1] ), .I1(\Kp[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4950));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n54844), 
            .I3(n207[22]), .O(n64605));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_581_2_lut (.I0(n20722[1]), .I1(n61219), .I2(GND_net), 
            .I3(GND_net), .O(n73003));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_581_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_956 (.I0(n53327), .I1(n64605), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n64609));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h9666;
    SB_LUT4 i37790_4_lut (.I0(n73003), .I1(\Kp[4] ), .I2(n6_adj_4953), 
            .I3(n207[22]), .O(n8_adj_4955));   // verilog/motorControl.v(61[20:26])
    defparam i37790_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i37743_4_lut (.I0(n20722[1]), .I1(\Kp[3] ), .I2(n64615), .I3(n207[23]), 
            .O(n6_adj_4956));   // verilog/motorControl.v(61[20:26])
    defparam i37743_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n6_adj_4956), .I1(n8_adj_4955), .I2(n64609), 
            .I3(n61219), .O(n62402));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4709));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4708));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4707));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4706));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4705));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n354), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4703));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4701));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4699));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4698));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4697));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52015_2_lut_4_lut (.I0(deadband[16]), .I1(n455[16]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n69105));
    defparam i52015_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53825_3_lut (.I0(n70914), .I1(n455[14]), .I2(n29_adj_4927), 
            .I3(GND_net), .O(n70915));   // verilog/motorControl.v(63[16:31])
    defparam i53825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4695));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5095_8_lut (.I0(GND_net), .I1(n19637[5]), .I2(n545_adj_4576), 
            .I3(n54072), .O(n19328[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51822_4_lut (.I0(n33_adj_4923), .I1(n31_adj_4920), .I2(n29_adj_4927), 
            .I3(n68939), .O(n68912));
    defparam i51822_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4693));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4692));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53970_4_lut (.I0(n30_adj_4938), .I1(n10_adj_4935), .I2(n35_adj_4861), 
            .I3(n68903), .O(n71060));   // verilog/motorControl.v(63[16:31])
    defparam i53970_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4690));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4687));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5095_8 (.CI(n54072), .I0(n19637[5]), .I1(n545_adj_4576), 
            .CO(n54073));
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4682));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5095_7_lut (.I0(GND_net), .I1(n19637[4]), .I2(n472_adj_4575), 
            .I3(n54071), .O(n19328[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52606_3_lut (.I0(n70915), .I1(n455[15]), .I2(n31_adj_4920), 
            .I3(GND_net), .O(n69696));   // verilog/motorControl.v(63[16:31])
    defparam i52606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4680));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4666));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4679));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4678));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4677));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4676));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4675));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n345), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4665));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4663));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54355_4_lut (.I0(n69696), .I1(n71060), .I2(n35_adj_4861), 
            .I3(n68912), .O(n71445));   // verilog/motorControl.v(63[16:31])
    defparam i54355_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54356_3_lut (.I0(n71445), .I1(n455[18]), .I2(n37_adj_4846), 
            .I3(GND_net), .O(n71446));   // verilog/motorControl.v(63[16:31])
    defparam i54356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4661));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5095_7 (.CI(n54071), .I0(n19637[4]), .I1(n472_adj_4575), 
            .CO(n54072));
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4672));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n342), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4671));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54273_3_lut (.I0(n71446), .I1(n455[19]), .I2(n39_adj_4798), 
            .I3(GND_net), .O(n71363));   // verilog/motorControl.v(63[16:31])
    defparam i54273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5095_6_lut (.I0(GND_net), .I1(n19637[3]), .I2(n399_adj_4574), 
            .I3(n54070), .O(n19328[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5095_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51780_4_lut (.I0(n43_adj_4929), .I1(n41_adj_4793), .I2(n39_adj_4798), 
            .I3(n71364), .O(n68870));
    defparam i51780_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5095_6 (.CI(n54070), .I0(n19637[3]), .I1(n399_adj_4574), 
            .CO(n54071));
    SB_LUT4 i53982_4_lut (.I0(n69694), .I1(n70784), .I2(n45_adj_4930), 
            .I3(n68863), .O(n71072));   // verilog/motorControl.v(63[16:31])
    defparam i53982_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4660));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4669));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4659));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4657));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4656));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4655));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4654));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4653));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n343), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4652));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4651));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52612_3_lut (.I0(n71363), .I1(n455[20]), .I2(n41_adj_4793), 
            .I3(GND_net), .O(n69702));   // verilog/motorControl.v(63[16:31])
    defparam i52612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4650));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54245_4_lut (.I0(n69702), .I1(n71072), .I2(n45_adj_4930), 
            .I3(n68870), .O(n71335));   // verilog/motorControl.v(63[16:31])
    defparam i54245_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n310[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4649));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i13_3_lut (.I0(n310[12]), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n347));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4648));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i26_2_lut (.I0(\Ki[0] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4438));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54246_3_lut (.I0(n71335), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(GND_net), .O(n508));   // verilog/motorControl.v(63[16:31])
    defparam i54246_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4647));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4646));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4645));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n355), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4644));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4643));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4642));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i45_2_lut (.I0(deadband[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4957));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4958));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i43_2_lut (.I0(deadband[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4959));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4641));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i39_2_lut (.I0(deadband[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4960));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4640));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(deadband[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4961));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4639));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4638));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4637));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4636));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4635));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4634));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i37_2_lut (.I0(deadband[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4962));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4633));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4632));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(deadband[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4963));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37810_2_lut (.I0(n22), .I1(control_update), .I2(GND_net), 
            .I3(GND_net), .O(n54838));
    defparam i37810_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4631));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51972_4_lut (.I0(n455[6]), .I1(n455[5]), .I2(n36[6]), .I3(n36[5]), 
            .O(n69062));
    defparam i51972_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52925_3_lut (.I0(n455[7]), .I1(n69062), .I2(n36[7]), .I3(GND_net), 
            .O(n70015));
    defparam i52925_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4630));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i27_rep_102_2_lut (.I0(n455[13]), .I1(n36[13]), 
            .I2(GND_net), .I3(GND_net), .O(n72524));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_rep_102_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4629));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52897_4_lut (.I0(n455[14]), .I1(n72524), .I2(n36[14]), .I3(n70015), 
            .O(n69987));
    defparam i52897_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i31_rep_97_2_lut (.I0(n455[15]), .I1(n36[15]), .I2(GND_net), 
            .I3(GND_net), .O(n72519));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_rep_97_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n356), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n356), .I2(GND_net), .I3(GND_net), 
            .O(n11_adj_4628));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51964_4_lut (.I0(n455[8]), .I1(n455[4]), .I2(n36[8]), .I3(n36[4]), 
            .O(n69054));
    defparam i51964_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i52917_3_lut (.I0(n455[9]), .I1(n69054), .I2(n36[9]), .I3(GND_net), 
            .O(n70007));
    defparam i52917_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4627));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i21_rep_117_2_lut (.I0(n455[10]), .I1(n36[10]), 
            .I2(GND_net), .I3(GND_net), .O(n72539));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_rep_117_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52911_4_lut (.I0(n455[11]), .I1(n72539), .I2(n36[11]), .I3(n70007), 
            .O(n70001));
    defparam i52911_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4626));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4624));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37590_2_lut_3_lut (.I0(\Kp[1] ), .I1(\Kp[0] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n54844));   // verilog/motorControl.v(61[20:26])
    defparam i37590_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 LessThan_28_i25_rep_112_2_lut (.I0(n455[12]), .I1(n36[12]), 
            .I2(GND_net), .I3(GND_net), .O(n72534));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_rep_112_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37584_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n53327));   // verilog/motorControl.v(61[20:26])
    defparam i37584_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n36[9]), .I1(n36[21]), .I2(n455[21]), 
            .I3(GND_net), .O(n16_adj_4964));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4623));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4620));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4619));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4616));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4614));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4613));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9971_bdd_4_lut_54852 (.I0(n9971), .I1(n68372), .I2(setpoint[17]), 
            .I3(n4743), .O(n71963));
    defparam n9971_bdd_4_lut_54852.LUT_INIT = 16'he4aa;
    SB_LUT4 i51895_4_lut (.I0(n455[21]), .I1(n455[9]), .I2(n36[21]), .I3(n36[9]), 
            .O(n68985));
    defparam i51895_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4611));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4610));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n36[4]), .I1(n36[8]), .I2(n455[8]), 
            .I3(GND_net), .O(n8_adj_4965));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4609));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4608));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4607));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51771_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(PWMLimit[9]), 
            .I3(n455[9]), .O(n68861));
    defparam i51771_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n357), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4605));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4604));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71963_bdd_4_lut (.I0(n71963), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4743), .O(n71966));
    defparam n71963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4603));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4602));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i24_3_lut (.I0(n16_adj_4964), .I1(n36[22]), .I2(n455[22]), 
            .I3(GND_net), .O(n24_adj_4966));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4601));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4600));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4596));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4595));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4592));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4590));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4589));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51976_4_lut (.I0(n455[3]), .I1(n455[2]), .I2(n36[3]), .I3(n36[2]), 
            .O(n69066));
    defparam i51976_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4587));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4586));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i9_rep_110_2_lut (.I0(n455[4]), .I1(n36[4]), .I2(GND_net), 
            .I3(GND_net), .O(n72532));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_rep_110_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4510));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4583));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51974_4_lut (.I0(n455[5]), .I1(n72532), .I2(n36[5]), .I3(n69066), 
            .O(n69064));
    defparam i51974_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4581));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4508));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4507));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4580));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n357), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4572));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i13_rep_138_2_lut (.I0(n455[6]), .I1(n36[6]), .I2(GND_net), 
            .I3(GND_net), .O(n72560));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_rep_138_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53469_4_lut (.I0(n455[7]), .I1(n72560), .I2(n36[7]), .I3(n69064), 
            .O(n70559));
    defparam i53469_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n358), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4571));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51711_2_lut (.I0(PWMLimit[11]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68368));
    defparam i51711_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n346), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4505));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51777_2_lut (.I0(PWMLimit[18]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68388));
    defparam i51777_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37606_2_lut_4_lut (.I0(\Ki[0] ), .I1(n339), .I2(n34395), 
            .I3(\Ki[1] ), .O(n20680[0]));   // verilog/motorControl.v(61[29:40])
    defparam i37606_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i51813_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(PWMLimit[7]), 
            .I3(n455[7]), .O(n68903));
    defparam i51813_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_28_i17_rep_135_2_lut (.I0(n455[8]), .I1(n36[8]), .I2(GND_net), 
            .I3(GND_net), .O(n72557));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_rep_135_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52919_4_lut (.I0(n455[9]), .I1(n72557), .I2(n36[9]), .I3(n70559), 
            .O(n70009));
    defparam i52919_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4499));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51776_2_lut (.I0(PWMLimit[19]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68389));
    defparam i51776_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53880_4_lut (.I0(n455[11]), .I1(n72539), .I2(n36[11]), .I3(n70009), 
            .O(n70970));
    defparam i53880_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51946_4_lut (.I0(n455[13]), .I1(n72534), .I2(n36[13]), .I3(n70970), 
            .O(n69036));
    defparam i51946_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i29_rep_100_2_lut (.I0(n455[14]), .I1(n36[14]), 
            .I2(GND_net), .I3(GND_net), .O(n72522));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_rep_100_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53459_4_lut (.I0(n455[15]), .I1(n72522), .I2(n36[15]), .I3(n69036), 
            .O(n70549));
    defparam i53459_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i33_rep_129_2_lut (.I0(n455[16]), .I1(n36[16]), 
            .I2(GND_net), .I3(GND_net), .O(n72551));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_rep_129_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37818_2_lut_3_lut (.I0(n39142), .I1(n22), .I2(control_update), 
            .I3(GND_net), .O(n54848));
    defparam i37818_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i54102_4_lut (.I0(n455[17]), .I1(n72551), .I2(n36[17]), .I3(n70549), 
            .O(n71192));
    defparam i54102_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i37_rep_91_2_lut (.I0(n455[18]), .I1(n36[18]), .I2(GND_net), 
            .I3(GND_net), .O(n72513));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i37_rep_91_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i54373_4_lut (.I0(n455[19]), .I1(n72513), .I2(n36[19]), .I3(n71192), 
            .O(n71463));
    defparam i54373_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i41_rep_88_2_lut (.I0(n455[20]), .I1(n36[20]), .I2(GND_net), 
            .I3(GND_net), .O(n72510));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i41_rep_88_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52034_4_lut (.I0(n27_adj_4567), .I1(n15_adj_4560), .I2(n13_adj_4559), 
            .I3(n11_adj_4558), .O(n69124));
    defparam i52034_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4569), 
            .I3(GND_net), .O(n12_adj_4967));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4559), 
            .I3(GND_net), .O(n10_adj_4968));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i30_3_lut (.I0(n12_adj_4967), .I1(n455[17]), .I2(n35_adj_4963), 
            .I3(GND_net), .O(n30_adj_4969));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4428_3_lut_4_lut (.I0(n131_c), .I1(n25205), .I2(n5190), .I3(n4743), 
            .O(n9971));
    defparam i4428_3_lut_4_lut.LUT_INIT = 16'h44f4;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n131_c), .I1(n25205), .I2(n508), 
            .I3(n54848), .O(n5_adj_4461));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hf444;
    SB_LUT4 i53009_4_lut (.I0(n13_adj_4559), .I1(n11_adj_4558), .I2(n9_adj_4561), 
            .I3(n69161), .O(n70099));
    defparam i53009_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i53001_4_lut (.I0(n19_adj_4563), .I1(n17_adj_4562), .I2(n15_adj_4560), 
            .I3(n70099), .O(n70091));
    defparam i53001_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n348), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4436));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54124_4_lut (.I0(n25_adj_4566), .I1(n23_adj_4565), .I2(n21_adj_4564), 
            .I3(n70091), .O(n71214));
    defparam i54124_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53503_4_lut (.I0(n31_adj_4961), .I1(n29_adj_4568), .I2(n27_adj_4567), 
            .I3(n71214), .O(n70593));
    defparam i53503_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i54282_4_lut (.I0(n37_adj_4962), .I1(n35_adj_4963), .I2(n33_adj_4569), 
            .I3(n70593), .O(n71372));
    defparam i54282_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4959), 
            .I3(GND_net), .O(n16_adj_4970));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4562), 
            .I3(GND_net), .O(n8_adj_4971));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i24_3_lut (.I0(n16_adj_4970), .I1(n455[22]), .I2(n45_adj_4957), 
            .I3(GND_net), .O(n24_adj_4972));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51826_2_lut (.I0(PWMLimit[20]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68426));
    defparam i51826_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i37761_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4954), 
            .I3(GND_net), .O(n20644[0]));   // verilog/motorControl.v(61[20:26])
    defparam i37761_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i53840_3_lut (.I0(n6_adj_4973), .I1(n455[10]), .I2(n21_adj_4564), 
            .I3(GND_net), .O(n70930));   // verilog/motorControl.v(62[14:31])
    defparam i53840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53841_3_lut (.I0(n70930), .I1(n455[11]), .I2(n23_adj_4565), 
            .I3(GND_net), .O(n70931));   // verilog/motorControl.v(62[14:31])
    defparam i53841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52046_4_lut (.I0(n21_adj_4564), .I1(n19_adj_4563), .I2(n17_adj_4562), 
            .I3(n9_adj_4561), .O(n69136));
    defparam i52046_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51982_4_lut (.I0(n43_adj_4959), .I1(n25_adj_4566), .I2(n23_adj_4565), 
            .I3(n69136), .O(n69072));
    defparam i51982_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4954), 
            .I3(n64619), .O(n20644[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i53690_4_lut (.I0(n24_adj_4972), .I1(n8_adj_4971), .I2(n45_adj_4957), 
            .I3(n69068), .O(n70780));   // verilog/motorControl.v(62[14:31])
    defparam i53690_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52584_3_lut (.I0(n70931), .I1(n455[12]), .I2(n25_adj_4566), 
            .I3(GND_net), .O(n69674));   // verilog/motorControl.v(62[14:31])
    defparam i52584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n68301), .I1(n36[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_4974));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53830_3_lut (.I0(n4_adj_4974), .I1(n36[13]), .I2(n455[13]), 
            .I3(GND_net), .O(n70920));   // verilog/motorControl.v(62[35:55])
    defparam i53830_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53831_3_lut (.I0(n70920), .I1(n36[14]), .I2(n455[14]), .I3(GND_net), 
            .O(n70921));   // verilog/motorControl.v(62[35:55])
    defparam i53831_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37530_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(n338), .I3(\Ki[1] ), 
            .O(n20738[0]));   // verilog/motorControl.v(61[29:40])
    defparam i37530_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i37532_3_lut_4_lut (.I0(\Ki[0] ), .I1(n337), .I2(n338), .I3(\Ki[1] ), 
            .O(n53272));   // verilog/motorControl.v(61[29:40])
    defparam i37532_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n36[7]), .I1(n36[16]), .I2(n455[16]), 
            .I3(GND_net), .O(n12_adj_4975));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n359), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51927_4_lut (.I0(n455[16]), .I1(n455[7]), .I2(n36[16]), .I3(n36[7]), 
            .O(n69017));
    defparam i51927_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i37559_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n338), .I2(n339), 
            .I3(\Ki[1] ), .O(n20717[0]));   // verilog/motorControl.v(61[29:40])
    defparam i37559_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i37561_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n338), .I2(n339), 
            .I3(\Ki[1] ), .O(n53302));   // verilog/motorControl.v(61[29:40])
    defparam i37561_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_28_i35_rep_123_2_lut (.I0(n455[17]), .I1(n36[17]), 
            .I2(GND_net), .I3(GND_net), .O(n72545));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_rep_123_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n36[5]), .I1(n36[6]), .I2(n455[6]), 
            .I3(GND_net), .O(n10_adj_4976));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_4975), .I1(n36[17]), .I2(n455[17]), 
            .I3(GND_net), .O(n30_adj_4977));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37702_3_lut_4_lut (.I0(\Ki[3] ), .I1(n341), .I2(n4_adj_4978), 
            .I3(n20680[1]), .O(n6_adj_4932));   // verilog/motorControl.v(61[29:40])
    defparam i37702_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i51936_4_lut (.I0(n455[16]), .I1(n72519), .I2(n36[16]), .I3(n69987), 
            .O(n69026));
    defparam i51936_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i1_3_lut_4_lut_adj_958 (.I0(\Ki[3] ), .I1(n341), .I2(n4_adj_4978), 
            .I3(n20680[1]), .O(n20623[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_958.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_959 (.I0(\Ki[2] ), .I1(n341), .I2(n53436), 
            .I3(n20680[0]), .O(n20623[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_959.LUT_INIT = 16'h8778;
    SB_LUT4 i37694_3_lut_4_lut (.I0(\Ki[2] ), .I1(n341), .I2(n53436), 
            .I3(n20680[0]), .O(n4_adj_4978));   // verilog/motorControl.v(61[29:40])
    defparam i37694_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i54183_4_lut (.I0(n30_adj_4977), .I1(n10_adj_4976), .I2(n72545), 
            .I3(n69017), .O(n71273));   // verilog/motorControl.v(62[35:55])
    defparam i54183_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52596_3_lut (.I0(n70921), .I1(n36[15]), .I2(n455[15]), .I3(GND_net), 
            .O(n69686));   // verilog/motorControl.v(62[35:55])
    defparam i52596_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54406_4_lut (.I0(n69686), .I1(n71273), .I2(n72545), .I3(n69026), 
            .O(n71496));   // verilog/motorControl.v(62[35:55])
    defparam i54406_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54407_3_lut (.I0(n71496), .I1(n36[18]), .I2(n455[18]), .I3(GND_net), 
            .O(n71497));   // verilog/motorControl.v(62[35:55])
    defparam i54407_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54362_3_lut (.I0(n71497), .I1(n36[19]), .I2(n455[19]), .I3(GND_net), 
            .O(n71452));   // verilog/motorControl.v(62[35:55])
    defparam i54362_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i6_3_lut (.I0(n36[2]), .I1(n36[3]), .I2(n455[3]), 
            .I3(GND_net), .O(n6_adj_4979));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53832_3_lut (.I0(n6_adj_4979), .I1(n36[10]), .I2(n455[10]), 
            .I3(GND_net), .O(n70922));   // verilog/motorControl.v(62[35:55])
    defparam i53832_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_960 (.I0(n62_adj_4934), .I1(n131), .I2(n204), 
            .I3(n20717[0]), .O(n20680[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_960.LUT_INIT = 16'h8778;
    SB_LUT4 i37619_3_lut_4_lut (.I0(n62_adj_4934), .I1(n131), .I2(n204), 
            .I3(n20717[0]), .O(n4));   // verilog/motorControl.v(61[29:40])
    defparam i37619_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i53833_3_lut (.I0(n70922), .I1(n36[11]), .I2(n455[11]), .I3(GND_net), 
            .O(n70923));   // verilog/motorControl.v(62[35:55])
    defparam i53833_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51897_4_lut (.I0(n455[21]), .I1(n72534), .I2(n36[21]), .I3(n70001), 
            .O(n68987));
    defparam i51897_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i45_rep_85_2_lut (.I0(n455[22]), .I1(n36[22]), .I2(GND_net), 
            .I3(GND_net), .O(n72507));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_rep_85_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53692_4_lut (.I0(n24_adj_4966), .I1(n8_adj_4965), .I2(n72507), 
            .I3(n68985), .O(n70782));   // verilog/motorControl.v(62[35:55])
    defparam i53692_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52594_3_lut (.I0(n70923), .I1(n36[12]), .I2(n455[12]), .I3(GND_net), 
            .O(n69684));   // verilog/motorControl.v(62[35:55])
    defparam i52594_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51901_4_lut (.I0(n455[21]), .I1(n72510), .I2(n36[21]), .I3(n71463), 
            .O(n68991));
    defparam i51901_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i52073_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n69163));
    defparam i52073_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i54241_4_lut (.I0(n69684), .I1(n70782), .I2(n72507), .I3(n68987), 
            .O(n71331));   // verilog/motorControl.v(62[35:55])
    defparam i54241_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52121_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n69211));
    defparam i52121_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52602_3_lut (.I0(n71452), .I1(n36[20]), .I2(n455[20]), .I3(GND_net), 
            .O(n69692));   // verilog/motorControl.v(62[35:55])
    defparam i52602_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i54243_4_lut (.I0(n69692), .I1(n71331), .I2(n72507), .I3(n68991), 
            .O(n71333));   // verilog/motorControl.v(62[35:55])
    defparam i54243_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51767_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n68857));   // verilog/motorControl.v(65[25:41])
    defparam i51767_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4491));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51416_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n68506));   // verilog/motorControl.v(47[25:43])
    defparam i51416_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_c));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52071_3_lut_4_lut (.I0(deadband[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(deadband[2]), .O(n69161));   // verilog/motorControl.v(62[14:31])
    defparam i52071_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_4982));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_26_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4973));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i53838_3_lut (.I0(n4_adj_4982), .I1(n455[13]), .I2(n27_adj_4567), 
            .I3(GND_net), .O(n70928));   // verilog/motorControl.v(62[14:31])
    defparam i53838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n336));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51893_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(PWMLimit[2]), .O(n68983));   // verilog/motorControl.v(63[16:31])
    defparam i51893_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_30_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4941));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i53839_3_lut (.I0(n70928), .I1(n455[14]), .I2(n29_adj_4568), 
            .I3(GND_net), .O(n70929));   // verilog/motorControl.v(62[14:31])
    defparam i53839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52187_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n69277));
    defparam i52187_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52024_4_lut (.I0(n33_adj_4569), .I1(n31_adj_4961), .I2(n29_adj_4568), 
            .I3(n69124), .O(n69114));
    defparam i52024_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54181_4_lut (.I0(n30_adj_4969), .I1(n10_adj_4968), .I2(n35_adj_4963), 
            .I3(n69105), .O(n71271));   // verilog/motorControl.v(62[14:31])
    defparam i54181_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52586_3_lut (.I0(n70929), .I1(n455[15]), .I2(n31_adj_4961), 
            .I3(GND_net), .O(n69676));   // verilog/motorControl.v(62[14:31])
    defparam i52586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52236_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n69326));
    defparam i52236_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51706_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n68796));
    defparam i51706_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n9971_bdd_4_lut_54847 (.I0(n9971), .I1(n68296), .I2(setpoint[16]), 
            .I3(n4743), .O(n71891));
    defparam n9971_bdd_4_lut_54847.LUT_INIT = 16'he4aa;
    SB_LUT4 i54404_4_lut (.I0(n69676), .I1(n71271), .I2(n35_adj_4963), 
            .I3(n69114), .O(n71494));   // verilog/motorControl.v(62[14:31])
    defparam i54404_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n71891_bdd_4_lut (.I0(n71891), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4743), .O(n71894));
    defparam n71891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i54405_3_lut (.I0(n71494), .I1(n455[18]), .I2(n37_adj_4962), 
            .I3(GND_net), .O(n71495));   // verilog/motorControl.v(62[14:31])
    defparam i54405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9971_bdd_4_lut_54790 (.I0(n9971), .I1(n68343), .I2(setpoint[10]), 
            .I3(n4743), .O(n71885));
    defparam n9971_bdd_4_lut_54790.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n347), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i54364_3_lut (.I0(n71495), .I1(n455[19]), .I2(n39_adj_4960), 
            .I3(GND_net), .O(n71454));   // verilog/motorControl.v(62[14:31])
    defparam i54364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52360_2_lut (.I0(PWMLimit[0]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68482));
    defparam i52360_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n71885_bdd_4_lut (.I0(n71885), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4743), .O(n71888));
    defparam n71885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9971_bdd_4_lut_54785 (.I0(n9971), .I1(n68284), .I2(setpoint[15]), 
            .I3(n4743), .O(n71879));
    defparam n9971_bdd_4_lut_54785.LUT_INIT = 16'he4aa;
    SB_LUT4 i51986_4_lut (.I0(n43_adj_4959), .I1(n41_adj_4958), .I2(n39_adj_4960), 
            .I3(n71372), .O(n69076));
    defparam i51986_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n71879_bdd_4_lut (.I0(n71879), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4743), .O(n71882));
    defparam n71879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i51734_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n68824));
    defparam i51734_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n9971_bdd_4_lut_54780 (.I0(n9971), .I1(n68271), .I2(setpoint[14]), 
            .I3(n4743), .O(n71861));
    defparam n9971_bdd_4_lut_54780.LUT_INIT = 16'he4aa;
    SB_LUT4 i52179_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n69269));   // verilog/motorControl.v(58[23:46])
    defparam i52179_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i54237_4_lut (.I0(n69674), .I1(n70780), .I2(n45_adj_4957), 
            .I3(n69072), .O(n71327));   // verilog/motorControl.v(62[14:31])
    defparam i54237_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52592_3_lut (.I0(n71454), .I1(n455[20]), .I2(n41_adj_4958), 
            .I3(GND_net), .O(n69682));   // verilog/motorControl.v(62[14:31])
    defparam i52592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54244_3_lut (.I0(n71333), .I1(n455[23]), .I2(n47_adj_4723), 
            .I3(GND_net), .O(n71334));   // verilog/motorControl.v(62[35:55])
    defparam i54244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n71861_bdd_4_lut (.I0(n71861), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4743), .O(n71864));
    defparam n71861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i54239_4_lut (.I0(n69682), .I1(n71327), .I2(n45_adj_4957), 
            .I3(n69076), .O(n71329));   // verilog/motorControl.v(62[14:31])
    defparam i54239_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4546));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5001[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23378_4_lut (.I0(n71329), .I1(n71334), .I2(deadband[23]), 
            .I3(n455[23]), .O(n39142));
    defparam i23378_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 i51413_2_lut (.I0(PWMLimit[1]), .I1(n5083), .I2(GND_net), 
            .I3(GND_net), .O(n68483));
    defparam i51413_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52302_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n69392));
    defparam i52302_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52365_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n69455));
    defparam i52365_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_9_i43_2_lut (.I0(PWMLimit[21]), .I1(setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i39_2_lut (.I0(PWMLimit[19]), .I1(setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4984));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9971_bdd_4_lut_54767 (.I0(n9971), .I1(n68252), .I2(setpoint[13]), 
            .I3(n4743), .O(n71855));
    defparam n9971_bdd_4_lut_54767.LUT_INIT = 16'he4aa;
    SB_LUT4 LessThan_9_i41_2_lut (.I0(PWMLimit[20]), .I1(setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4985));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i17_2_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4986));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n71855_bdd_4_lut (.I0(n71855), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4743), .O(n71858));
    defparam n71855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i53317_3_lut (.I0(n4_adj_3), .I1(setpoint[2]), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n70407));   // verilog/motorControl.v(45[16:33])
    defparam i53317_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i53318_3_lut (.I0(n70407), .I1(setpoint[3]), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(45[16:33])
    defparam i53318_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_9_i16_3_lut (.I0(n14), .I1(setpoint[8]), .I2(n17_adj_4986), 
            .I3(GND_net), .O(n16_adj_4989));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53319_4_lut (.I0(n16_adj_4989), .I1(n12), .I2(n17_adj_4986), 
            .I3(n68680), .O(n70409));   // verilog/motorControl.v(45[16:33])
    defparam i53319_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 n9971_bdd_4_lut_54762 (.I0(n9971), .I1(n68266), .I2(setpoint[9]), 
            .I3(n4743), .O(n71843));
    defparam n9971_bdd_4_lut_54762.LUT_INIT = 16'he4aa;
    SB_LUT4 i53320_3_lut (.I0(n70409), .I1(setpoint[9]), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(45[16:33])
    defparam i53320_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n71843_bdd_4_lut (.I0(n71843), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4743), .O(n71846));
    defparam n71843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_9_i33_2_lut (.I0(PWMLimit[16]), .I1(setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4992));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i35_2_lut (.I0(PWMLimit[17]), .I1(setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4993));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i25_2_lut (.I0(PWMLimit[12]), .I1(setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4994));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4995));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4996));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4997));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52290_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n69380));   // verilog/motorControl.v(56[14:36])
    defparam i52290_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_adj_4506));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51566_4_lut (.I0(n29_adj_4996), .I1(n27_adj_4995), .I2(n25_adj_4994), 
            .I3(n23_adj_4997), .O(n68656));
    defparam i51566_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51554_4_lut (.I0(n35_adj_4993), .I1(n33_adj_4992), .I2(n31), 
            .I3(n68656), .O(n68644));
    defparam i51554_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_9_i30_3_lut (.I0(n28), .I1(setpoint[16]), .I2(n33_adj_4992), 
            .I3(GND_net), .O(n30_adj_4999));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_9_i34_3_lut (.I0(n26_adj_4926), .I1(setpoint[18]), 
            .I2(n37), .I3(GND_net), .O(n34));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54309_4_lut (.I0(n34), .I1(n24_adj_4925), .I2(n37), .I3(n68640), 
            .O(n71399));   // verilog/motorControl.v(45[16:33])
    defparam i54309_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i54310_3_lut (.I0(n71399), .I1(setpoint[19]), .I2(n39_adj_4984), 
            .I3(GND_net), .O(n71400));   // verilog/motorControl.v(45[16:33])
    defparam i54310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54220_3_lut (.I0(n71400), .I1(setpoint[20]), .I2(n41_adj_4985), 
            .I3(GND_net), .O(n71310));   // verilog/motorControl.v(45[16:33])
    defparam i54220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53651_4_lut (.I0(n41_adj_4985), .I1(n39_adj_4984), .I2(n37), 
            .I3(n68644), .O(n70741));
    defparam i53651_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53718_4_lut (.I0(n30_adj_4999), .I1(n34791), .I2(n33_adj_4992), 
            .I3(n68652), .O(n70808));   // verilog/motorControl.v(45[16:33])
    defparam i53718_4_lut.LUT_INIT = 16'haaac;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (GND_net, \pwm_counter[16] , \pwm_counter[19] , \pwm_counter[15] , 
            \pwm_counter[22] , \pwm_counter[21] , \pwm_counter[20] , n2881, 
            pwm_out, clk32MHz, pwm_setpoint, n31, n33, n45, n43, 
            VCC_net, n39, n41, reset, \data_in_frame[10][7] , \rx_data[7] , 
            n60771, n29190, \data_in_frame[10][6] , n25647, n25732, 
            n60896) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \pwm_counter[16] ;
    output \pwm_counter[19] ;
    output \pwm_counter[15] ;
    output \pwm_counter[22] ;
    output \pwm_counter[21] ;
    output \pwm_counter[20] ;
    input n2881;
    output pwm_out;
    input clk32MHz;
    input [23:0]pwm_setpoint;
    input n31;
    input n33;
    input n45;
    input n43;
    input VCC_net;
    input n39;
    input n41;
    input reset;
    input \data_in_frame[10][7] ;
    input \rx_data[7] ;
    input n60771;
    output n29190;
    input \data_in_frame[10][6] ;
    input n25647;
    input n25732;
    output n60896;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n63329, n22, n15, n20, n24, n19, n45_c, pwm_out_N_577, 
        n37, n23, n25, n29, n35, n11, n13, n27, n9, n17, 
        n19_adj_4430, n21, n15_adj_4431, n69216, n69167, n12, n30, 
        n69237, n70165, n59268, n54483, n59308, n54482, n70161, 
        n59340, n54481, n59380, n54480, n71225, n70611, n59420, 
        n54479, n59462, n54478, n71376, n59496, n54477, n59536, 
        n54476, n59568, n54475, n59604, n54474, n6, n70954, n70955, 
        n59630, n54473, n59656, n54472, n16, n24_adj_4433, n69013, 
        n59690, n54471, n8, n68970, n70756, n59730, n54470, n59780, 
        n54469, n59826, n54468, n69618, n59874, n54467, n59928, 
        n54466, n60018, n54465, n60132, n54464, n4, n60222, n54463, 
        n60220, n54462, n70760, n70761, n69147, n60218, n54461, 
        n60210, n10, n69134, n71235, n69616, n71486, n71487, n71391, 
        n69020, n71313, n70759, n71422;
    
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n63329));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[11]), .I1(\pwm_counter[16] ), .I2(\pwm_counter[19] ), 
            .I3(pwm_counter[18]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n63329), .I1(\pwm_counter[15] ), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(\pwm_counter[22] ), .I1(\pwm_counter[21] ), .I2(pwm_counter[14]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(\pwm_counter[20] ), .I3(pwm_counter[12]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[13]), .I1(pwm_counter[17]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(n45_c));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2881), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4430));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4431));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52126_4_lut (.I0(n21), .I1(n19_adj_4430), .I2(n17), .I3(n9), 
            .O(n69216));
    defparam i52126_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52077_4_lut (.I0(n27), .I1(n15_adj_4431), .I2(n13), .I3(n11), 
            .O(n69167));
    defparam i52077_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53075_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n69237), 
            .O(n70165));
    defparam i53075_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 pwm_counter_2040_add_4_25_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n54483), .O(n59268)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2040_add_4_24_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n54482), .O(n59308)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i53071_4_lut (.I0(n19_adj_4430), .I1(n17), .I2(n15_adj_4431), 
            .I3(n70165), .O(n70161));
    defparam i53071_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY pwm_counter_2040_add_4_24 (.CI(n54482), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n54483));
    SB_LUT4 pwm_counter_2040_add_4_23_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n54481), .O(n59340)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_23 (.CI(n54481), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n54482));
    SB_LUT4 pwm_counter_2040_add_4_22_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[20] ), 
            .I3(n54480), .O(n59380)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_22 (.CI(n54480), .I0(GND_net), .I1(\pwm_counter[20] ), 
            .CO(n54481));
    SB_LUT4 i54135_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n70161), 
            .O(n71225));
    defparam i54135_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53521_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n71225), 
            .O(n70611));
    defparam i53521_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 pwm_counter_2040_add_4_21_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n54479), .O(n59420)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_21 (.CI(n54479), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n54480));
    SB_LUT4 pwm_counter_2040_add_4_20_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n54478), .O(n59462)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_20 (.CI(n54478), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n54479));
    SB_LUT4 i54286_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n70611), 
            .O(n71376));
    defparam i54286_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_counter_2040_add_4_19_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n54477), .O(n59496)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_19 (.CI(n54477), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n54478));
    SB_LUT4 pwm_counter_2040_add_4_18_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[16] ), 
            .I3(n54476), .O(n59536)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_18 (.CI(n54476), .I0(GND_net), .I1(\pwm_counter[16] ), 
            .CO(n54477));
    SB_LUT4 pwm_counter_2040_add_4_17_lut (.I0(n45_c), .I1(GND_net), .I2(\pwm_counter[15] ), 
            .I3(n54475), .O(n59568)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_17 (.CI(n54475), .I0(GND_net), .I1(\pwm_counter[15] ), 
            .CO(n54476));
    SB_LUT4 pwm_counter_2040_add_4_16_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n54474), .O(n59604)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i53864_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n70954));   // verilog/pwm.v(21[8:24])
    defparam i53864_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY pwm_counter_2040_add_4_16 (.CI(n54474), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n54475));
    SB_LUT4 i53865_3_lut (.I0(n70954), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n70955));   // verilog/pwm.v(21[8:24])
    defparam i53865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_counter_2040_add_4_15_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n54473), .O(n59630)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_15 (.CI(n54473), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n54474));
    SB_LUT4 pwm_counter_2040_add_4_14_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n54472), .O(n59656)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4433));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY pwm_counter_2040_add_4_14 (.CI(n54472), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n54473));
    SB_LUT4 i51923_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n69216), 
            .O(n69013));
    defparam i51923_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_counter_2040_add_4_13_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n54471), .O(n59690)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_13 (.CI(n54471), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n54472));
    SB_LUT4 i53666_4_lut (.I0(n24_adj_4433), .I1(n8), .I2(n45), .I3(n68970), 
            .O(n70756));   // verilog/pwm.v(21[8:24])
    defparam i53666_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 pwm_counter_2040_add_4_12_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n54470), .O(n59730)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_12 (.CI(n54470), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n54471));
    SB_LUT4 pwm_counter_2040_add_4_11_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n54469), .O(n59780)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_11 (.CI(n54469), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n54470));
    SB_LUT4 pwm_counter_2040_add_4_10_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n54468), .O(n59826)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i52528_3_lut (.I0(n70955), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n69618));   // verilog/pwm.v(21[8:24])
    defparam i52528_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY pwm_counter_2040_add_4_10 (.CI(n54468), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n54469));
    SB_LUT4 pwm_counter_2040_add_4_9_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n54467), .O(n59874)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_9 (.CI(n54467), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n54468));
    SB_LUT4 pwm_counter_2040_add_4_8_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n54466), .O(n59928)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_8 (.CI(n54466), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n54467));
    SB_LUT4 pwm_counter_2040_add_4_7_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n54465), .O(n60018)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_7 (.CI(n54465), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n54466));
    SB_LUT4 pwm_counter_2040_add_4_6_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n54464), .O(n60132)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_6 (.CI(n54464), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n54465));
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 pwm_counter_2040_add_4_5_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n54463), .O(n60222)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_5 (.CI(n54463), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n54464));
    SB_LUT4 pwm_counter_2040_add_4_4_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n54462), .O(n60220)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i53670_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n70760));   // verilog/pwm.v(21[8:24])
    defparam i53670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53671_3_lut (.I0(n70760), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n70761));   // verilog/pwm.v(21[8:24])
    defparam i53671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52057_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n69167), 
            .O(n69147));
    defparam i52057_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY pwm_counter_2040_add_4_4 (.CI(n54462), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n54463));
    SB_LUT4 pwm_counter_2040_add_4_3_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n54461), .O(n60218)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_3 (.CI(n54461), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n54462));
    SB_LUT4 pwm_counter_2040_add_4_2_lut (.I0(n45_c), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n60210)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n54461));
    SB_LUT4 i54145_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n69134), 
            .O(n71235));   // verilog/pwm.v(21[8:24])
    defparam i54145_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52526_3_lut (.I0(n70761), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n69616));   // verilog/pwm.v(21[8:24])
    defparam i52526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54396_4_lut (.I0(n69616), .I1(n71235), .I2(n35), .I3(n69147), 
            .O(n71486));   // verilog/pwm.v(21[8:24])
    defparam i54396_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54397_3_lut (.I0(n71486), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n71487));   // verilog/pwm.v(21[8:24])
    defparam i54397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54301_3_lut (.I0(n71487), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n71391));   // verilog/pwm.v(21[8:24])
    defparam i54301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51930_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n71376), 
            .O(n69020));
    defparam i51930_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i54223_4_lut (.I0(n69618), .I1(n70756), .I2(n45), .I3(n69013), 
            .O(n71313));   // verilog/pwm.v(21[8:24])
    defparam i54223_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i53669_3_lut (.I0(n71391), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n70759));   // verilog/pwm.v(21[8:24])
    defparam i53669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i54332_4_lut (.I0(n70759), .I1(n71313), .I2(n45), .I3(n69020), 
            .O(n71422));   // verilog/pwm.v(21[8:24])
    defparam i54332_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i54333_3_lut (.I0(n71422), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i54333_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52147_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n69237));   // verilog/pwm.v(21[8:24])
    defparam i52147_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_DFFR pwm_counter_2040__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n60210), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_DFFR pwm_counter_2040__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n60218), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n60220), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n60222), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n60132), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n60018), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n59928), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n59874), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n59826), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n59780), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n59730), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n59690), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n59656), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n59630), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n59604), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i15 (.Q(\pwm_counter[15] ), .C(clk32MHz), 
            .D(n59568), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i16 (.Q(\pwm_counter[16] ), .C(clk32MHz), 
            .D(n59536), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n59496), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n59462), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n59420), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i20 (.Q(\pwm_counter[20] ), .C(clk32MHz), 
            .D(n59380), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n59340), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n59308), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n59268), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i13329_3_lut (.I0(\data_in_frame[10][7] ), .I1(\rx_data[7] ), 
            .I2(n60771), .I3(GND_net), .O(n29190));   // verilog/coms.v(130[12] 305[6])
    defparam i13329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51880_2_lut_4_lut (.I0(\pwm_counter[21] ), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n68970));
    defparam i51880_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(\pwm_counter[21] ), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52044_2_lut_4_lut (.I0(\pwm_counter[16] ), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n69134));
    defparam i52044_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(\pwm_counter[16] ), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[10][6] ), .I1(n25647), .I2(n25732), 
            .I3(GND_net), .O(n60896));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    
endmodule
